*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=0
.PARAM TCLOCK=1e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.1E-12 0.5E-09
ROUT Q 0  1
IT1|T 0 CLK  PWL(0 0 -3e-12 0 0 0.00105 3e-12 0 9.7e-11 0 1e-10 0.00105 1.03e-10 0 1.97e-10 0 2e-10 0.00105 2.03e-10 0 2.97e-10 0 3e-10 0.00105 3.03e-10 0 3.97e-10 0 4e-10 0.00105 4.03e-10 0 4.97e-10 0 5e-10 0.00105 5.03e-10 0 5.97e-10 0 6e-10 0.00105 6.03e-10 0 6.97e-10 0 7e-10 0.00105 7.03e-10 0 7.97e-10 0 8e-10 0.00105 8.03e-10 0 8.97e-10 0 9e-10 0.00105 9.03e-10 0 9.97e-10 0 1e-09 0.00105 1.003e-09 0 1.097e-09 0 1.1e-09 0.00105 1.103e-09 0 1.197e-09 0 1.2e-09 0.00105 1.203e-09 0 1.297e-09 0 1.3e-09 0.00105 1.303e-09 0 1.397e-09 0 1.4e-09 0.00105 1.403e-09 0 1.497e-09 0 1.5e-09 0.00105 1.503e-09 0 1.597e-09 0 1.6e-09 0.00105 1.603e-09 0 1.697e-09 0 1.7e-09 0.00105 1.703e-09 0 1.797e-09 0 1.8e-09 0.00105 1.803e-09 0 1.897e-09 0 1.9e-09 0.00105 1.903e-09 0 1.997e-09 0 2e-09 0.00105 2.003e-09 0 2.097e-09 0 2.1e-09 0.00105 2.103e-09 0 2.197e-09 0 2.2e-09 0.00105 2.203e-09 0 2.297e-09 0 2.3e-09 0.00105 2.303e-09 0 2.397e-09 0 2.4e-09 0.00105 2.403e-09 0 2.497e-09 0 2.5e-09 0.00105 2.503e-09 0 2.597e-09 0 2.6e-09 0.00105 2.603e-09 0 2.697e-09 0 2.7e-09 0.00105 2.703e-09 0 2.797e-09 0 2.8e-09 0.00105 2.803e-09 0 2.897e-09 0 2.9e-09 0.00105 2.903e-09 0 2.997e-09 0 3e-09 0.00105 3.003e-09 0 3.097e-09 0 3.1e-09 0.00105 3.103e-09 0 3.197e-09 0 3.2e-09 0.00105 3.203e-09 0 3.297e-09 0 3.3e-09 0.00105 3.303e-09 0 3.397e-09 0 3.4e-09 0.00105 3.403e-09 0 3.497e-09 0 3.5e-09 0.00105 3.503e-09 0 3.597e-09 0 3.6e-09 0.00105 3.603e-09 0 3.697e-09 0 3.7e-09 0.00105 3.703e-09 0 3.797e-09 0 3.8e-09 0.00105 3.803e-09 0 3.897e-09 0 3.9e-09 0.00105 3.903e-09 0 3.997e-09 0 4e-09 0.00105 4.003e-09 0 4.097e-09 0 4.1e-09 0.00105 4.103e-09 0 4.197e-09 0 4.2e-09 0.00105 4.203e-09 0 4.297e-09 0 4.3e-09 0.00105 4.303e-09 0 4.397e-09 0 4.4e-09 0.00105 4.403e-09 0 4.497e-09 0 4.5e-09 0.00105 4.503e-09 0 4.597e-09 0 4.6e-09 0.00105 4.603e-09 0 4.697e-09 0 4.7e-09 0.00105 4.703e-09 0 4.797e-09 0 4.8e-09 0.00105 4.803e-09 0 4.897e-09 0 4.9e-09 0.00105 4.903e-09 0 4.997e-09 0 5e-09 0.00105 5.003e-09 0 5.097e-09 0 5.1e-09 0.00105 5.103e-09 0 5.197e-09 0 5.2e-09 0.00105 5.203e-09 0 5.297e-09 0 5.3e-09 0.00105 5.303e-09 0 5.397e-09 0 5.4e-09 0.00105 5.403e-09 0 5.497e-09 0 5.5e-09 0.00105 5.503e-09 0 5.597e-09 0 5.6e-09 0.00105 5.603e-09 0 5.697e-09 0 5.7e-09 0.00105 5.703e-09 0 5.797e-09 0 5.8e-09 0.00105 5.803e-09 0 5.897e-09 0 5.9e-09 0.00105 5.903e-09 0 5.997e-09 0 6e-09 0.00105 6.003e-09 0 6.097e-09 0 6.1e-09 0.00105 6.103e-09 0 6.197e-09 0 6.2e-09 0.00105 6.203e-09 0 6.297e-09 0 6.3e-09 0.00105 6.303e-09 0 6.397e-09 0 6.4e-09 0.00105 6.403e-09 0 6.497e-09 0 6.5e-09 0.00105 6.503e-09 0 6.597e-09 0 6.6e-09 0.00105 6.603e-09 0 6.697e-09 0 6.7e-09 0.00105 6.703e-09 0 6.797e-09 0 6.8e-09 0.00105 6.803e-09 0 6.897e-09 0 6.9e-09 0.00105 6.903e-09 0 6.997e-09 0 7e-09 0.00105 7.003e-09 0 7.097e-09 0 7.1e-09 0.00105 7.103e-09 0 7.197e-09 0 7.2e-09 0.00105 7.203e-09 0 7.297e-09 0 7.3e-09 0.00105 7.303e-09 0 7.397e-09 0 7.4e-09 0.00105 7.403e-09 0 7.497e-09 0 7.5e-09 0.00105 7.503e-09 0 7.597e-09 0 7.6e-09 0.00105 7.603e-09 0 7.697e-09 0 7.7e-09 0.00105 7.703e-09 0 7.797e-09 0 7.8e-09 0.00105 7.803e-09 0 7.897e-09 0 7.9e-09 0.00105 7.903e-09 0 7.997e-09 0 8e-09 0.00105 8.003e-09 0 8.097e-09 0 8.1e-09 0.00105 8.103e-09 0 8.197e-09 0 8.2e-09 0.00105 8.203e-09 0 8.297e-09 0 8.3e-09 0.00105 8.303e-09 0 8.397e-09 0 8.4e-09 0.00105 8.403e-09 0 8.497e-09 0 8.5e-09 0.00105 8.503e-09 0 8.597e-09 0 8.6e-09 0.00105 8.603e-09 0 8.697e-09 0 8.7e-09 0.00105 8.703e-09 0 8.797e-09 0 8.8e-09 0.00105 8.803e-09 0 8.897e-09 0 8.9e-09 0.00105 8.903e-09 0 8.997e-09 0 9e-09 0.00105 9.003e-09 0 9.097e-09 0 9.1e-09 0.00105 9.103e-09 0 9.197e-09 0 9.2e-09 0.00105 9.203e-09 0 9.297e-09 0 9.3e-09 0.00105 9.303e-09 0 9.397e-09 0 9.4e-09 0.00105 9.403e-09 0 9.497e-09 0 9.5e-09 0.00105 9.503e-09 0 9.597e-09 0 9.6e-09 0.00105 9.603e-09 0 9.697e-09 0 9.7e-09 0.00105 9.703e-09 0 9.797e-09 0 9.8e-09 0.00105 9.803e-09 0 9.897e-09 0 9.9e-09 0.00105 9.903e-09 0 9.997e-09 0 1e-08 0.00105 1.0003e-08 0 1.0097e-08 0 1.01e-08 0.00105 1.0103e-08 0 1.0197e-08 0 1.02e-08 0.00105 1.0203e-08 0 1.0297e-08 0 1.03e-08 0.00105 1.0303e-08 0 1.0397e-08 0 1.04e-08 0.00105 1.0403e-08 0 1.0497e-08 0 1.05e-08 0.00105 1.0503e-08 0 1.0597e-08 0 1.06e-08 0.00105 1.0603e-08 0 1.0697e-08 0 1.07e-08 0.00105 1.0703e-08 0 1.0797e-08 0 1.08e-08 0.00105 1.0803e-08 0 1.0897e-08 0 1.09e-08 0.00105 1.0903e-08 0 1.0997e-08 0 1.1e-08 0.00105 1.1003e-08 0 1.1097e-08 0 1.11e-08 0.00105 1.1103e-08 0 1.1197e-08 0 1.12e-08 0.00105 1.1203e-08 0 1.1297e-08 0 1.13e-08 0.00105 1.1303e-08 0 1.1397e-08 0 1.14e-08 0.00105 1.1403e-08 0 1.1497e-08 0 1.15e-08 0.00105 1.1503e-08 0 1.1597e-08 0 1.16e-08 0.00105 1.1603e-08 0 1.1697e-08 0 1.17e-08 0.00105 1.1703e-08 0 1.1797e-08 0 1.18e-08 0.00105 1.1803e-08 0 1.1897e-08 0 1.19e-08 0.00105 1.1903e-08 0 1.1997e-08 0 1.2e-08 0.00105 1.2003e-08 0 1.2097e-08 0 1.21e-08 0.00105 1.2103e-08 0 1.2197e-08 0 1.22e-08 0.00105 1.2203e-08 0 1.2297e-08 0 1.23e-08 0.00105 1.2303e-08 0 1.2397e-08 0 1.24e-08 0.00105 1.2403e-08 0 1.2497e-08 0 1.25e-08 0.00105 1.2503e-08 0 1.2597e-08 0 1.26e-08 0.00105 1.2603e-08 0 1.2697e-08 0 1.27e-08 0.00105 1.2703e-08 0 1.2797e-08 0 1.28e-08 0.00105 1.2803e-08 0 1.2897e-08 0 1.29e-08 0.00105 1.2903e-08 0 1.2997e-08 0 1.3e-08 0.00105 1.3003e-08 0 1.3097e-08 0 1.31e-08 0.00105 1.3103e-08 0 1.3197e-08 0 1.32e-08 0.00105 1.3203e-08 0 1.3297e-08 0 1.33e-08 0.00105 1.3303e-08 0 1.3397e-08 0 1.34e-08 0.00105 1.3403e-08 0 1.3497e-08 0 1.35e-08 0.00105 1.3503e-08 0 1.3597e-08 0 1.36e-08 0.00105 1.3603e-08 0 1.3697e-08 0 1.37e-08 0.00105 1.3703e-08 0 1.3797e-08 0 1.38e-08 0.00105 1.3803e-08 0 1.3897e-08 0 1.39e-08 0.00105 1.3903e-08 0 1.3997e-08 0 1.4e-08 0.00105 1.4003e-08 0 1.4097e-08 0 1.41e-08 0.00105 1.4103e-08 0 1.4197e-08 0 1.42e-08 0.00105 1.4203e-08 0 1.4297e-08 0 1.43e-08 0.00105 1.4303e-08 0 1.4397e-08 0 1.44e-08 0.00105 1.4403e-08 0 1.4497e-08 0 1.45e-08 0.00105 1.4503e-08 0 1.4597e-08 0 1.46e-08 0.00105 1.4603e-08 0 1.4697e-08 0 1.47e-08 0.00105 1.4703e-08 0 1.4797e-08 0 1.48e-08 0.00105 1.4803e-08 0 1.4897e-08 0 1.49e-08 0.00105 1.4903e-08 0 1.4997e-08 0 1.5e-08 0.00105 1.5003e-08 0 1.5097e-08 0 1.51e-08 0.00105 1.5103e-08 0 1.5197e-08 0 1.52e-08 0.00105 1.5203e-08 0 1.5297e-08 0 1.53e-08 0.00105 1.5303e-08 0 1.5397e-08 0 1.54e-08 0.00105 1.5403e-08 0 1.5497e-08 0 1.55e-08 0.00105 1.5503e-08 0 1.5597e-08 0 1.56e-08 0.00105 1.5603e-08 0 1.5697e-08 0 1.57e-08 0.00105 1.5703e-08 0 1.5797e-08 0 1.58e-08 0.00105 1.5803e-08 0 1.5897e-08 0 1.59e-08 0.00105 1.5903e-08 0 1.5997e-08 0 1.6e-08 0.00105 1.6003e-08 0 1.6097e-08 0 1.61e-08 0.00105 1.6103e-08 0 1.6197e-08 0 1.62e-08 0.00105 1.6203e-08 0 1.6297e-08 0 1.63e-08 0.00105 1.6303e-08 0 1.6397e-08 0 1.64e-08 0.00105 1.6403e-08 0 1.6497e-08 0 1.65e-08 0.00105 1.6503e-08 0 1.6597e-08 0 1.66e-08 0.00105 1.6603e-08 0 1.6697e-08 0 1.67e-08 0.00105 1.6703e-08 0 1.6797e-08 0 1.68e-08 0.00105 1.6803e-08 0 1.6897e-08 0 1.69e-08 0.00105 1.6903e-08 0 1.6997e-08 0 1.7e-08 0.00105 1.7003e-08 0 1.7097e-08 0 1.71e-08 0.00105 1.7103e-08 0 1.7197e-08 0 1.72e-08 0.00105 1.7203e-08 0 1.7297e-08 0 1.73e-08 0.00105 1.7303e-08 0 1.7397e-08 0 1.74e-08 0.00105 1.7403e-08 0 1.7497e-08 0 1.75e-08 0.00105 1.7503e-08 0 1.7597e-08 0 1.76e-08 0.00105 1.7603e-08 0 1.7697e-08 0 1.77e-08 0.00105 1.7703e-08 0 1.7797e-08 0 1.78e-08 0.00105 1.7803e-08 0 1.7897e-08 0 1.79e-08 0.00105 1.7903e-08 0 1.7997e-08 0 1.8e-08 0.00105 1.8003e-08 0 1.8097e-08 0 1.81e-08 0.00105 1.8103e-08 0 1.8197e-08 0 1.82e-08 0.00105 1.8203e-08 0 1.8297e-08 0 1.83e-08 0.00105 1.8303e-08 0 1.8397e-08 0 1.84e-08 0.00105 1.8403e-08 0 1.8497e-08 0 1.85e-08 0.00105 1.8503e-08 0 1.8597e-08 0 1.86e-08 0.00105 1.8603e-08 0 1.8697e-08 0 1.87e-08 0.00105 1.8703e-08 0 1.8797e-08 0 1.88e-08 0.00105 1.8803e-08 0 1.8897e-08 0 1.89e-08 0.00105 1.8903e-08 0 1.8997e-08 0 1.9e-08 0.00105 1.9003e-08 0 1.9097e-08 0 1.91e-08 0.00105 1.9103e-08 0 1.9197e-08 0 1.92e-08 0.00105 1.9203e-08 0 1.9297e-08 0 1.93e-08 0.00105 1.9303e-08 0 1.9397e-08 0 1.94e-08 0.00105 1.9403e-08 0 1.9497e-08 0 1.95e-08 0.00105 1.9503e-08 0 1.9597e-08 0 1.96e-08 0.00105 1.9603e-08 0 1.9697e-08 0 1.97e-08 0.00105 1.9703e-08 0 1.9797e-08 0 1.98e-08 0.00105 1.9803e-08 0 1.9897e-08 0 1.99e-08 0.00105 1.9903e-08 0 1.9997e-08 0 2e-08 0.00105 2.0003e-08 0 2.0097e-08 0 2.01e-08 0.00105 2.0103e-08 0 2.0197e-08 0 2.02e-08 0.00105 2.0203e-08 0 2.0297e-08 0 2.03e-08 0.00105 2.0303e-08 0 2.0397e-08 0 2.04e-08 0.00105 2.0403e-08 0 2.0497e-08 0 2.05e-08 0.00105 2.0503e-08 0 2.0597e-08 0 2.06e-08 0.00105 2.0603e-08 0 2.0697e-08 0 2.07e-08 0.00105 2.0703e-08 0 2.0797e-08 0 2.08e-08 0.00105 2.0803e-08 0 2.0897e-08 0 2.09e-08 0.00105 2.0903e-08 0 2.0997e-08 0 2.1e-08 0.00105 2.1003e-08 0 2.1097e-08 0 2.11e-08 0.00105 2.1103e-08 0 2.1197e-08 0 2.12e-08 0.00105 2.1203e-08 0 2.1297e-08 0 2.13e-08 0.00105 2.1303e-08 0 2.1397e-08 0 2.14e-08 0.00105 2.1403e-08 0 2.1497e-08 0 2.15e-08 0.00105 2.1503e-08 0 2.1597e-08 0 2.16e-08 0.00105 2.1603e-08 0 2.1697e-08 0 2.17e-08 0.00105 2.1703e-08 0 2.1797e-08 0 2.18e-08 0.00105 2.1803e-08 0 2.1897e-08 0 2.19e-08 0.00105 2.1903e-08 0 2.1997e-08 0 2.2e-08 0.00105 2.2003e-08 0 2.2097e-08 0 2.21e-08 0.00105 2.2103e-08 0 2.2197e-08 0 2.22e-08 0.00105 2.2203e-08 0 2.2297e-08 0 2.23e-08 0.00105 2.2303e-08 0 2.2397e-08 0 2.24e-08 0.00105 2.2403e-08 0 2.2497e-08 0 2.25e-08 0.00105 2.2503e-08 0 2.2597e-08 0 2.26e-08 0.00105 2.2603e-08 0 2.2697e-08 0 2.27e-08 0.00105 2.2703e-08 0 2.2797e-08 0 2.28e-08 0.00105 2.2803e-08 0 2.2897e-08 0 2.29e-08 0.00105 2.2903e-08 0 2.2997e-08 0 2.3e-08 0.00105 2.3003e-08 0 2.3097e-08 0 2.31e-08 0.00105 2.3103e-08 0 2.3197e-08 0 2.32e-08 0.00105 2.3203e-08 0 2.3297e-08 0 2.33e-08 0.00105 2.3303e-08 0 2.3397e-08 0 2.34e-08 0.00105 2.3403e-08 0 2.3497e-08 0 2.35e-08 0.00105 2.3503e-08 0 2.3597e-08 0 2.36e-08 0.00105 2.3603e-08 0 2.3697e-08 0 2.37e-08 0.00105 2.3703e-08 0 2.3797e-08 0 2.38e-08 0.00105 2.3803e-08 0 2.3897e-08 0 2.39e-08 0.00105 2.3903e-08 0 2.3997e-08 0 2.4e-08 0.00105 2.4003e-08 0 2.4097e-08 0 2.41e-08 0.00105 2.4103e-08 0 2.4197e-08 0 2.42e-08 0.00105 2.4203e-08 0 2.4297e-08 0 2.43e-08 0.00105 2.4303e-08 0 2.4397e-08 0 2.44e-08 0.00105 2.4403e-08 0 2.4497e-08 0 2.45e-08 0.00105 2.4503e-08 0 2.4597e-08 0 2.46e-08 0.00105 2.4603e-08 0 2.4697e-08 0 2.47e-08 0.00105 2.4703e-08 0 2.4797e-08 0 2.48e-08 0.00105 2.4803e-08 0 2.4897e-08 0 2.49e-08 0.00105 2.4903e-08 0 2.4997e-08 0 2.5e-08 0.00105 2.5003e-08 0 2.5097e-08 0 2.51e-08 0.00105 2.5103e-08 0 2.5197e-08 0 2.52e-08 0.00105 2.5203e-08 0 2.5297e-08 0 2.53e-08 0.00105 2.5303e-08 0 2.5397e-08 0 2.54e-08 0.00105 2.5403e-08 0 2.5497e-08 0 2.55e-08 0.00105 2.5503e-08 0 2.5597e-08 0 2.56e-08 0.00105 2.5603e-08 0 2.5697e-08 0 2.57e-08 0.00105 2.5703e-08 0 2.5797e-08 0 2.58e-08 0.00105 2.5803e-08 0 2.5897e-08 0 2.59e-08 0.00105 2.5903e-08 0 2.5997e-08 0 2.6e-08 0.00105 2.6003e-08 0 2.6097e-08 0 2.61e-08 0.00105 2.6103e-08 0 2.6197e-08 0 2.62e-08 0.00105 2.6203e-08 0 2.6297e-08 0 2.63e-08 0.00105 2.6303e-08 0 2.6397e-08 0 2.64e-08 0.00105 2.6403e-08 0 2.6497e-08 0 2.65e-08 0.00105 2.6503e-08 0 2.6597e-08 0 2.66e-08 0.00105 2.6603e-08 0 2.6697e-08 0 2.67e-08 0.00105 2.6703e-08 0 2.6797e-08 0 2.68e-08 0.00105 2.6803e-08 0 2.6897e-08 0 2.69e-08 0.00105 2.6903e-08 0 2.6997e-08 0 2.7e-08 0.00105 2.7003e-08 0 2.7097e-08 0 2.71e-08 0.00105 2.7103e-08 0 2.7197e-08 0 2.72e-08 0.00105 2.7203e-08 0 2.7297e-08 0 2.73e-08 0.00105 2.7303e-08 0 2.7397e-08 0 2.74e-08 0.00105 2.7403e-08 0 2.7497e-08 0 2.75e-08 0.00105 2.7503e-08 0 2.7597e-08 0 2.76e-08 0.00105 2.7603e-08 0 2.7697e-08 0 2.77e-08 0.00105 2.7703e-08 0 2.7797e-08 0 2.78e-08 0.00105 2.7803e-08 0 2.7897e-08 0 2.79e-08 0.00105 2.7903e-08 0 2.7997e-08 0 2.8e-08 0.00105 2.8003e-08 0 2.8097e-08 0 2.81e-08 0.00105 2.8103e-08 0 2.8197e-08 0 2.82e-08 0.00105 2.8203e-08 0 2.8297e-08 0 2.83e-08 0.00105 2.8303e-08 0 2.8397e-08 0 2.84e-08 0.00105 2.8403e-08 0 2.8497e-08 0 2.85e-08 0.00105 2.8503e-08 0 2.8597e-08 0 2.86e-08 0.00105 2.8603e-08 0 2.8697e-08 0 2.87e-08 0.00105 2.8703e-08 0 2.8797e-08 0 2.88e-08 0.00105 2.8803e-08 0 2.8897e-08 0 2.89e-08 0.00105 2.8903e-08 0 2.8997e-08 0 2.9e-08 0.00105 2.9003e-08 0 2.9097e-08 0 2.91e-08 0.00105 2.9103e-08 0 2.9197e-08 0 2.92e-08 0.00105 2.9203e-08 0 2.9297e-08 0 2.93e-08 0.00105 2.9303e-08 0 2.9397e-08 0 2.94e-08 0.00105 2.9403e-08 0 2.9497e-08 0 2.95e-08 0.00105 2.9503e-08 0 2.9597e-08 0 2.96e-08 0.00105 2.9603e-08 0 2.9697e-08 0 2.97e-08 0.00105 2.9703e-08 0 2.9797e-08 0 2.98e-08 0.00105 2.9803e-08 0 2.9897e-08 0 2.99e-08 0.00105 2.9903e-08 0 2.9997e-08 0 3e-08 0.00105 3.0003e-08 0 3.0097e-08 0 3.01e-08 0.00105 3.0103e-08 0 3.0197e-08 0 3.02e-08 0.00105 3.0203e-08 0 3.0297e-08 0 3.03e-08 0.00105 3.0303e-08 0 3.0397e-08 0 3.04e-08 0.00105 3.0403e-08 0 3.0497e-08 0 3.05e-08 0.00105 3.0503e-08 0 3.0597e-08 0 3.06e-08 0.00105 3.0603e-08 0 3.0697e-08 0 3.07e-08 0.00105 3.0703e-08 0 3.0797e-08 0 3.08e-08 0.00105 3.0803e-08 0 3.0897e-08 0 3.09e-08 0.00105 3.0903e-08 0 3.0997e-08 0 3.1e-08 0.00105 3.1003e-08 0 3.1097e-08 0 3.11e-08 0.00105 3.1103e-08 0 3.1197e-08 0 3.12e-08 0.00105 3.1203e-08 0 3.1297e-08 0 3.13e-08 0.00105 3.1303e-08 0 3.1397e-08 0 3.14e-08 0.00105 3.1403e-08 0 3.1497e-08 0 3.15e-08 0.00105 3.1503e-08 0 3.1597e-08 0 3.16e-08 0.00105 3.1603e-08 0 3.1697e-08 0 3.17e-08 0.00105 3.1703e-08 0 3.1797e-08 0 3.18e-08 0.00105 3.1803e-08 0 3.1897e-08 0 3.19e-08 0.00105 3.1903e-08 0 3.1997e-08 0 3.2e-08 0.00105 3.2003e-08 0 3.2097e-08 0 3.21e-08 0.00105 3.2103e-08 0 3.2197e-08 0 3.22e-08 0.00105 3.2203e-08 0 3.2297e-08 0 3.23e-08 0.00105 3.2303e-08 0 3.2397e-08 0 3.24e-08 0.00105 3.2403e-08 0 3.2497e-08 0 3.25e-08 0.00105 3.2503e-08 0 3.2597e-08 0 3.26e-08 0.00105 3.2603e-08 0 3.2697e-08 0 3.27e-08 0.00105 3.2703e-08 0 3.2797e-08 0 3.28e-08 0.00105 3.2803e-08 0 3.2897e-08 0 3.29e-08 0.00105 3.2903e-08 0 3.2997e-08 0 3.3e-08 0.00105 3.3003e-08 0 3.3097e-08 0 3.31e-08 0.00105 3.3103e-08 0 3.3197e-08 0 3.32e-08 0.00105 3.3203e-08 0 3.3297e-08 0 3.33e-08 0.00105 3.3303e-08 0 3.3397e-08 0 3.34e-08 0.00105 3.3403e-08 0 3.3497e-08 0 3.35e-08 0.00105 3.3503e-08 0 3.3597e-08 0 3.36e-08 0.00105 3.3603e-08 0 3.3697e-08 0 3.37e-08 0.00105 3.3703e-08 0 3.3797e-08 0 3.38e-08 0.00105 3.3803e-08 0 3.3897e-08 0 3.39e-08 0.00105 3.3903e-08 0 3.3997e-08 0 3.4e-08 0.00105 3.4003e-08 0 3.4097e-08 0 3.41e-08 0.00105 3.4103e-08 0 3.4197e-08 0 3.42e-08 0.00105 3.4203e-08 0 3.4297e-08 0 3.43e-08 0.00105 3.4303e-08 0 3.4397e-08 0 3.44e-08 0.00105 3.4403e-08 0 3.4497e-08 0 3.45e-08 0.00105 3.4503e-08 0 3.4597e-08 0 3.46e-08 0.00105 3.4603e-08 0 3.4697e-08 0 3.47e-08 0.00105 3.4703e-08 0 3.4797e-08 0 3.48e-08 0.00105 3.4803e-08 0 3.4897e-08 0 3.49e-08 0.00105 3.4903e-08 0 3.4997e-08 0 3.5e-08 0.00105 3.5003e-08 0 3.5097e-08 0 3.51e-08 0.00105 3.5103e-08 0 3.5197e-08 0 3.52e-08 0.00105 3.5203e-08 0 3.5297e-08 0 3.53e-08 0.00105 3.5303e-08 0 3.5397e-08 0 3.54e-08 0.00105 3.5403e-08 0 3.5497e-08 0 3.55e-08 0.00105 3.5503e-08 0 3.5597e-08 0 3.56e-08 0.00105 3.5603e-08 0 3.5697e-08 0 3.57e-08 0.00105 3.5703e-08 0 3.5797e-08 0 3.58e-08 0.00105 3.5803e-08 0 3.5897e-08 0 3.59e-08 0.00105 3.5903e-08 0 3.5997e-08 0 3.6e-08 0.00105 3.6003e-08 0 3.6097e-08 0 3.61e-08 0.00105 3.6103e-08 0 3.6197e-08 0 3.62e-08 0.00105 3.6203e-08 0 3.6297e-08 0 3.63e-08 0.00105 3.6303e-08 0 3.6397e-08 0 3.64e-08 0.00105 3.6403e-08 0 3.6497e-08 0 3.65e-08 0.00105 3.6503e-08 0 3.6597e-08 0 3.66e-08 0.00105 3.6603e-08 0 3.6697e-08 0 3.67e-08 0.00105 3.6703e-08 0 3.6797e-08 0 3.68e-08 0.00105 3.6803e-08 0 3.6897e-08 0 3.69e-08 0.00105 3.6903e-08 0 3.6997e-08 0 3.7e-08 0.00105 3.7003e-08 0 3.7097e-08 0 3.71e-08 0.00105 3.7103e-08 0 3.7197e-08 0 3.72e-08 0.00105 3.7203e-08 0 3.7297e-08 0 3.73e-08 0.00105 3.7303e-08 0 3.7397e-08 0 3.74e-08 0.00105 3.7403e-08 0 3.7497e-08 0 3.75e-08 0.00105 3.7503e-08 0 3.7597e-08 0 3.76e-08 0.00105 3.7603e-08 0 3.7697e-08 0 3.77e-08 0.00105 3.7703e-08 0 3.7797e-08 0 3.78e-08 0.00105 3.7803e-08 0 3.7897e-08 0 3.79e-08 0.00105 3.7903e-08 0 3.7997e-08 0 3.8e-08 0.00105 3.8003e-08 0 3.8097e-08 0 3.81e-08 0.00105 3.8103e-08 0 3.8197e-08 0 3.82e-08 0.00105 3.8203e-08 0 3.8297e-08 0 3.83e-08 0.00105 3.8303e-08 0 3.8397e-08 0 3.84e-08 0.00105 3.8403e-08 0 3.8497e-08 0 3.85e-08 0.00105 3.8503e-08 0 3.8597e-08 0 3.86e-08 0.00105 3.8603e-08 0 3.8697e-08 0 3.87e-08 0.00105 3.8703e-08 0 3.8797e-08 0 3.88e-08 0.00105 3.8803e-08 0 3.8897e-08 0 3.89e-08 0.00105 3.8903e-08 0 3.8997e-08 0 3.9e-08 0.00105 3.9003e-08 0 3.9097e-08 0 3.91e-08 0.00105 3.9103e-08 0 3.9197e-08 0 3.92e-08 0.00105 3.9203e-08 0 3.9297e-08 0 3.93e-08 0.00105 3.9303e-08 0 3.9397e-08 0 3.94e-08 0.00105 3.9403e-08 0 3.9497e-08 0 3.95e-08 0.00105 3.9503e-08 0 3.9597e-08 0 3.96e-08 0.00105 3.9603e-08 0 3.9697e-08 0 3.97e-08 0.00105 3.9703e-08 0 3.9797e-08 0 3.98e-08 0.00105 3.9803e-08 0)
IDATA_A1|A 0 A  PWL(0 0 1.637e-10 0 1.667e-10 0.0007 1.697e-10 0 3.637e-10 0 3.667e-10 0.0007 3.697e-10 0 5.637e-10 0 5.667e-10 0.0007 5.697e-10 0 7.637e-10 0 7.667e-10 0.0007 7.697e-10 0 9.637e-10 0 9.667e-10 0.0007 9.697e-10 0 1.1637e-09 0 1.1667e-09 0.0007 1.1697e-09 0 1.3637e-09 0 1.3667e-09 0.0007 1.3697e-09 0 1.5637e-09 0 1.5667e-09 0.0007 1.5697e-09 0 1.7637e-09 0 1.7667e-09 0.0007 1.7697e-09 0 1.9637e-09 0 1.9667e-09 0.0007 1.9697e-09 0 2.1637e-09 0 2.1667e-09 0.0007 2.1697e-09 0 2.3637e-09 0 2.3667e-09 0.0007 2.3697e-09 0 2.5637e-09 0 2.5667e-09 0.0007 2.5697e-09 0 2.7637e-09 0 2.7667e-09 0.0007 2.7697e-09 0 2.9637e-09 0 2.9667e-09 0.0007 2.9697e-09 0 3.1637e-09 0 3.1667e-09 0.0007 3.1697e-09 0 3.3637e-09 0 3.3667e-09 0.0007 3.3697e-09 0 3.5637e-09 0 3.5667e-09 0.0007 3.5697e-09 0 3.7637e-09 0 3.7667e-09 0.0007 3.7697e-09 0 3.9637e-09 0 3.9667e-09 0.0007 3.9697e-09 0 4.1637e-09 0 4.1667e-09 0.0007 4.1697e-09 0 4.3637e-09 0 4.3667e-09 0.0007 4.3697e-09 0 4.5637e-09 0 4.5667e-09 0.0007 4.5697e-09 0 4.7637e-09 0 4.7667e-09 0.0007 4.7697e-09 0 4.9637e-09 0 4.9667e-09 0.0007 4.9697e-09 0 5.1637e-09 0 5.1667e-09 0.0007 5.1697e-09 0 5.3637e-09 0 5.3667e-09 0.0007 5.3697e-09 0 5.5637e-09 0 5.5667e-09 0.0007 5.5697e-09 0 5.7637e-09 0 5.7667e-09 0.0007 5.7697e-09 0 5.9637e-09 0 5.9667e-09 0.0007 5.9697e-09 0 6.1637e-09 0 6.1667e-09 0.0007 6.1697e-09 0 6.3637e-09 0 6.3667e-09 0.0007 6.3697e-09 0 6.5637e-09 0 6.5667e-09 0.0007 6.5697e-09 0 6.7637e-09 0 6.7667e-09 0.0007 6.7697e-09 0 6.9637e-09 0 6.9667e-09 0.0007 6.9697e-09 0 7.1637e-09 0 7.1667e-09 0.0007 7.1697e-09 0 7.3637e-09 0 7.3667e-09 0.0007 7.3697e-09 0 7.5637e-09 0 7.5667e-09 0.0007 7.5697e-09 0 7.7637e-09 0 7.7667e-09 0.0007 7.7697e-09 0 7.9637e-09 0 7.9667e-09 0.0007 7.9697e-09 0 8.1637e-09 0 8.1667e-09 0.0007 8.1697e-09 0 8.3637e-09 0 8.3667e-09 0.0007 8.3697e-09 0 8.5637e-09 0 8.5667e-09 0.0007 8.5697e-09 0 8.7637e-09 0 8.7667e-09 0.0007 8.7697e-09 0 8.9637e-09 0 8.9667e-09 0.0007 8.9697e-09 0 9.1637e-09 0 9.1667e-09 0.0007 9.1697e-09 0 9.3637e-09 0 9.3667e-09 0.0007 9.3697e-09 0 9.5637e-09 0 9.5667e-09 0.0007 9.5697e-09 0 9.7637e-09 0 9.7667e-09 0.0007 9.7697e-09 0 9.9637e-09 0 9.9667e-09 0.0007 9.9697e-09 0 1.01637e-08 0 1.01667e-08 0.0007 1.01697e-08 0 1.03637e-08 0 1.03667e-08 0.0007 1.03697e-08 0 1.05637e-08 0 1.05667e-08 0.0007 1.05697e-08 0 1.07637e-08 0 1.07667e-08 0.0007 1.07697e-08 0 1.09637e-08 0 1.09667e-08 0.0007 1.09697e-08 0 1.11637e-08 0 1.11667e-08 0.0007 1.11697e-08 0 1.13637e-08 0 1.13667e-08 0.0007 1.13697e-08 0 1.15637e-08 0 1.15667e-08 0.0007 1.15697e-08 0 1.17637e-08 0 1.17667e-08 0.0007 1.17697e-08 0 1.19637e-08 0 1.19667e-08 0.0007 1.19697e-08 0 1.21637e-08 0 1.21667e-08 0.0007 1.21697e-08 0 1.23637e-08 0 1.23667e-08 0.0007 1.23697e-08 0 1.25637e-08 0 1.25667e-08 0.0007 1.25697e-08 0 1.27637e-08 0 1.27667e-08 0.0007 1.27697e-08 0 1.29637e-08 0 1.29667e-08 0.0007 1.29697e-08 0 1.31637e-08 0 1.31667e-08 0.0007 1.31697e-08 0 1.33637e-08 0 1.33667e-08 0.0007 1.33697e-08 0 1.35637e-08 0 1.35667e-08 0.0007 1.35697e-08 0 1.37637e-08 0 1.37667e-08 0.0007 1.37697e-08 0 1.39637e-08 0 1.39667e-08 0.0007 1.39697e-08 0 1.41637e-08 0 1.41667e-08 0.0007 1.41697e-08 0 1.43637e-08 0 1.43667e-08 0.0007 1.43697e-08 0 1.45637e-08 0 1.45667e-08 0.0007 1.45697e-08 0 1.47637e-08 0 1.47667e-08 0.0007 1.47697e-08 0 1.49637e-08 0 1.49667e-08 0.0007 1.49697e-08 0 1.51637e-08 0 1.51667e-08 0.0007 1.51697e-08 0 1.53637e-08 0 1.53667e-08 0.0007 1.53697e-08 0 1.55637e-08 0 1.55667e-08 0.0007 1.55697e-08 0 1.57637e-08 0 1.57667e-08 0.0007 1.57697e-08 0 1.59637e-08 0 1.59667e-08 0.0007 1.59697e-08 0 1.61637e-08 0 1.61667e-08 0.0007 1.61697e-08 0 1.63637e-08 0 1.63667e-08 0.0007 1.63697e-08 0 1.65637e-08 0 1.65667e-08 0.0007 1.65697e-08 0 1.67637e-08 0 1.67667e-08 0.0007 1.67697e-08 0 1.69637e-08 0 1.69667e-08 0.0007 1.69697e-08 0 1.71637e-08 0 1.71667e-08 0.0007 1.71697e-08 0 1.73637e-08 0 1.73667e-08 0.0007 1.73697e-08 0 1.75637e-08 0 1.75667e-08 0.0007 1.75697e-08 0 1.77637e-08 0 1.77667e-08 0.0007 1.77697e-08 0 1.79637e-08 0 1.79667e-08 0.0007 1.79697e-08 0 1.81637e-08 0 1.81667e-08 0.0007 1.81697e-08 0 1.83637e-08 0 1.83667e-08 0.0007 1.83697e-08 0 1.85637e-08 0 1.85667e-08 0.0007 1.85697e-08 0 1.87637e-08 0 1.87667e-08 0.0007 1.87697e-08 0 1.89637e-08 0 1.89667e-08 0.0007 1.89697e-08 0 1.91637e-08 0 1.91667e-08 0.0007 1.91697e-08 0 1.93637e-08 0 1.93667e-08 0.0007 1.93697e-08 0 1.95637e-08 0 1.95667e-08 0.0007 1.95697e-08 0 1.97637e-08 0 1.97667e-08 0.0007 1.97697e-08 0 1.99637e-08 0 1.99667e-08 0.0007 1.99697e-08 0 2.01637e-08 0 2.01667e-08 0.0007 2.01697e-08 0 2.03637e-08 0 2.03667e-08 0.0007 2.03697e-08 0 2.05637e-08 0 2.05667e-08 0.0007 2.05697e-08 0 2.07637e-08 0 2.07667e-08 0.0007 2.07697e-08 0 2.09637e-08 0 2.09667e-08 0.0007 2.09697e-08 0 2.11637e-08 0 2.11667e-08 0.0007 2.11697e-08 0 2.13637e-08 0 2.13667e-08 0.0007 2.13697e-08 0 2.15637e-08 0 2.15667e-08 0.0007 2.15697e-08 0 2.17637e-08 0 2.17667e-08 0.0007 2.17697e-08 0 2.19637e-08 0 2.19667e-08 0.0007 2.19697e-08 0 2.21637e-08 0 2.21667e-08 0.0007 2.21697e-08 0 2.23637e-08 0 2.23667e-08 0.0007 2.23697e-08 0 2.25637e-08 0 2.25667e-08 0.0007 2.25697e-08 0 2.27637e-08 0 2.27667e-08 0.0007 2.27697e-08 0 2.29637e-08 0 2.29667e-08 0.0007 2.29697e-08 0 2.31637e-08 0 2.31667e-08 0.0007 2.31697e-08 0 2.33637e-08 0 2.33667e-08 0.0007 2.33697e-08 0 2.35637e-08 0 2.35667e-08 0.0007 2.35697e-08 0 2.37637e-08 0 2.37667e-08 0.0007 2.37697e-08 0 2.39637e-08 0 2.39667e-08 0.0007 2.39697e-08 0 2.41637e-08 0 2.41667e-08 0.0007 2.41697e-08 0 2.43637e-08 0 2.43667e-08 0.0007 2.43697e-08 0 2.45637e-08 0 2.45667e-08 0.0007 2.45697e-08 0 2.47637e-08 0 2.47667e-08 0.0007 2.47697e-08 0 2.49637e-08 0 2.49667e-08 0.0007 2.49697e-08 0 2.51637e-08 0 2.51667e-08 0.0007 2.51697e-08 0 2.53637e-08 0 2.53667e-08 0.0007 2.53697e-08 0 2.55637e-08 0 2.55667e-08 0.0007 2.55697e-08 0)
IDATA_B1|B 0 B  PWL(0 0 2.303e-10 0 2.333e-10 0.0007 2.363e-10 0 3.303e-10 0 3.333e-10 0.0007 3.363e-10 0 6.303e-10 0 6.333e-10 0.0007 6.363e-10 0 7.303e-10 0 7.333e-10 0.0007 7.363e-10 0 1.0303e-09 0 1.0333e-09 0.0007 1.0363e-09 0 1.1303e-09 0 1.1333e-09 0.0007 1.1363e-09 0 1.4303e-09 0 1.4333e-09 0.0007 1.4363e-09 0 1.5303e-09 0 1.5333e-09 0.0007 1.5363e-09 0 1.8303e-09 0 1.8333e-09 0.0007 1.8363e-09 0 1.9303e-09 0 1.9333e-09 0.0007 1.9363e-09 0 2.2303e-09 0 2.2333e-09 0.0007 2.2363e-09 0 2.3303e-09 0 2.3333e-09 0.0007 2.3363e-09 0 2.6303e-09 0 2.6333e-09 0.0007 2.6363e-09 0 2.7303e-09 0 2.7333e-09 0.0007 2.7363e-09 0 3.0303e-09 0 3.0333e-09 0.0007 3.0363e-09 0 3.1303e-09 0 3.1333e-09 0.0007 3.1363e-09 0 3.4303e-09 0 3.4333e-09 0.0007 3.4363e-09 0 3.5303e-09 0 3.5333e-09 0.0007 3.5363e-09 0 3.8303e-09 0 3.8333e-09 0.0007 3.8363e-09 0 3.9303e-09 0 3.9333e-09 0.0007 3.9363e-09 0 4.2303e-09 0 4.2333e-09 0.0007 4.2363e-09 0 4.3303e-09 0 4.3333e-09 0.0007 4.3363e-09 0 4.6303e-09 0 4.6333e-09 0.0007 4.6363e-09 0 4.7303e-09 0 4.7333e-09 0.0007 4.7363e-09 0 5.0303e-09 0 5.0333e-09 0.0007 5.0363e-09 0 5.1303e-09 0 5.1333e-09 0.0007 5.1363e-09 0 5.4303e-09 0 5.4333e-09 0.0007 5.4363e-09 0 5.5303e-09 0 5.5333e-09 0.0007 5.5363e-09 0 5.8303e-09 0 5.8333e-09 0.0007 5.8363e-09 0 5.9303e-09 0 5.9333e-09 0.0007 5.9363e-09 0 6.2303e-09 0 6.2333e-09 0.0007 6.2363e-09 0 6.3303e-09 0 6.3333e-09 0.0007 6.3363e-09 0 6.6303e-09 0 6.6333e-09 0.0007 6.6363e-09 0 6.7303e-09 0 6.7333e-09 0.0007 6.7363e-09 0 7.0303e-09 0 7.0333e-09 0.0007 7.0363e-09 0 7.1303e-09 0 7.1333e-09 0.0007 7.1363e-09 0 7.4303e-09 0 7.4333e-09 0.0007 7.4363e-09 0 7.5303e-09 0 7.5333e-09 0.0007 7.5363e-09 0 7.8303e-09 0 7.8333e-09 0.0007 7.8363e-09 0 7.9303e-09 0 7.9333e-09 0.0007 7.9363e-09 0 8.2303e-09 0 8.2333e-09 0.0007 8.2363e-09 0 8.3303e-09 0 8.3333e-09 0.0007 8.3363e-09 0 8.6303e-09 0 8.6333e-09 0.0007 8.6363e-09 0 8.7303e-09 0 8.7333e-09 0.0007 8.7363e-09 0 9.0303e-09 0 9.0333e-09 0.0007 9.0363e-09 0 9.1303e-09 0 9.1333e-09 0.0007 9.1363e-09 0 9.4303e-09 0 9.4333e-09 0.0007 9.4363e-09 0 9.5303e-09 0 9.5333e-09 0.0007 9.5363e-09 0 9.8303e-09 0 9.8333e-09 0.0007 9.8363e-09 0 9.9303e-09 0 9.9333e-09 0.0007 9.9363e-09 0 1.02303e-08 0 1.02333e-08 0.0007 1.02363e-08 0 1.03303e-08 0 1.03333e-08 0.0007 1.03363e-08 0 1.06303e-08 0 1.06333e-08 0.0007 1.06363e-08 0 1.07303e-08 0 1.07333e-08 0.0007 1.07363e-08 0 1.10303e-08 0 1.10333e-08 0.0007 1.10363e-08 0 1.11303e-08 0 1.11333e-08 0.0007 1.11363e-08 0 1.14303e-08 0 1.14333e-08 0.0007 1.14363e-08 0 1.15303e-08 0 1.15333e-08 0.0007 1.15363e-08 0 1.18303e-08 0 1.18333e-08 0.0007 1.18363e-08 0 1.19303e-08 0 1.19333e-08 0.0007 1.19363e-08 0 1.22303e-08 0 1.22333e-08 0.0007 1.22363e-08 0 1.23303e-08 0 1.23333e-08 0.0007 1.23363e-08 0 1.26303e-08 0 1.26333e-08 0.0007 1.26363e-08 0 1.27303e-08 0 1.27333e-08 0.0007 1.27363e-08 0 1.30303e-08 0 1.30333e-08 0.0007 1.30363e-08 0 1.31303e-08 0 1.31333e-08 0.0007 1.31363e-08 0 1.34303e-08 0 1.34333e-08 0.0007 1.34363e-08 0 1.35303e-08 0 1.35333e-08 0.0007 1.35363e-08 0 1.38303e-08 0 1.38333e-08 0.0007 1.38363e-08 0 1.39303e-08 0 1.39333e-08 0.0007 1.39363e-08 0 1.42303e-08 0 1.42333e-08 0.0007 1.42363e-08 0 1.43303e-08 0 1.43333e-08 0.0007 1.43363e-08 0 1.46303e-08 0 1.46333e-08 0.0007 1.46363e-08 0 1.47303e-08 0 1.47333e-08 0.0007 1.47363e-08 0 1.50303e-08 0 1.50333e-08 0.0007 1.50363e-08 0 1.51303e-08 0 1.51333e-08 0.0007 1.51363e-08 0 1.54303e-08 0 1.54333e-08 0.0007 1.54363e-08 0 1.55303e-08 0 1.55333e-08 0.0007 1.55363e-08 0 1.58303e-08 0 1.58333e-08 0.0007 1.58363e-08 0 1.59303e-08 0 1.59333e-08 0.0007 1.59363e-08 0 1.62303e-08 0 1.62333e-08 0.0007 1.62363e-08 0 1.63303e-08 0 1.63333e-08 0.0007 1.63363e-08 0 1.66303e-08 0 1.66333e-08 0.0007 1.66363e-08 0 1.67303e-08 0 1.67333e-08 0.0007 1.67363e-08 0 1.70303e-08 0 1.70333e-08 0.0007 1.70363e-08 0 1.71303e-08 0 1.71333e-08 0.0007 1.71363e-08 0 1.74303e-08 0 1.74333e-08 0.0007 1.74363e-08 0 1.75303e-08 0 1.75333e-08 0.0007 1.75363e-08 0 1.78303e-08 0 1.78333e-08 0.0007 1.78363e-08 0 1.79303e-08 0 1.79333e-08 0.0007 1.79363e-08 0 1.82303e-08 0 1.82333e-08 0.0007 1.82363e-08 0 1.83303e-08 0 1.83333e-08 0.0007 1.83363e-08 0 1.86303e-08 0 1.86333e-08 0.0007 1.86363e-08 0 1.87303e-08 0 1.87333e-08 0.0007 1.87363e-08 0 1.90303e-08 0 1.90333e-08 0.0007 1.90363e-08 0 1.91303e-08 0 1.91333e-08 0.0007 1.91363e-08 0 1.94303e-08 0 1.94333e-08 0.0007 1.94363e-08 0 1.95303e-08 0 1.95333e-08 0.0007 1.95363e-08 0 1.98303e-08 0 1.98333e-08 0.0007 1.98363e-08 0 1.99303e-08 0 1.99333e-08 0.0007 1.99363e-08 0 2.02303e-08 0 2.02333e-08 0.0007 2.02363e-08 0 2.03303e-08 0 2.03333e-08 0.0007 2.03363e-08 0 2.06303e-08 0 2.06333e-08 0.0007 2.06363e-08 0 2.07303e-08 0 2.07333e-08 0.0007 2.07363e-08 0 2.10303e-08 0 2.10333e-08 0.0007 2.10363e-08 0 2.11303e-08 0 2.11333e-08 0.0007 2.11363e-08 0 2.14303e-08 0 2.14333e-08 0.0007 2.14363e-08 0 2.15303e-08 0 2.15333e-08 0.0007 2.15363e-08 0 2.18303e-08 0 2.18333e-08 0.0007 2.18363e-08 0 2.19303e-08 0 2.19333e-08 0.0007 2.19363e-08 0 2.22303e-08 0 2.22333e-08 0.0007 2.22363e-08 0 2.23303e-08 0 2.23333e-08 0.0007 2.23363e-08 0 2.26303e-08 0 2.26333e-08 0.0007 2.26363e-08 0 2.27303e-08 0 2.27333e-08 0.0007 2.27363e-08 0 2.30303e-08 0 2.30333e-08 0.0007 2.30363e-08 0 2.31303e-08 0 2.31333e-08 0.0007 2.31363e-08 0 2.34303e-08 0 2.34333e-08 0.0007 2.34363e-08 0 2.35303e-08 0 2.35333e-08 0.0007 2.35363e-08 0 2.38303e-08 0 2.38333e-08 0.0007 2.38363e-08 0 2.39303e-08 0 2.39333e-08 0.0007 2.39363e-08 0 2.42303e-08 0 2.42333e-08 0.0007 2.42363e-08 0 2.43303e-08 0 2.43333e-08 0.0007 2.43363e-08 0 2.46303e-08 0 2.46333e-08 0.0007 2.46363e-08 0 2.47303e-08 0 2.47333e-08 0.0007 2.47363e-08 0 2.50303e-08 0 2.50333e-08 0.0007 2.50363e-08 0 2.51303e-08 0 2.51333e-08 0.0007 2.51363e-08 0 2.54303e-08 0 2.54333e-08 0.0007 2.54363e-08 0 2.55303e-08 0 2.55333e-08 0.0007 2.55363e-08 0)
L_DFF|1 A _DFF|A1  2.067833848e-12
L_DFF|2 _DFF|A1 _DFF|A2  4.135667696e-12
L_DFF|3 _DFF|A3 _DFF|A4  8.271335392e-12
L_DFF|T CLK _DFF|T1  2.067833848e-12
L_DFF|4 _DFF|T1 _DFF|T2  4.135667696e-12
L_DFF|5 _DFF|A4 _DFF|Q1  4.135667696e-12
L_DFF|6 _DFF|Q1 DFF_A  2.067833848e-12
L_NOT|1 B _NOT|A1  2.067833848e-12
L_NOT|2 _NOT|A1 _NOT|A2  4.135667696e-12
L_NOT|3 _NOT|A2 _NOT|A3  4.135667696e-12
L_NOT|4 CLK _NOT|T1  2.067833848e-12
L_NOT|5 _NOT|T1 _NOT|T2  1e-12
L_NOT|7 _NOT|T2 _NOT|CW1  2e-12
L_NOT|8 _NOT|CW1 _NOT|CW2  1e-12
L_NOT|9 _NOT|CW2 _NOT|A4  8.271335392e-12
L_NOT|10 _NOT|A4 _NOT|CW3  1e-12
L_NOT|6 _NOT|T2 _NOT|CCW  4.135667696e-12
L_NOT|11 _NOT|Q2 _NOT|Q1  4.135667696e-12
L_NOT|12 _NOT|Q1 NOT_B  2.067833848e-12
L_NOT|RD _NOT|CW1 _NOT|112  2e-12
R_NOT|D _NOT|112 0  4
L_MERGE|A1 DFF_A _MERGE|A1  2.067833848e-12
L_MERGE|A2 _MERGE|A1 _MERGE|A2  4.135667696e-12
L_MERGE|A3 _MERGE|A3 _MERGE|Q3  1.2e-12
L_MERGE|B1 NOT_B _MERGE|B1  2.067833848e-12
L_MERGE|B2 _MERGE|B1 _MERGE|B2  4.135667696e-12
L_MERGE|B3 _MERGE|B3 _MERGE|Q3  1.2e-12
L_MERGE|Q3 _MERGE|Q3 _MERGE|Q2  4.135667696e-12
L_MERGE|Q2 _MERGE|Q2 _MERGE|Q1  4.135667696e-12
L_MERGE|Q1 _MERGE|Q1 Q  2.067833848e-12
L_DFF|I_1|B _DFF|A1 _DFF|I_1|MID  2e-12
I_DFF|I_1|B 0 _DFF|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF|I_3|B _DFF|A3 _DFF|I_3|MID  2e-12
I_DFF|I_3|B 0 _DFF|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF|I_T|B _DFF|T1 _DFF|I_T|MID  2e-12
I_DFF|I_T|B 0 _DFF|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF|I_6|B _DFF|Q1 _DFF|I_6|MID  2e-12
I_DFF|I_6|B 0 _DFF|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF|1|1 _DFF|A1 _DFF|1|MID_SERIES JJMIT AREA=2.5
L_DFF|1|P _DFF|1|MID_SERIES 0  2e-13
R_DFF|1|B _DFF|A1 _DFF|1|MID_SHUNT  2.7439617672
L_DFF|1|RB _DFF|1|MID_SHUNT 0  1.550338398468e-12
B_DFF|23|1 _DFF|A2 _DFF|A3 JJMIT AREA=1.7857142857142858
R_DFF|23|B _DFF|A2 _DFF|23|MID_SHUNT  3.84154647408
L_DFF|23|RB _DFF|23|MID_SHUNT _DFF|A3  2.1704737578552e-12
B_DFF|3|1 _DFF|A3 _DFF|3|MID_SERIES JJMIT AREA=2.5
L_DFF|3|P _DFF|3|MID_SERIES 0  2e-13
R_DFF|3|B _DFF|A3 _DFF|3|MID_SHUNT  2.7439617672
L_DFF|3|RB _DFF|3|MID_SHUNT 0  1.550338398468e-12
B_DFF|4|1 _DFF|A4 _DFF|4|MID_SERIES JJMIT AREA=2.5
L_DFF|4|P _DFF|4|MID_SERIES 0  2e-13
R_DFF|4|B _DFF|A4 _DFF|4|MID_SHUNT  2.7439617672
L_DFF|4|RB _DFF|4|MID_SHUNT 0  1.550338398468e-12
B_DFF|T|1 _DFF|T1 _DFF|T|MID_SERIES JJMIT AREA=2.5
L_DFF|T|P _DFF|T|MID_SERIES 0  2e-13
R_DFF|T|B _DFF|T1 _DFF|T|MID_SHUNT  2.7439617672
L_DFF|T|RB _DFF|T|MID_SHUNT 0  1.550338398468e-12
B_DFF|45|1 _DFF|T2 _DFF|A4 JJMIT AREA=1.7857142857142858
R_DFF|45|B _DFF|T2 _DFF|45|MID_SHUNT  3.84154647408
L_DFF|45|RB _DFF|45|MID_SHUNT _DFF|A4  2.1704737578552e-12
B_DFF|6|1 _DFF|Q1 _DFF|6|MID_SERIES JJMIT AREA=2.5
L_DFF|6|P _DFF|6|MID_SERIES 0  2e-13
R_DFF|6|B _DFF|Q1 _DFF|6|MID_SHUNT  2.7439617672
L_DFF|6|RB _DFF|6|MID_SHUNT 0  1.550338398468e-12
B_NOT|1|1 _NOT|A1 _NOT|1|MID_SERIES JJMIT AREA=2.5
L_NOT|1|P _NOT|1|MID_SERIES 0  2e-13
R_NOT|1|B _NOT|A1 _NOT|1|MID_SHUNT  2.7439617672
L_NOT|1|RB _NOT|1|MID_SHUNT 0  1.550338398468e-12
B_NOT|2|1 _NOT|A2 _NOT|2|B_JCT JJMIT AREA=1.7857142857142858
R_NOT|2|B _NOT|A2 _NOT|2|MID_SHUNT  3.84154647408
L_NOT|2|RB _NOT|2|MID_SHUNT _NOT|2|B_JCT  2.1704737578552e-12
L_NOT|2|P_SERIES _NOT|2|B_JCT 0  2e-13
B_NOT|3|1 _NOT|A3 _NOT|A4 JJMIT AREA=1.7857142857142858
R_NOT|3|B _NOT|A3 _NOT|3|MID_SHUNT  3.84154647408
L_NOT|3|RB _NOT|3|MID_SHUNT _NOT|A4  2.1704737578552e-12
B_NOT|4|1 _NOT|T1 _NOT|4|MID_SERIES JJMIT AREA=2.5
L_NOT|4|P _NOT|4|MID_SERIES 0  2e-13
R_NOT|4|B _NOT|T1 _NOT|4|MID_SHUNT  2.7439617672
L_NOT|4|RB _NOT|4|MID_SHUNT 0  1.550338398468e-12
B_NOT|6|1 _NOT|CW2 _NOT|6|MID_SERIES JJMIT AREA=2.5
L_NOT|6|P _NOT|6|MID_SERIES 0  2e-13
R_NOT|6|B _NOT|CW2 _NOT|6|MID_SHUNT  2.7439617672
L_NOT|6|RB _NOT|6|MID_SHUNT 0  1.550338398468e-12
B_NOT|7|1 _NOT|CW3 _NOT|Q2 JJMIT AREA=1.7857142857142858
R_NOT|7|B _NOT|CW3 _NOT|7|MID_SHUNT  3.84154647408
L_NOT|7|RB _NOT|7|MID_SHUNT _NOT|Q2  2.1704737578552e-12
B_NOT|5|1 _NOT|CCW _NOT|Q2 JJMIT AREA=1.7857142857142858
R_NOT|5|B _NOT|CCW _NOT|5|MID_SHUNT  3.84154647408
L_NOT|5|RB _NOT|5|MID_SHUNT _NOT|Q2  2.1704737578552e-12
B_NOT|8|1 _NOT|Q2 _NOT|8|MID_SERIES JJMIT AREA=2.5
L_NOT|8|P _NOT|8|MID_SERIES 0  2e-13
R_NOT|8|B _NOT|Q2 _NOT|8|MID_SHUNT  2.7439617672
L_NOT|8|RB _NOT|8|MID_SHUNT 0  1.550338398468e-12
B_NOT|9|1 _NOT|Q1 _NOT|9|MID_SERIES JJMIT AREA=2.5
L_NOT|9|P _NOT|9|MID_SERIES 0  2e-13
R_NOT|9|B _NOT|Q1 _NOT|9|MID_SHUNT  2.7439617672
L_NOT|9|RB _NOT|9|MID_SHUNT 0  1.550338398468e-12
L_NOT|I_A1|B _NOT|A1 _NOT|I_A1|MID  2e-12
I_NOT|I_A1|B 0 _NOT|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_NOT|I_A2|B _NOT|A2 _NOT|I_A2|MID  2e-12
I_NOT|I_A2|B 0 _NOT|I_A2|MID  PWL(0 0 5e-12 0.000125)
L_NOT|I_A4|B _NOT|A4 _NOT|I_A4|MID  2e-12
I_NOT|I_A4|B 0 _NOT|I_A4|MID  PWL(0 0 5e-12 0.000175)
L_NOT|I_T1|B _NOT|T1 _NOT|I_T1|MID  2e-12
I_NOT|I_T1|B 0 _NOT|I_T1|MID  PWL(0 0 5e-12 0.000175)
L_NOT|I_Q1|B _NOT|Q1 _NOT|I_Q1|MID  2e-12
I_NOT|I_Q1|B 0 _NOT|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_MERGE|I_A1|B _MERGE|A1 _MERGE|I_A1|MID  2e-12
I_MERGE|I_A1|B 0 _MERGE|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_MERGE|I_B1|B _MERGE|B1 _MERGE|I_B1|MID  2e-12
I_MERGE|I_B1|B 0 _MERGE|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_MERGE|I_Q3|B _MERGE|Q3 _MERGE|I_Q3|MID  2e-12
I_MERGE|I_Q3|B 0 _MERGE|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_MERGE|I_Q2|B _MERGE|Q2 _MERGE|I_Q2|MID  2e-12
I_MERGE|I_Q2|B 0 _MERGE|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_MERGE|I_Q1|B _MERGE|Q1 _MERGE|I_Q1|MID  2e-12
I_MERGE|I_Q1|B 0 _MERGE|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_MERGE|A1|1 _MERGE|A1 _MERGE|A1|MID_SERIES JJMIT AREA=2.5
L_MERGE|A1|P _MERGE|A1|MID_SERIES 0  2e-13
R_MERGE|A1|B _MERGE|A1 _MERGE|A1|MID_SHUNT  2.7439617672
L_MERGE|A1|RB _MERGE|A1|MID_SHUNT 0  1.550338398468e-12
B_MERGE|A2|1 _MERGE|A2 _MERGE|A2|MID_SERIES JJMIT AREA=2.5
L_MERGE|A2|P _MERGE|A2|MID_SERIES 0  2e-13
R_MERGE|A2|B _MERGE|A2 _MERGE|A2|MID_SHUNT  2.7439617672
L_MERGE|A2|RB _MERGE|A2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|A12|1 _MERGE|A2 _MERGE|A3 JJMIT AREA=1.7857142857142858
R_MERGE|A12|B _MERGE|A2 _MERGE|A12|MID_SHUNT  3.84154647408
L_MERGE|A12|RB _MERGE|A12|MID_SHUNT _MERGE|A3  2.1704737578552e-12
B_MERGE|B1|1 _MERGE|B1 _MERGE|B1|MID_SERIES JJMIT AREA=2.5
L_MERGE|B1|P _MERGE|B1|MID_SERIES 0  2e-13
R_MERGE|B1|B _MERGE|B1 _MERGE|B1|MID_SHUNT  2.7439617672
L_MERGE|B1|RB _MERGE|B1|MID_SHUNT 0  1.550338398468e-12
B_MERGE|B2|1 _MERGE|B2 _MERGE|B2|MID_SERIES JJMIT AREA=2.5
L_MERGE|B2|P _MERGE|B2|MID_SERIES 0  2e-13
R_MERGE|B2|B _MERGE|B2 _MERGE|B2|MID_SHUNT  2.7439617672
L_MERGE|B2|RB _MERGE|B2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|B12|1 _MERGE|B2 _MERGE|B3 JJMIT AREA=1.7857142857142858
R_MERGE|B12|B _MERGE|B2 _MERGE|B12|MID_SHUNT  3.84154647408
L_MERGE|B12|RB _MERGE|B12|MID_SHUNT _MERGE|B3  2.1704737578552e-12
B_MERGE|Q2|1 _MERGE|Q2 _MERGE|Q2|MID_SERIES JJMIT AREA=2.5
L_MERGE|Q2|P _MERGE|Q2|MID_SERIES 0  2e-13
R_MERGE|Q2|B _MERGE|Q2 _MERGE|Q2|MID_SHUNT  2.7439617672
L_MERGE|Q2|RB _MERGE|Q2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|Q1|1 _MERGE|Q1 _MERGE|Q1|MID_SERIES JJMIT AREA=2.5
L_MERGE|Q1|P _MERGE|Q1|MID_SERIES 0  2e-13
R_MERGE|Q1|B _MERGE|Q1 _MERGE|Q1|MID_SHUNT  2.7439617672
L_MERGE|Q1|RB _MERGE|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI ROUT
.print DEVI IT1|T
.print DEVI IDATA_A1|A
.print DEVI IDATA_B1|B
.print DEVI L_DFF|1
.print DEVI L_DFF|2
.print DEVI L_DFF|3
.print DEVI L_DFF|T
.print DEVI L_DFF|4
.print DEVI L_DFF|5
.print DEVI L_DFF|6
.print DEVI L_NOT|1
.print DEVI L_NOT|2
.print DEVI L_NOT|3
.print DEVI L_NOT|4
.print DEVI L_NOT|5
.print DEVI L_NOT|7
.print DEVI L_NOT|8
.print DEVI L_NOT|9
.print DEVI L_NOT|10
.print DEVI L_NOT|6
.print DEVI L_NOT|11
.print DEVI L_NOT|12
.print DEVI L_NOT|RD
.print DEVI R_NOT|D
.print DEVI L_MERGE|A1
.print DEVI L_MERGE|A2
.print DEVI L_MERGE|A3
.print DEVI L_MERGE|B1
.print DEVI L_MERGE|B2
.print DEVI L_MERGE|B3
.print DEVI L_MERGE|Q3
.print DEVI L_MERGE|Q2
.print DEVI L_MERGE|Q1
.print V _NOT|A1
.print V _NOT|A3
.print V _NOT|A2
.print V _MERGE|B1
.print V A
.print V _MERGE|B2
.print V _NOT|T1
.print V _DFF|A4
.print V _DFF|Q1
.print V _MERGE|Q3
.print V _NOT|CCW
.print V _DFF|A1
.print V _DFF|T2
.print V _NOT|T2
.print V _MERGE|Q1
.print V _MERGE|Q2
.print V _MERGE|A3
.print V CLK
.print V _MERGE|A1
.print V _NOT|CW3
.print V DFF_A
.print V _MERGE|B3
.print V _DFF|A2
.print V Q
.print V NOT_B
.print V _NOT|CW1
.print V _MERGE|A2
.print V _DFF|A3
.print V _NOT|112
.print V _NOT|CW2
.print V _DFF|T1
.print V B
.print V _NOT|Q2
.print V _NOT|Q1
.print V _NOT|A4
.print DEVP B_DFF|1|1
.print DEVP B_DFF|23|1
.print DEVP B_DFF|3|1
.print DEVP B_DFF|4|1
.print DEVP B_DFF|T|1
.print DEVP B_DFF|45|1
.print DEVP B_DFF|6|1
.print DEVP B_NOT|1|1
.print DEVP B_NOT|2|1
.print DEVP B_NOT|3|1
.print DEVP B_NOT|4|1
.print DEVP B_NOT|6|1
.print DEVP B_NOT|7|1
.print DEVP B_NOT|5|1
.print DEVP B_NOT|8|1
.print DEVP B_NOT|9|1
.print DEVP B_MERGE|A1|1
.print DEVP B_MERGE|A2|1
.print DEVP B_MERGE|A12|1
.print DEVP B_MERGE|B1|1
.print DEVP B_MERGE|B2|1
.print DEVP B_MERGE|B12|1
.print DEVP B_MERGE|Q2|1
.print DEVP B_MERGE|Q1|1
