*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM DCBIAS=1
.PARAM TCLOCK=1.8e-10
.PARAM OS=4.5e-12
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 52000E-12/200*180
R_S0 S0 0  1
R_S1 S1 0  1
R_S2 S2 0  1
R_S3 S3 0  1
R_S4 S4 0  1
IA0|A 0 A0  PWL(0 0 2.103e-10 0 2.133e-10 0.0007 2.163e-10 0 5.703e-10 0 5.733e-10 0.0007 5.763e-10 0 9.303e-10 0 9.333e-10 0.0007 9.363e-10 0 1.2903e-09 0 1.2933e-09 0.0007 1.2963e-09 0 1.6503e-09 0 1.6533e-09 0.0007 1.6563e-09 0 2.0103e-09 0 2.0133e-09 0.0007 2.0163e-09 0 2.3703e-09 0 2.3733e-09 0.0007 2.3763e-09 0 2.7303e-09 0 2.7333e-09 0.0007 2.7363e-09 0 3.0903e-09 0 3.0933e-09 0.0007 3.0963e-09 0 3.4503e-09 0 3.4533e-09 0.0007 3.4563e-09 0 3.8103e-09 0 3.8133e-09 0.0007 3.8163e-09 0 4.1703e-09 0 4.1733e-09 0.0007 4.1763e-09 0 4.5303e-09 0 4.5333e-09 0.0007 4.5363e-09 0 4.8903e-09 0 4.8933e-09 0.0007 4.8963e-09 0 5.2503e-09 0 5.2533e-09 0.0007 5.2563e-09 0 5.6103e-09 0 5.6133e-09 0.0007 5.6163e-09 0 5.9703e-09 0 5.9733e-09 0.0007 5.9763e-09 0 6.3303e-09 0 6.3333e-09 0.0007 6.3363e-09 0 6.6903e-09 0 6.6933e-09 0.0007 6.6963e-09 0 7.0503e-09 0 7.0533e-09 0.0007 7.0563e-09 0 7.4103e-09 0 7.4133e-09 0.0007 7.4163e-09 0 7.7703e-09 0 7.7733e-09 0.0007 7.7763e-09 0 8.1303e-09 0 8.1333e-09 0.0007 8.1363e-09 0 8.4903e-09 0 8.4933e-09 0.0007 8.4963e-09 0 8.8503e-09 0 8.8533e-09 0.0007 8.8563e-09 0 9.2103e-09 0 9.2133e-09 0.0007 9.2163e-09 0 9.5703e-09 0 9.5733e-09 0.0007 9.5763e-09 0 9.9303e-09 0 9.9333e-09 0.0007 9.9363e-09 0 1.02903e-08 0 1.02933e-08 0.0007 1.02963e-08 0 1.06503e-08 0 1.06533e-08 0.0007 1.06563e-08 0 1.10103e-08 0 1.10133e-08 0.0007 1.10163e-08 0 1.13703e-08 0 1.13733e-08 0.0007 1.13763e-08 0 1.17303e-08 0 1.17333e-08 0.0007 1.17363e-08 0 1.20903e-08 0 1.20933e-08 0.0007 1.20963e-08 0 1.24503e-08 0 1.24533e-08 0.0007 1.24563e-08 0 1.28103e-08 0 1.28133e-08 0.0007 1.28163e-08 0 1.31703e-08 0 1.31733e-08 0.0007 1.31763e-08 0 1.35303e-08 0 1.35333e-08 0.0007 1.35363e-08 0 1.38903e-08 0 1.38933e-08 0.0007 1.38963e-08 0 1.42503e-08 0 1.42533e-08 0.0007 1.42563e-08 0 1.46103e-08 0 1.46133e-08 0.0007 1.46163e-08 0 1.49703e-08 0 1.49733e-08 0.0007 1.49763e-08 0 1.53303e-08 0 1.53333e-08 0.0007 1.53363e-08 0 1.56903e-08 0 1.56933e-08 0.0007 1.56963e-08 0 1.60503e-08 0 1.60533e-08 0.0007 1.60563e-08 0 1.64103e-08 0 1.64133e-08 0.0007 1.64163e-08 0 1.67703e-08 0 1.67733e-08 0.0007 1.67763e-08 0 1.71303e-08 0 1.71333e-08 0.0007 1.71363e-08 0 1.74903e-08 0 1.74933e-08 0.0007 1.74963e-08 0 1.78503e-08 0 1.78533e-08 0.0007 1.78563e-08 0 1.82103e-08 0 1.82133e-08 0.0007 1.82163e-08 0 1.85703e-08 0 1.85733e-08 0.0007 1.85763e-08 0 1.89303e-08 0 1.89333e-08 0.0007 1.89363e-08 0 1.92903e-08 0 1.92933e-08 0.0007 1.92963e-08 0 1.96503e-08 0 1.96533e-08 0.0007 1.96563e-08 0 2.00103e-08 0 2.00133e-08 0.0007 2.00163e-08 0 2.03703e-08 0 2.03733e-08 0.0007 2.03763e-08 0 2.07303e-08 0 2.07333e-08 0.0007 2.07363e-08 0 2.10903e-08 0 2.10933e-08 0.0007 2.10963e-08 0 2.14503e-08 0 2.14533e-08 0.0007 2.14563e-08 0 2.18103e-08 0 2.18133e-08 0.0007 2.18163e-08 0 2.21703e-08 0 2.21733e-08 0.0007 2.21763e-08 0 2.25303e-08 0 2.25333e-08 0.0007 2.25363e-08 0 2.28903e-08 0 2.28933e-08 0.0007 2.28963e-08 0 2.32503e-08 0 2.32533e-08 0.0007 2.32563e-08 0 2.36103e-08 0 2.36133e-08 0.0007 2.36163e-08 0 2.39703e-08 0 2.39733e-08 0.0007 2.39763e-08 0 2.43303e-08 0 2.43333e-08 0.0007 2.43363e-08 0 2.46903e-08 0 2.46933e-08 0.0007 2.46963e-08 0 2.50503e-08 0 2.50533e-08 0.0007 2.50563e-08 0 2.54103e-08 0 2.54133e-08 0.0007 2.54163e-08 0 2.57703e-08 0 2.57733e-08 0.0007 2.57763e-08 0 2.61303e-08 0 2.61333e-08 0.0007 2.61363e-08 0 2.64903e-08 0 2.64933e-08 0.0007 2.64963e-08 0 2.68503e-08 0 2.68533e-08 0.0007 2.68563e-08 0 2.72103e-08 0 2.72133e-08 0.0007 2.72163e-08 0 2.75703e-08 0 2.75733e-08 0.0007 2.75763e-08 0 2.79303e-08 0 2.79333e-08 0.0007 2.79363e-08 0 2.82903e-08 0 2.82933e-08 0.0007 2.82963e-08 0 2.86503e-08 0 2.86533e-08 0.0007 2.86563e-08 0 2.90103e-08 0 2.90133e-08 0.0007 2.90163e-08 0 2.93703e-08 0 2.93733e-08 0.0007 2.93763e-08 0 2.97303e-08 0 2.97333e-08 0.0007 2.97363e-08 0 3.00903e-08 0 3.00933e-08 0.0007 3.00963e-08 0 3.04503e-08 0 3.04533e-08 0.0007 3.04563e-08 0 3.08103e-08 0 3.08133e-08 0.0007 3.08163e-08 0 3.11703e-08 0 3.11733e-08 0.0007 3.11763e-08 0 3.15303e-08 0 3.15333e-08 0.0007 3.15363e-08 0 3.18903e-08 0 3.18933e-08 0.0007 3.18963e-08 0 3.22503e-08 0 3.22533e-08 0.0007 3.22563e-08 0 3.26103e-08 0 3.26133e-08 0.0007 3.26163e-08 0 3.29703e-08 0 3.29733e-08 0.0007 3.29763e-08 0 3.33303e-08 0 3.33333e-08 0.0007 3.33363e-08 0 3.36903e-08 0 3.36933e-08 0.0007 3.36963e-08 0 3.40503e-08 0 3.40533e-08 0.0007 3.40563e-08 0 3.44103e-08 0 3.44133e-08 0.0007 3.44163e-08 0 3.47703e-08 0 3.47733e-08 0.0007 3.47763e-08 0 3.51303e-08 0 3.51333e-08 0.0007 3.51363e-08 0 3.54903e-08 0 3.54933e-08 0.0007 3.54963e-08 0 3.58503e-08 0 3.58533e-08 0.0007 3.58563e-08 0 3.62103e-08 0 3.62133e-08 0.0007 3.62163e-08 0 3.65703e-08 0 3.65733e-08 0.0007 3.65763e-08 0 3.69303e-08 0 3.69333e-08 0.0007 3.69363e-08 0 3.72903e-08 0 3.72933e-08 0.0007 3.72963e-08 0 3.76503e-08 0 3.76533e-08 0.0007 3.76563e-08 0 3.80103e-08 0 3.80133e-08 0.0007 3.80163e-08 0 3.83703e-08 0 3.83733e-08 0.0007 3.83763e-08 0 3.87303e-08 0 3.87333e-08 0.0007 3.87363e-08 0 3.90903e-08 0 3.90933e-08 0.0007 3.90963e-08 0 3.94503e-08 0 3.94533e-08 0.0007 3.94563e-08 0 3.98103e-08 0 3.98133e-08 0.0007 3.98163e-08 0 4.01703e-08 0 4.01733e-08 0.0007 4.01763e-08 0 4.05303e-08 0 4.05333e-08 0.0007 4.05363e-08 0 4.08903e-08 0 4.08933e-08 0.0007 4.08963e-08 0 4.12503e-08 0 4.12533e-08 0.0007 4.12563e-08 0 4.16103e-08 0 4.16133e-08 0.0007 4.16163e-08 0 4.19703e-08 0 4.19733e-08 0.0007 4.19763e-08 0 4.23303e-08 0 4.23333e-08 0.0007 4.23363e-08 0 4.26903e-08 0 4.26933e-08 0.0007 4.26963e-08 0 4.30503e-08 0 4.30533e-08 0.0007 4.30563e-08 0 4.34103e-08 0 4.34133e-08 0.0007 4.34163e-08 0 4.37703e-08 0 4.37733e-08 0.0007 4.37763e-08 0 4.41303e-08 0 4.41333e-08 0.0007 4.41363e-08 0 4.44903e-08 0 4.44933e-08 0.0007 4.44963e-08 0 4.48503e-08 0 4.48533e-08 0.0007 4.48563e-08 0 4.52103e-08 0 4.52133e-08 0.0007 4.52163e-08 0 4.55703e-08 0 4.55733e-08 0.0007 4.55763e-08 0 4.59303e-08 0 4.59333e-08 0.0007 4.59363e-08 0)
IB0|B 0 B0  PWL(0 0 4.047e-10 0 4.077e-10 0.0007 4.107e-10 0 5.847e-10 0 5.877e-10 0.0007 5.907e-10 0 1.1247e-09 0 1.1277e-09 0.0007 1.1307e-09 0 1.3047e-09 0 1.3077e-09 0.0007 1.3107e-09 0 1.8447e-09 0 1.8477e-09 0.0007 1.8507e-09 0 2.0247e-09 0 2.0277e-09 0.0007 2.0307e-09 0 2.5647e-09 0 2.5677e-09 0.0007 2.5707e-09 0 2.7447e-09 0 2.7477e-09 0.0007 2.7507e-09 0 3.2847e-09 0 3.2877e-09 0.0007 3.2907e-09 0 3.4647e-09 0 3.4677e-09 0.0007 3.4707e-09 0 4.0047e-09 0 4.0077e-09 0.0007 4.0107e-09 0 4.1847e-09 0 4.1877e-09 0.0007 4.1907e-09 0 4.7247e-09 0 4.7277e-09 0.0007 4.7307e-09 0 4.9047e-09 0 4.9077e-09 0.0007 4.9107e-09 0 5.4447e-09 0 5.4477e-09 0.0007 5.4507e-09 0 5.6247e-09 0 5.6277e-09 0.0007 5.6307e-09 0 6.1647e-09 0 6.1677e-09 0.0007 6.1707e-09 0 6.3447e-09 0 6.3477e-09 0.0007 6.3507e-09 0 6.8847e-09 0 6.8877e-09 0.0007 6.8907e-09 0 7.0647e-09 0 7.0677e-09 0.0007 7.0707e-09 0 7.6047e-09 0 7.6077e-09 0.0007 7.6107e-09 0 7.7847e-09 0 7.7877e-09 0.0007 7.7907e-09 0 8.3247e-09 0 8.3277e-09 0.0007 8.3307e-09 0 8.5047e-09 0 8.5077e-09 0.0007 8.5107e-09 0 9.0447e-09 0 9.0477e-09 0.0007 9.0507e-09 0 9.2247e-09 0 9.2277e-09 0.0007 9.2307e-09 0 9.7647e-09 0 9.7677e-09 0.0007 9.7707e-09 0 9.9447e-09 0 9.9477e-09 0.0007 9.9507e-09 0 1.04847e-08 0 1.04877e-08 0.0007 1.04907e-08 0 1.06647e-08 0 1.06677e-08 0.0007 1.06707e-08 0 1.12047e-08 0 1.12077e-08 0.0007 1.12107e-08 0 1.13847e-08 0 1.13877e-08 0.0007 1.13907e-08 0 1.19247e-08 0 1.19277e-08 0.0007 1.19307e-08 0 1.21047e-08 0 1.21077e-08 0.0007 1.21107e-08 0 1.26447e-08 0 1.26477e-08 0.0007 1.26507e-08 0 1.28247e-08 0 1.28277e-08 0.0007 1.28307e-08 0 1.33647e-08 0 1.33677e-08 0.0007 1.33707e-08 0 1.35447e-08 0 1.35477e-08 0.0007 1.35507e-08 0 1.40847e-08 0 1.40877e-08 0.0007 1.40907e-08 0 1.42647e-08 0 1.42677e-08 0.0007 1.42707e-08 0 1.48047e-08 0 1.48077e-08 0.0007 1.48107e-08 0 1.49847e-08 0 1.49877e-08 0.0007 1.49907e-08 0 1.55247e-08 0 1.55277e-08 0.0007 1.55307e-08 0 1.57047e-08 0 1.57077e-08 0.0007 1.57107e-08 0 1.62447e-08 0 1.62477e-08 0.0007 1.62507e-08 0 1.64247e-08 0 1.64277e-08 0.0007 1.64307e-08 0 1.69647e-08 0 1.69677e-08 0.0007 1.69707e-08 0 1.71447e-08 0 1.71477e-08 0.0007 1.71507e-08 0 1.76847e-08 0 1.76877e-08 0.0007 1.76907e-08 0 1.78647e-08 0 1.78677e-08 0.0007 1.78707e-08 0 1.84047e-08 0 1.84077e-08 0.0007 1.84107e-08 0 1.85847e-08 0 1.85877e-08 0.0007 1.85907e-08 0 1.91247e-08 0 1.91277e-08 0.0007 1.91307e-08 0 1.93047e-08 0 1.93077e-08 0.0007 1.93107e-08 0 1.98447e-08 0 1.98477e-08 0.0007 1.98507e-08 0 2.00247e-08 0 2.00277e-08 0.0007 2.00307e-08 0 2.05647e-08 0 2.05677e-08 0.0007 2.05707e-08 0 2.07447e-08 0 2.07477e-08 0.0007 2.07507e-08 0 2.12847e-08 0 2.12877e-08 0.0007 2.12907e-08 0 2.14647e-08 0 2.14677e-08 0.0007 2.14707e-08 0 2.20047e-08 0 2.20077e-08 0.0007 2.20107e-08 0 2.21847e-08 0 2.21877e-08 0.0007 2.21907e-08 0 2.27247e-08 0 2.27277e-08 0.0007 2.27307e-08 0 2.29047e-08 0 2.29077e-08 0.0007 2.29107e-08 0 2.34447e-08 0 2.34477e-08 0.0007 2.34507e-08 0 2.36247e-08 0 2.36277e-08 0.0007 2.36307e-08 0 2.41647e-08 0 2.41677e-08 0.0007 2.41707e-08 0 2.43447e-08 0 2.43477e-08 0.0007 2.43507e-08 0 2.48847e-08 0 2.48877e-08 0.0007 2.48907e-08 0 2.50647e-08 0 2.50677e-08 0.0007 2.50707e-08 0 2.56047e-08 0 2.56077e-08 0.0007 2.56107e-08 0 2.57847e-08 0 2.57877e-08 0.0007 2.57907e-08 0 2.63247e-08 0 2.63277e-08 0.0007 2.63307e-08 0 2.65047e-08 0 2.65077e-08 0.0007 2.65107e-08 0 2.70447e-08 0 2.70477e-08 0.0007 2.70507e-08 0 2.72247e-08 0 2.72277e-08 0.0007 2.72307e-08 0 2.77647e-08 0 2.77677e-08 0.0007 2.77707e-08 0 2.79447e-08 0 2.79477e-08 0.0007 2.79507e-08 0 2.84847e-08 0 2.84877e-08 0.0007 2.84907e-08 0 2.86647e-08 0 2.86677e-08 0.0007 2.86707e-08 0 2.92047e-08 0 2.92077e-08 0.0007 2.92107e-08 0 2.93847e-08 0 2.93877e-08 0.0007 2.93907e-08 0 2.99247e-08 0 2.99277e-08 0.0007 2.99307e-08 0 3.01047e-08 0 3.01077e-08 0.0007 3.01107e-08 0 3.06447e-08 0 3.06477e-08 0.0007 3.06507e-08 0 3.08247e-08 0 3.08277e-08 0.0007 3.08307e-08 0 3.13647e-08 0 3.13677e-08 0.0007 3.13707e-08 0 3.15447e-08 0 3.15477e-08 0.0007 3.15507e-08 0 3.20847e-08 0 3.20877e-08 0.0007 3.20907e-08 0 3.22647e-08 0 3.22677e-08 0.0007 3.22707e-08 0 3.28047e-08 0 3.28077e-08 0.0007 3.28107e-08 0 3.29847e-08 0 3.29877e-08 0.0007 3.29907e-08 0 3.35247e-08 0 3.35277e-08 0.0007 3.35307e-08 0 3.37047e-08 0 3.37077e-08 0.0007 3.37107e-08 0 3.42447e-08 0 3.42477e-08 0.0007 3.42507e-08 0 3.44247e-08 0 3.44277e-08 0.0007 3.44307e-08 0 3.49647e-08 0 3.49677e-08 0.0007 3.49707e-08 0 3.51447e-08 0 3.51477e-08 0.0007 3.51507e-08 0 3.56847e-08 0 3.56877e-08 0.0007 3.56907e-08 0 3.58647e-08 0 3.58677e-08 0.0007 3.58707e-08 0 3.64047e-08 0 3.64077e-08 0.0007 3.64107e-08 0 3.65847e-08 0 3.65877e-08 0.0007 3.65907e-08 0 3.71247e-08 0 3.71277e-08 0.0007 3.71307e-08 0 3.73047e-08 0 3.73077e-08 0.0007 3.73107e-08 0 3.78447e-08 0 3.78477e-08 0.0007 3.78507e-08 0 3.80247e-08 0 3.80277e-08 0.0007 3.80307e-08 0 3.85647e-08 0 3.85677e-08 0.0007 3.85707e-08 0 3.87447e-08 0 3.87477e-08 0.0007 3.87507e-08 0 3.92847e-08 0 3.92877e-08 0.0007 3.92907e-08 0 3.94647e-08 0 3.94677e-08 0.0007 3.94707e-08 0 4.00047e-08 0 4.00077e-08 0.0007 4.00107e-08 0 4.01847e-08 0 4.01877e-08 0.0007 4.01907e-08 0 4.07247e-08 0 4.07277e-08 0.0007 4.07307e-08 0 4.09047e-08 0 4.09077e-08 0.0007 4.09107e-08 0 4.14447e-08 0 4.14477e-08 0.0007 4.14507e-08 0 4.16247e-08 0 4.16277e-08 0.0007 4.16307e-08 0 4.21647e-08 0 4.21677e-08 0.0007 4.21707e-08 0 4.23447e-08 0 4.23477e-08 0.0007 4.23507e-08 0 4.28847e-08 0 4.28877e-08 0.0007 4.28907e-08 0 4.30647e-08 0 4.30677e-08 0.0007 4.30707e-08 0 4.36047e-08 0 4.36077e-08 0.0007 4.36107e-08 0 4.37847e-08 0 4.37877e-08 0.0007 4.37907e-08 0 4.43247e-08 0 4.43277e-08 0.0007 4.43307e-08 0 4.45047e-08 0 4.45077e-08 0.0007 4.45107e-08 0 4.50447e-08 0 4.50477e-08 0.0007 4.50507e-08 0 4.52247e-08 0 4.52277e-08 0.0007 4.52307e-08 0 4.57647e-08 0 4.57677e-08 0.0007 4.57707e-08 0 4.59447e-08 0 4.59477e-08 0.0007 4.59507e-08 0)
IA1|C 0 A1  PWL(0 0 7.791e-10 0 7.821e-10 0.0007 7.851e-10 0 9.591e-10 0 9.621e-10 0.0007 9.651e-10 0 1.1391e-09 0 1.1421e-09 0.0007 1.1451e-09 0 1.3191e-09 0 1.3221e-09 0.0007 1.3251e-09 0 2.2191e-09 0 2.2221e-09 0.0007 2.2251e-09 0 2.3991e-09 0 2.4021e-09 0.0007 2.4051e-09 0 2.5791e-09 0 2.5821e-09 0.0007 2.5851e-09 0 2.7591e-09 0 2.7621e-09 0.0007 2.7651e-09 0 3.6591e-09 0 3.6621e-09 0.0007 3.6651e-09 0 3.8391e-09 0 3.8421e-09 0.0007 3.8451e-09 0 4.0191e-09 0 4.0221e-09 0.0007 4.0251e-09 0 4.1991e-09 0 4.2021e-09 0.0007 4.2051e-09 0 5.0991e-09 0 5.1021e-09 0.0007 5.1051e-09 0 5.2791e-09 0 5.2821e-09 0.0007 5.2851e-09 0 5.4591e-09 0 5.4621e-09 0.0007 5.4651e-09 0 5.6391e-09 0 5.6421e-09 0.0007 5.6451e-09 0 6.5391e-09 0 6.5421e-09 0.0007 6.5451e-09 0 6.7191e-09 0 6.7221e-09 0.0007 6.7251e-09 0 6.8991e-09 0 6.9021e-09 0.0007 6.9051e-09 0 7.0791e-09 0 7.0821e-09 0.0007 7.0851e-09 0 7.9791e-09 0 7.9821e-09 0.0007 7.9851e-09 0 8.1591e-09 0 8.1621e-09 0.0007 8.1651e-09 0 8.3391e-09 0 8.3421e-09 0.0007 8.3451e-09 0 8.5191e-09 0 8.5221e-09 0.0007 8.5251e-09 0 9.4191e-09 0 9.4221e-09 0.0007 9.4251e-09 0 9.5991e-09 0 9.6021e-09 0.0007 9.6051e-09 0 9.7791e-09 0 9.7821e-09 0.0007 9.7851e-09 0 9.9591e-09 0 9.9621e-09 0.0007 9.9651e-09 0 1.08591e-08 0 1.08621e-08 0.0007 1.08651e-08 0 1.10391e-08 0 1.10421e-08 0.0007 1.10451e-08 0 1.12191e-08 0 1.12221e-08 0.0007 1.12251e-08 0 1.13991e-08 0 1.14021e-08 0.0007 1.14051e-08 0 1.22991e-08 0 1.23021e-08 0.0007 1.23051e-08 0 1.24791e-08 0 1.24821e-08 0.0007 1.24851e-08 0 1.26591e-08 0 1.26621e-08 0.0007 1.26651e-08 0 1.28391e-08 0 1.28421e-08 0.0007 1.28451e-08 0 1.37391e-08 0 1.37421e-08 0.0007 1.37451e-08 0 1.39191e-08 0 1.39221e-08 0.0007 1.39251e-08 0 1.40991e-08 0 1.41021e-08 0.0007 1.41051e-08 0 1.42791e-08 0 1.42821e-08 0.0007 1.42851e-08 0 1.51791e-08 0 1.51821e-08 0.0007 1.51851e-08 0 1.53591e-08 0 1.53621e-08 0.0007 1.53651e-08 0 1.55391e-08 0 1.55421e-08 0.0007 1.55451e-08 0 1.57191e-08 0 1.57221e-08 0.0007 1.57251e-08 0 1.66191e-08 0 1.66221e-08 0.0007 1.66251e-08 0 1.67991e-08 0 1.68021e-08 0.0007 1.68051e-08 0 1.69791e-08 0 1.69821e-08 0.0007 1.69851e-08 0 1.71591e-08 0 1.71621e-08 0.0007 1.71651e-08 0 1.80591e-08 0 1.80621e-08 0.0007 1.80651e-08 0 1.82391e-08 0 1.82421e-08 0.0007 1.82451e-08 0 1.84191e-08 0 1.84221e-08 0.0007 1.84251e-08 0 1.85991e-08 0 1.86021e-08 0.0007 1.86051e-08 0 1.94991e-08 0 1.95021e-08 0.0007 1.95051e-08 0 1.96791e-08 0 1.96821e-08 0.0007 1.96851e-08 0 1.98591e-08 0 1.98621e-08 0.0007 1.98651e-08 0 2.00391e-08 0 2.00421e-08 0.0007 2.00451e-08 0 2.09391e-08 0 2.09421e-08 0.0007 2.09451e-08 0 2.11191e-08 0 2.11221e-08 0.0007 2.11251e-08 0 2.12991e-08 0 2.13021e-08 0.0007 2.13051e-08 0 2.14791e-08 0 2.14821e-08 0.0007 2.14851e-08 0 2.23791e-08 0 2.23821e-08 0.0007 2.23851e-08 0 2.25591e-08 0 2.25621e-08 0.0007 2.25651e-08 0 2.27391e-08 0 2.27421e-08 0.0007 2.27451e-08 0 2.29191e-08 0 2.29221e-08 0.0007 2.29251e-08 0 2.38191e-08 0 2.38221e-08 0.0007 2.38251e-08 0 2.39991e-08 0 2.40021e-08 0.0007 2.40051e-08 0 2.41791e-08 0 2.41821e-08 0.0007 2.41851e-08 0 2.43591e-08 0 2.43621e-08 0.0007 2.43651e-08 0 2.52591e-08 0 2.52621e-08 0.0007 2.52651e-08 0 2.54391e-08 0 2.54421e-08 0.0007 2.54451e-08 0 2.56191e-08 0 2.56221e-08 0.0007 2.56251e-08 0 2.57991e-08 0 2.58021e-08 0.0007 2.58051e-08 0 2.66991e-08 0 2.67021e-08 0.0007 2.67051e-08 0 2.68791e-08 0 2.68821e-08 0.0007 2.68851e-08 0 2.70591e-08 0 2.70621e-08 0.0007 2.70651e-08 0 2.72391e-08 0 2.72421e-08 0.0007 2.72451e-08 0 2.81391e-08 0 2.81421e-08 0.0007 2.81451e-08 0 2.83191e-08 0 2.83221e-08 0.0007 2.83251e-08 0 2.84991e-08 0 2.85021e-08 0.0007 2.85051e-08 0 2.86791e-08 0 2.86821e-08 0.0007 2.86851e-08 0 2.95791e-08 0 2.95821e-08 0.0007 2.95851e-08 0 2.97591e-08 0 2.97621e-08 0.0007 2.97651e-08 0 2.99391e-08 0 2.99421e-08 0.0007 2.99451e-08 0 3.01191e-08 0 3.01221e-08 0.0007 3.01251e-08 0 3.10191e-08 0 3.10221e-08 0.0007 3.10251e-08 0 3.11991e-08 0 3.12021e-08 0.0007 3.12051e-08 0 3.13791e-08 0 3.13821e-08 0.0007 3.13851e-08 0 3.15591e-08 0 3.15621e-08 0.0007 3.15651e-08 0 3.24591e-08 0 3.24621e-08 0.0007 3.24651e-08 0 3.26391e-08 0 3.26421e-08 0.0007 3.26451e-08 0 3.28191e-08 0 3.28221e-08 0.0007 3.28251e-08 0 3.29991e-08 0 3.30021e-08 0.0007 3.30051e-08 0 3.38991e-08 0 3.39021e-08 0.0007 3.39051e-08 0 3.40791e-08 0 3.40821e-08 0.0007 3.40851e-08 0 3.42591e-08 0 3.42621e-08 0.0007 3.42651e-08 0 3.44391e-08 0 3.44421e-08 0.0007 3.44451e-08 0 3.53391e-08 0 3.53421e-08 0.0007 3.53451e-08 0 3.55191e-08 0 3.55221e-08 0.0007 3.55251e-08 0 3.56991e-08 0 3.57021e-08 0.0007 3.57051e-08 0 3.58791e-08 0 3.58821e-08 0.0007 3.58851e-08 0 3.67791e-08 0 3.67821e-08 0.0007 3.67851e-08 0 3.69591e-08 0 3.69621e-08 0.0007 3.69651e-08 0 3.71391e-08 0 3.71421e-08 0.0007 3.71451e-08 0 3.73191e-08 0 3.73221e-08 0.0007 3.73251e-08 0 3.82191e-08 0 3.82221e-08 0.0007 3.82251e-08 0 3.83991e-08 0 3.84021e-08 0.0007 3.84051e-08 0 3.85791e-08 0 3.85821e-08 0.0007 3.85851e-08 0 3.87591e-08 0 3.87621e-08 0.0007 3.87651e-08 0 3.96591e-08 0 3.96621e-08 0.0007 3.96651e-08 0 3.98391e-08 0 3.98421e-08 0.0007 3.98451e-08 0 4.00191e-08 0 4.00221e-08 0.0007 4.00251e-08 0 4.01991e-08 0 4.02021e-08 0.0007 4.02051e-08 0 4.10991e-08 0 4.11021e-08 0.0007 4.11051e-08 0 4.12791e-08 0 4.12821e-08 0.0007 4.12851e-08 0 4.14591e-08 0 4.14621e-08 0.0007 4.14651e-08 0 4.16391e-08 0 4.16421e-08 0.0007 4.16451e-08 0 4.25391e-08 0 4.25421e-08 0.0007 4.25451e-08 0 4.27191e-08 0 4.27221e-08 0.0007 4.27251e-08 0 4.28991e-08 0 4.29021e-08 0.0007 4.29051e-08 0 4.30791e-08 0 4.30821e-08 0.0007 4.30851e-08 0 4.39791e-08 0 4.39821e-08 0.0007 4.39851e-08 0 4.41591e-08 0 4.41621e-08 0.0007 4.41651e-08 0 4.43391e-08 0 4.43421e-08 0.0007 4.43451e-08 0 4.45191e-08 0 4.45221e-08 0.0007 4.45251e-08 0 4.54191e-08 0 4.54221e-08 0.0007 4.54251e-08 0 4.55991e-08 0 4.56021e-08 0.0007 4.56051e-08 0 4.57791e-08 0 4.57821e-08 0.0007 4.57851e-08 0 4.59591e-08 0 4.59621e-08 0.0007 4.59651e-08 0)
IB1|D 0 B1  PWL(0 0 1.5135e-09 0 1.5165e-09 0.0007 1.5195e-09 0 1.6935e-09 0 1.6965e-09 0.0007 1.6995e-09 0 1.8735e-09 0 1.8765e-09 0.0007 1.8795e-09 0 2.0535e-09 0 2.0565e-09 0.0007 2.0595e-09 0 2.2335e-09 0 2.2365e-09 0.0007 2.2395e-09 0 2.4135e-09 0 2.4165e-09 0.0007 2.4195e-09 0 2.5935e-09 0 2.5965e-09 0.0007 2.5995e-09 0 2.7735e-09 0 2.7765e-09 0.0007 2.7795e-09 0 4.3935e-09 0 4.3965e-09 0.0007 4.3995e-09 0 4.5735e-09 0 4.5765e-09 0.0007 4.5795e-09 0 4.7535e-09 0 4.7565e-09 0.0007 4.7595e-09 0 4.9335e-09 0 4.9365e-09 0.0007 4.9395e-09 0 5.1135e-09 0 5.1165e-09 0.0007 5.1195e-09 0 5.2935e-09 0 5.2965e-09 0.0007 5.2995e-09 0 5.4735e-09 0 5.4765e-09 0.0007 5.4795e-09 0 5.6535e-09 0 5.6565e-09 0.0007 5.6595e-09 0 7.2735e-09 0 7.2765e-09 0.0007 7.2795e-09 0 7.4535e-09 0 7.4565e-09 0.0007 7.4595e-09 0 7.6335e-09 0 7.6365e-09 0.0007 7.6395e-09 0 7.8135e-09 0 7.8165e-09 0.0007 7.8195e-09 0 7.9935e-09 0 7.9965e-09 0.0007 7.9995e-09 0 8.1735e-09 0 8.1765e-09 0.0007 8.1795e-09 0 8.3535e-09 0 8.3565e-09 0.0007 8.3595e-09 0 8.5335e-09 0 8.5365e-09 0.0007 8.5395e-09 0 1.01535e-08 0 1.01565e-08 0.0007 1.01595e-08 0 1.03335e-08 0 1.03365e-08 0.0007 1.03395e-08 0 1.05135e-08 0 1.05165e-08 0.0007 1.05195e-08 0 1.06935e-08 0 1.06965e-08 0.0007 1.06995e-08 0 1.08735e-08 0 1.08765e-08 0.0007 1.08795e-08 0 1.10535e-08 0 1.10565e-08 0.0007 1.10595e-08 0 1.12335e-08 0 1.12365e-08 0.0007 1.12395e-08 0 1.14135e-08 0 1.14165e-08 0.0007 1.14195e-08 0 1.30335e-08 0 1.30365e-08 0.0007 1.30395e-08 0 1.32135e-08 0 1.32165e-08 0.0007 1.32195e-08 0 1.33935e-08 0 1.33965e-08 0.0007 1.33995e-08 0 1.35735e-08 0 1.35765e-08 0.0007 1.35795e-08 0 1.37535e-08 0 1.37565e-08 0.0007 1.37595e-08 0 1.39335e-08 0 1.39365e-08 0.0007 1.39395e-08 0 1.41135e-08 0 1.41165e-08 0.0007 1.41195e-08 0 1.42935e-08 0 1.42965e-08 0.0007 1.42995e-08 0 1.59135e-08 0 1.59165e-08 0.0007 1.59195e-08 0 1.60935e-08 0 1.60965e-08 0.0007 1.60995e-08 0 1.62735e-08 0 1.62765e-08 0.0007 1.62795e-08 0 1.64535e-08 0 1.64565e-08 0.0007 1.64595e-08 0 1.66335e-08 0 1.66365e-08 0.0007 1.66395e-08 0 1.68135e-08 0 1.68165e-08 0.0007 1.68195e-08 0 1.69935e-08 0 1.69965e-08 0.0007 1.69995e-08 0 1.71735e-08 0 1.71765e-08 0.0007 1.71795e-08 0 1.87935e-08 0 1.87965e-08 0.0007 1.87995e-08 0 1.89735e-08 0 1.89765e-08 0.0007 1.89795e-08 0 1.91535e-08 0 1.91565e-08 0.0007 1.91595e-08 0 1.93335e-08 0 1.93365e-08 0.0007 1.93395e-08 0 1.95135e-08 0 1.95165e-08 0.0007 1.95195e-08 0 1.96935e-08 0 1.96965e-08 0.0007 1.96995e-08 0 1.98735e-08 0 1.98765e-08 0.0007 1.98795e-08 0 2.00535e-08 0 2.00565e-08 0.0007 2.00595e-08 0 2.16735e-08 0 2.16765e-08 0.0007 2.16795e-08 0 2.18535e-08 0 2.18565e-08 0.0007 2.18595e-08 0 2.20335e-08 0 2.20365e-08 0.0007 2.20395e-08 0 2.22135e-08 0 2.22165e-08 0.0007 2.22195e-08 0 2.23935e-08 0 2.23965e-08 0.0007 2.23995e-08 0 2.25735e-08 0 2.25765e-08 0.0007 2.25795e-08 0 2.27535e-08 0 2.27565e-08 0.0007 2.27595e-08 0 2.29335e-08 0 2.29365e-08 0.0007 2.29395e-08 0 2.45535e-08 0 2.45565e-08 0.0007 2.45595e-08 0 2.47335e-08 0 2.47365e-08 0.0007 2.47395e-08 0 2.49135e-08 0 2.49165e-08 0.0007 2.49195e-08 0 2.50935e-08 0 2.50965e-08 0.0007 2.50995e-08 0 2.52735e-08 0 2.52765e-08 0.0007 2.52795e-08 0 2.54535e-08 0 2.54565e-08 0.0007 2.54595e-08 0 2.56335e-08 0 2.56365e-08 0.0007 2.56395e-08 0 2.58135e-08 0 2.58165e-08 0.0007 2.58195e-08 0 2.74335e-08 0 2.74365e-08 0.0007 2.74395e-08 0 2.76135e-08 0 2.76165e-08 0.0007 2.76195e-08 0 2.77935e-08 0 2.77965e-08 0.0007 2.77995e-08 0 2.79735e-08 0 2.79765e-08 0.0007 2.79795e-08 0 2.81535e-08 0 2.81565e-08 0.0007 2.81595e-08 0 2.83335e-08 0 2.83365e-08 0.0007 2.83395e-08 0 2.85135e-08 0 2.85165e-08 0.0007 2.85195e-08 0 2.86935e-08 0 2.86965e-08 0.0007 2.86995e-08 0 3.03135e-08 0 3.03165e-08 0.0007 3.03195e-08 0 3.04935e-08 0 3.04965e-08 0.0007 3.04995e-08 0 3.06735e-08 0 3.06765e-08 0.0007 3.06795e-08 0 3.08535e-08 0 3.08565e-08 0.0007 3.08595e-08 0 3.10335e-08 0 3.10365e-08 0.0007 3.10395e-08 0 3.12135e-08 0 3.12165e-08 0.0007 3.12195e-08 0 3.13935e-08 0 3.13965e-08 0.0007 3.13995e-08 0 3.15735e-08 0 3.15765e-08 0.0007 3.15795e-08 0 3.31935e-08 0 3.31965e-08 0.0007 3.31995e-08 0 3.33735e-08 0 3.33765e-08 0.0007 3.33795e-08 0 3.35535e-08 0 3.35565e-08 0.0007 3.35595e-08 0 3.37335e-08 0 3.37365e-08 0.0007 3.37395e-08 0 3.39135e-08 0 3.39165e-08 0.0007 3.39195e-08 0 3.40935e-08 0 3.40965e-08 0.0007 3.40995e-08 0 3.42735e-08 0 3.42765e-08 0.0007 3.42795e-08 0 3.44535e-08 0 3.44565e-08 0.0007 3.44595e-08 0 3.60735e-08 0 3.60765e-08 0.0007 3.60795e-08 0 3.62535e-08 0 3.62565e-08 0.0007 3.62595e-08 0 3.64335e-08 0 3.64365e-08 0.0007 3.64395e-08 0 3.66135e-08 0 3.66165e-08 0.0007 3.66195e-08 0 3.67935e-08 0 3.67965e-08 0.0007 3.67995e-08 0 3.69735e-08 0 3.69765e-08 0.0007 3.69795e-08 0 3.71535e-08 0 3.71565e-08 0.0007 3.71595e-08 0 3.73335e-08 0 3.73365e-08 0.0007 3.73395e-08 0 3.89535e-08 0 3.89565e-08 0.0007 3.89595e-08 0 3.91335e-08 0 3.91365e-08 0.0007 3.91395e-08 0 3.93135e-08 0 3.93165e-08 0.0007 3.93195e-08 0 3.94935e-08 0 3.94965e-08 0.0007 3.94995e-08 0 3.96735e-08 0 3.96765e-08 0.0007 3.96795e-08 0 3.98535e-08 0 3.98565e-08 0.0007 3.98595e-08 0 4.00335e-08 0 4.00365e-08 0.0007 4.00395e-08 0 4.02135e-08 0 4.02165e-08 0.0007 4.02195e-08 0 4.18335e-08 0 4.18365e-08 0.0007 4.18395e-08 0 4.20135e-08 0 4.20165e-08 0.0007 4.20195e-08 0 4.21935e-08 0 4.21965e-08 0.0007 4.21995e-08 0 4.23735e-08 0 4.23765e-08 0.0007 4.23795e-08 0 4.25535e-08 0 4.25565e-08 0.0007 4.25595e-08 0 4.27335e-08 0 4.27365e-08 0.0007 4.27395e-08 0 4.29135e-08 0 4.29165e-08 0.0007 4.29195e-08 0 4.30935e-08 0 4.30965e-08 0.0007 4.30995e-08 0 4.47135e-08 0 4.47165e-08 0.0007 4.47195e-08 0 4.48935e-08 0 4.48965e-08 0.0007 4.48995e-08 0 4.50735e-08 0 4.50765e-08 0.0007 4.50795e-08 0 4.52535e-08 0 4.52565e-08 0.0007 4.52595e-08 0 4.54335e-08 0 4.54365e-08 0.0007 4.54395e-08 0 4.56135e-08 0 4.56165e-08 0.0007 4.56195e-08 0 4.57935e-08 0 4.57965e-08 0.0007 4.57995e-08 0 4.59735e-08 0 4.59765e-08 0.0007 4.59795e-08 0)
IA2|E 0 A2  PWL(0 0 2.9679e-09 0 2.9709e-09 0.0007 2.9739e-09 0 3.1479e-09 0 3.1509e-09 0.0007 3.1539e-09 0 3.3279e-09 0 3.3309e-09 0.0007 3.3339e-09 0 3.5079e-09 0 3.5109e-09 0.0007 3.5139e-09 0 3.6879e-09 0 3.6909e-09 0.0007 3.6939e-09 0 3.8679e-09 0 3.8709e-09 0.0007 3.8739e-09 0 4.0479e-09 0 4.0509e-09 0.0007 4.0539e-09 0 4.2279e-09 0 4.2309e-09 0.0007 4.2339e-09 0 4.4079e-09 0 4.4109e-09 0.0007 4.4139e-09 0 4.5879e-09 0 4.5909e-09 0.0007 4.5939e-09 0 4.7679e-09 0 4.7709e-09 0.0007 4.7739e-09 0 4.9479e-09 0 4.9509e-09 0.0007 4.9539e-09 0 5.1279e-09 0 5.1309e-09 0.0007 5.1339e-09 0 5.3079e-09 0 5.3109e-09 0.0007 5.3139e-09 0 5.4879e-09 0 5.4909e-09 0.0007 5.4939e-09 0 5.6679e-09 0 5.6709e-09 0.0007 5.6739e-09 0 8.7279e-09 0 8.7309e-09 0.0007 8.7339e-09 0 8.9079e-09 0 8.9109e-09 0.0007 8.9139e-09 0 9.0879e-09 0 9.0909e-09 0.0007 9.0939e-09 0 9.2679e-09 0 9.2709e-09 0.0007 9.2739e-09 0 9.4479e-09 0 9.4509e-09 0.0007 9.4539e-09 0 9.6279e-09 0 9.6309e-09 0.0007 9.6339e-09 0 9.8079e-09 0 9.8109e-09 0.0007 9.8139e-09 0 9.9879e-09 0 9.9909e-09 0.0007 9.9939e-09 0 1.01679e-08 0 1.01709e-08 0.0007 1.01739e-08 0 1.03479e-08 0 1.03509e-08 0.0007 1.03539e-08 0 1.05279e-08 0 1.05309e-08 0.0007 1.05339e-08 0 1.07079e-08 0 1.07109e-08 0.0007 1.07139e-08 0 1.08879e-08 0 1.08909e-08 0.0007 1.08939e-08 0 1.10679e-08 0 1.10709e-08 0.0007 1.10739e-08 0 1.12479e-08 0 1.12509e-08 0.0007 1.12539e-08 0 1.14279e-08 0 1.14309e-08 0.0007 1.14339e-08 0 1.44879e-08 0 1.44909e-08 0.0007 1.44939e-08 0 1.46679e-08 0 1.46709e-08 0.0007 1.46739e-08 0 1.48479e-08 0 1.48509e-08 0.0007 1.48539e-08 0 1.50279e-08 0 1.50309e-08 0.0007 1.50339e-08 0 1.52079e-08 0 1.52109e-08 0.0007 1.52139e-08 0 1.53879e-08 0 1.53909e-08 0.0007 1.53939e-08 0 1.55679e-08 0 1.55709e-08 0.0007 1.55739e-08 0 1.57479e-08 0 1.57509e-08 0.0007 1.57539e-08 0 1.59279e-08 0 1.59309e-08 0.0007 1.59339e-08 0 1.61079e-08 0 1.61109e-08 0.0007 1.61139e-08 0 1.62879e-08 0 1.62909e-08 0.0007 1.62939e-08 0 1.64679e-08 0 1.64709e-08 0.0007 1.64739e-08 0 1.66479e-08 0 1.66509e-08 0.0007 1.66539e-08 0 1.68279e-08 0 1.68309e-08 0.0007 1.68339e-08 0 1.70079e-08 0 1.70109e-08 0.0007 1.70139e-08 0 1.71879e-08 0 1.71909e-08 0.0007 1.71939e-08 0 2.02479e-08 0 2.02509e-08 0.0007 2.02539e-08 0 2.04279e-08 0 2.04309e-08 0.0007 2.04339e-08 0 2.06079e-08 0 2.06109e-08 0.0007 2.06139e-08 0 2.07879e-08 0 2.07909e-08 0.0007 2.07939e-08 0 2.09679e-08 0 2.09709e-08 0.0007 2.09739e-08 0 2.11479e-08 0 2.11509e-08 0.0007 2.11539e-08 0 2.13279e-08 0 2.13309e-08 0.0007 2.13339e-08 0 2.15079e-08 0 2.15109e-08 0.0007 2.15139e-08 0 2.16879e-08 0 2.16909e-08 0.0007 2.16939e-08 0 2.18679e-08 0 2.18709e-08 0.0007 2.18739e-08 0 2.20479e-08 0 2.20509e-08 0.0007 2.20539e-08 0 2.22279e-08 0 2.22309e-08 0.0007 2.22339e-08 0 2.24079e-08 0 2.24109e-08 0.0007 2.24139e-08 0 2.25879e-08 0 2.25909e-08 0.0007 2.25939e-08 0 2.27679e-08 0 2.27709e-08 0.0007 2.27739e-08 0 2.29479e-08 0 2.29509e-08 0.0007 2.29539e-08 0 2.60079e-08 0 2.60109e-08 0.0007 2.60139e-08 0 2.61879e-08 0 2.61909e-08 0.0007 2.61939e-08 0 2.63679e-08 0 2.63709e-08 0.0007 2.63739e-08 0 2.65479e-08 0 2.65509e-08 0.0007 2.65539e-08 0 2.67279e-08 0 2.67309e-08 0.0007 2.67339e-08 0 2.69079e-08 0 2.69109e-08 0.0007 2.69139e-08 0 2.70879e-08 0 2.70909e-08 0.0007 2.70939e-08 0 2.72679e-08 0 2.72709e-08 0.0007 2.72739e-08 0 2.74479e-08 0 2.74509e-08 0.0007 2.74539e-08 0 2.76279e-08 0 2.76309e-08 0.0007 2.76339e-08 0 2.78079e-08 0 2.78109e-08 0.0007 2.78139e-08 0 2.79879e-08 0 2.79909e-08 0.0007 2.79939e-08 0 2.81679e-08 0 2.81709e-08 0.0007 2.81739e-08 0 2.83479e-08 0 2.83509e-08 0.0007 2.83539e-08 0 2.85279e-08 0 2.85309e-08 0.0007 2.85339e-08 0 2.87079e-08 0 2.87109e-08 0.0007 2.87139e-08 0 3.17679e-08 0 3.17709e-08 0.0007 3.17739e-08 0 3.19479e-08 0 3.19509e-08 0.0007 3.19539e-08 0 3.21279e-08 0 3.21309e-08 0.0007 3.21339e-08 0 3.23079e-08 0 3.23109e-08 0.0007 3.23139e-08 0 3.24879e-08 0 3.24909e-08 0.0007 3.24939e-08 0 3.26679e-08 0 3.26709e-08 0.0007 3.26739e-08 0 3.28479e-08 0 3.28509e-08 0.0007 3.28539e-08 0 3.30279e-08 0 3.30309e-08 0.0007 3.30339e-08 0 3.32079e-08 0 3.32109e-08 0.0007 3.32139e-08 0 3.33879e-08 0 3.33909e-08 0.0007 3.33939e-08 0 3.35679e-08 0 3.35709e-08 0.0007 3.35739e-08 0 3.37479e-08 0 3.37509e-08 0.0007 3.37539e-08 0 3.39279e-08 0 3.39309e-08 0.0007 3.39339e-08 0 3.41079e-08 0 3.41109e-08 0.0007 3.41139e-08 0 3.42879e-08 0 3.42909e-08 0.0007 3.42939e-08 0 3.44679e-08 0 3.44709e-08 0.0007 3.44739e-08 0 3.75279e-08 0 3.75309e-08 0.0007 3.75339e-08 0 3.77079e-08 0 3.77109e-08 0.0007 3.77139e-08 0 3.78879e-08 0 3.78909e-08 0.0007 3.78939e-08 0 3.80679e-08 0 3.80709e-08 0.0007 3.80739e-08 0 3.82479e-08 0 3.82509e-08 0.0007 3.82539e-08 0 3.84279e-08 0 3.84309e-08 0.0007 3.84339e-08 0 3.86079e-08 0 3.86109e-08 0.0007 3.86139e-08 0 3.87879e-08 0 3.87909e-08 0.0007 3.87939e-08 0 3.89679e-08 0 3.89709e-08 0.0007 3.89739e-08 0 3.91479e-08 0 3.91509e-08 0.0007 3.91539e-08 0 3.93279e-08 0 3.93309e-08 0.0007 3.93339e-08 0 3.95079e-08 0 3.95109e-08 0.0007 3.95139e-08 0 3.96879e-08 0 3.96909e-08 0.0007 3.96939e-08 0 3.98679e-08 0 3.98709e-08 0.0007 3.98739e-08 0 4.00479e-08 0 4.00509e-08 0.0007 4.00539e-08 0 4.02279e-08 0 4.02309e-08 0.0007 4.02339e-08 0 4.32879e-08 0 4.32909e-08 0.0007 4.32939e-08 0 4.34679e-08 0 4.34709e-08 0.0007 4.34739e-08 0 4.36479e-08 0 4.36509e-08 0.0007 4.36539e-08 0 4.38279e-08 0 4.38309e-08 0.0007 4.38339e-08 0 4.40079e-08 0 4.40109e-08 0.0007 4.40139e-08 0 4.41879e-08 0 4.41909e-08 0.0007 4.41939e-08 0 4.43679e-08 0 4.43709e-08 0.0007 4.43739e-08 0 4.45479e-08 0 4.45509e-08 0.0007 4.45539e-08 0 4.47279e-08 0 4.47309e-08 0.0007 4.47339e-08 0 4.49079e-08 0 4.49109e-08 0.0007 4.49139e-08 0 4.50879e-08 0 4.50909e-08 0.0007 4.50939e-08 0 4.52679e-08 0 4.52709e-08 0.0007 4.52739e-08 0 4.54479e-08 0 4.54509e-08 0.0007 4.54539e-08 0 4.56279e-08 0 4.56309e-08 0.0007 4.56339e-08 0 4.58079e-08 0 4.58109e-08 0.0007 4.58139e-08 0 4.59879e-08 0 4.59909e-08 0.0007 4.59939e-08 0)
IB2|F 0 B2  PWL(0 0 5.8623e-09 0 5.8653e-09 0.0007 5.8683e-09 0 6.0423e-09 0 6.0453e-09 0.0007 6.0483e-09 0 6.2223e-09 0 6.2253e-09 0.0007 6.2283e-09 0 6.4023e-09 0 6.4053e-09 0.0007 6.4083e-09 0 6.5823e-09 0 6.5853e-09 0.0007 6.5883e-09 0 6.7623e-09 0 6.7653e-09 0.0007 6.7683e-09 0 6.9423e-09 0 6.9453e-09 0.0007 6.9483e-09 0 7.1223e-09 0 7.1253e-09 0.0007 7.1283e-09 0 7.3023e-09 0 7.3053e-09 0.0007 7.3083e-09 0 7.4823e-09 0 7.4853e-09 0.0007 7.4883e-09 0 7.6623e-09 0 7.6653e-09 0.0007 7.6683e-09 0 7.8423e-09 0 7.8453e-09 0.0007 7.8483e-09 0 8.0223e-09 0 8.0253e-09 0.0007 8.0283e-09 0 8.2023e-09 0 8.2053e-09 0.0007 8.2083e-09 0 8.3823e-09 0 8.3853e-09 0.0007 8.3883e-09 0 8.5623e-09 0 8.5653e-09 0.0007 8.5683e-09 0 8.7423e-09 0 8.7453e-09 0.0007 8.7483e-09 0 8.9223e-09 0 8.9253e-09 0.0007 8.9283e-09 0 9.1023e-09 0 9.1053e-09 0.0007 9.1083e-09 0 9.2823e-09 0 9.2853e-09 0.0007 9.2883e-09 0 9.4623e-09 0 9.4653e-09 0.0007 9.4683e-09 0 9.6423e-09 0 9.6453e-09 0.0007 9.6483e-09 0 9.8223e-09 0 9.8253e-09 0.0007 9.8283e-09 0 1.00023e-08 0 1.00053e-08 0.0007 1.00083e-08 0 1.01823e-08 0 1.01853e-08 0.0007 1.01883e-08 0 1.03623e-08 0 1.03653e-08 0.0007 1.03683e-08 0 1.05423e-08 0 1.05453e-08 0.0007 1.05483e-08 0 1.07223e-08 0 1.07253e-08 0.0007 1.07283e-08 0 1.09023e-08 0 1.09053e-08 0.0007 1.09083e-08 0 1.10823e-08 0 1.10853e-08 0.0007 1.10883e-08 0 1.12623e-08 0 1.12653e-08 0.0007 1.12683e-08 0 1.14423e-08 0 1.14453e-08 0.0007 1.14483e-08 0 1.73823e-08 0 1.73853e-08 0.0007 1.73883e-08 0 1.75623e-08 0 1.75653e-08 0.0007 1.75683e-08 0 1.77423e-08 0 1.77453e-08 0.0007 1.77483e-08 0 1.79223e-08 0 1.79253e-08 0.0007 1.79283e-08 0 1.81023e-08 0 1.81053e-08 0.0007 1.81083e-08 0 1.82823e-08 0 1.82853e-08 0.0007 1.82883e-08 0 1.84623e-08 0 1.84653e-08 0.0007 1.84683e-08 0 1.86423e-08 0 1.86453e-08 0.0007 1.86483e-08 0 1.88223e-08 0 1.88253e-08 0.0007 1.88283e-08 0 1.90023e-08 0 1.90053e-08 0.0007 1.90083e-08 0 1.91823e-08 0 1.91853e-08 0.0007 1.91883e-08 0 1.93623e-08 0 1.93653e-08 0.0007 1.93683e-08 0 1.95423e-08 0 1.95453e-08 0.0007 1.95483e-08 0 1.97223e-08 0 1.97253e-08 0.0007 1.97283e-08 0 1.99023e-08 0 1.99053e-08 0.0007 1.99083e-08 0 2.00823e-08 0 2.00853e-08 0.0007 2.00883e-08 0 2.02623e-08 0 2.02653e-08 0.0007 2.02683e-08 0 2.04423e-08 0 2.04453e-08 0.0007 2.04483e-08 0 2.06223e-08 0 2.06253e-08 0.0007 2.06283e-08 0 2.08023e-08 0 2.08053e-08 0.0007 2.08083e-08 0 2.09823e-08 0 2.09853e-08 0.0007 2.09883e-08 0 2.11623e-08 0 2.11653e-08 0.0007 2.11683e-08 0 2.13423e-08 0 2.13453e-08 0.0007 2.13483e-08 0 2.15223e-08 0 2.15253e-08 0.0007 2.15283e-08 0 2.17023e-08 0 2.17053e-08 0.0007 2.17083e-08 0 2.18823e-08 0 2.18853e-08 0.0007 2.18883e-08 0 2.20623e-08 0 2.20653e-08 0.0007 2.20683e-08 0 2.22423e-08 0 2.22453e-08 0.0007 2.22483e-08 0 2.24223e-08 0 2.24253e-08 0.0007 2.24283e-08 0 2.26023e-08 0 2.26053e-08 0.0007 2.26083e-08 0 2.27823e-08 0 2.27853e-08 0.0007 2.27883e-08 0 2.29623e-08 0 2.29653e-08 0.0007 2.29683e-08 0 2.89023e-08 0 2.89053e-08 0.0007 2.89083e-08 0 2.90823e-08 0 2.90853e-08 0.0007 2.90883e-08 0 2.92623e-08 0 2.92653e-08 0.0007 2.92683e-08 0 2.94423e-08 0 2.94453e-08 0.0007 2.94483e-08 0 2.96223e-08 0 2.96253e-08 0.0007 2.96283e-08 0 2.98023e-08 0 2.98053e-08 0.0007 2.98083e-08 0 2.99823e-08 0 2.99853e-08 0.0007 2.99883e-08 0 3.01623e-08 0 3.01653e-08 0.0007 3.01683e-08 0 3.03423e-08 0 3.03453e-08 0.0007 3.03483e-08 0 3.05223e-08 0 3.05253e-08 0.0007 3.05283e-08 0 3.07023e-08 0 3.07053e-08 0.0007 3.07083e-08 0 3.08823e-08 0 3.08853e-08 0.0007 3.08883e-08 0 3.10623e-08 0 3.10653e-08 0.0007 3.10683e-08 0 3.12423e-08 0 3.12453e-08 0.0007 3.12483e-08 0 3.14223e-08 0 3.14253e-08 0.0007 3.14283e-08 0 3.16023e-08 0 3.16053e-08 0.0007 3.16083e-08 0 3.17823e-08 0 3.17853e-08 0.0007 3.17883e-08 0 3.19623e-08 0 3.19653e-08 0.0007 3.19683e-08 0 3.21423e-08 0 3.21453e-08 0.0007 3.21483e-08 0 3.23223e-08 0 3.23253e-08 0.0007 3.23283e-08 0 3.25023e-08 0 3.25053e-08 0.0007 3.25083e-08 0 3.26823e-08 0 3.26853e-08 0.0007 3.26883e-08 0 3.28623e-08 0 3.28653e-08 0.0007 3.28683e-08 0 3.30423e-08 0 3.30453e-08 0.0007 3.30483e-08 0 3.32223e-08 0 3.32253e-08 0.0007 3.32283e-08 0 3.34023e-08 0 3.34053e-08 0.0007 3.34083e-08 0 3.35823e-08 0 3.35853e-08 0.0007 3.35883e-08 0 3.37623e-08 0 3.37653e-08 0.0007 3.37683e-08 0 3.39423e-08 0 3.39453e-08 0.0007 3.39483e-08 0 3.41223e-08 0 3.41253e-08 0.0007 3.41283e-08 0 3.43023e-08 0 3.43053e-08 0.0007 3.43083e-08 0 3.44823e-08 0 3.44853e-08 0.0007 3.44883e-08 0 4.04223e-08 0 4.04253e-08 0.0007 4.04283e-08 0 4.06023e-08 0 4.06053e-08 0.0007 4.06083e-08 0 4.07823e-08 0 4.07853e-08 0.0007 4.07883e-08 0 4.09623e-08 0 4.09653e-08 0.0007 4.09683e-08 0 4.11423e-08 0 4.11453e-08 0.0007 4.11483e-08 0 4.13223e-08 0 4.13253e-08 0.0007 4.13283e-08 0 4.15023e-08 0 4.15053e-08 0.0007 4.15083e-08 0 4.16823e-08 0 4.16853e-08 0.0007 4.16883e-08 0 4.18623e-08 0 4.18653e-08 0.0007 4.18683e-08 0 4.20423e-08 0 4.20453e-08 0.0007 4.20483e-08 0 4.22223e-08 0 4.22253e-08 0.0007 4.22283e-08 0 4.24023e-08 0 4.24053e-08 0.0007 4.24083e-08 0 4.25823e-08 0 4.25853e-08 0.0007 4.25883e-08 0 4.27623e-08 0 4.27653e-08 0.0007 4.27683e-08 0 4.29423e-08 0 4.29453e-08 0.0007 4.29483e-08 0 4.31223e-08 0 4.31253e-08 0.0007 4.31283e-08 0 4.33023e-08 0 4.33053e-08 0.0007 4.33083e-08 0 4.34823e-08 0 4.34853e-08 0.0007 4.34883e-08 0 4.36623e-08 0 4.36653e-08 0.0007 4.36683e-08 0 4.38423e-08 0 4.38453e-08 0.0007 4.38483e-08 0 4.40223e-08 0 4.40253e-08 0.0007 4.40283e-08 0 4.42023e-08 0 4.42053e-08 0.0007 4.42083e-08 0 4.43823e-08 0 4.43853e-08 0.0007 4.43883e-08 0 4.45623e-08 0 4.45653e-08 0.0007 4.45683e-08 0 4.47423e-08 0 4.47453e-08 0.0007 4.47483e-08 0 4.49223e-08 0 4.49253e-08 0.0007 4.49283e-08 0 4.51023e-08 0 4.51053e-08 0.0007 4.51083e-08 0 4.52823e-08 0 4.52853e-08 0.0007 4.52883e-08 0 4.54623e-08 0 4.54653e-08 0.0007 4.54683e-08 0 4.56423e-08 0 4.56453e-08 0.0007 4.56483e-08 0 4.58223e-08 0 4.58253e-08 0.0007 4.58283e-08 0 4.60023e-08 0 4.60053e-08 0.0007 4.60083e-08 0)
IA3|G 0 A3  PWL(0 0 1.16367e-08 0 1.16397e-08 0.0007 1.16427e-08 0 1.18167e-08 0 1.18197e-08 0.0007 1.18227e-08 0 1.19967e-08 0 1.19997e-08 0.0007 1.20027e-08 0 1.21767e-08 0 1.21797e-08 0.0007 1.21827e-08 0 1.23567e-08 0 1.23597e-08 0.0007 1.23627e-08 0 1.25367e-08 0 1.25397e-08 0.0007 1.25427e-08 0 1.27167e-08 0 1.27197e-08 0.0007 1.27227e-08 0 1.28967e-08 0 1.28997e-08 0.0007 1.29027e-08 0 1.30767e-08 0 1.30797e-08 0.0007 1.30827e-08 0 1.32567e-08 0 1.32597e-08 0.0007 1.32627e-08 0 1.34367e-08 0 1.34397e-08 0.0007 1.34427e-08 0 1.36167e-08 0 1.36197e-08 0.0007 1.36227e-08 0 1.37967e-08 0 1.37997e-08 0.0007 1.38027e-08 0 1.39767e-08 0 1.39797e-08 0.0007 1.39827e-08 0 1.41567e-08 0 1.41597e-08 0.0007 1.41627e-08 0 1.43367e-08 0 1.43397e-08 0.0007 1.43427e-08 0 1.45167e-08 0 1.45197e-08 0.0007 1.45227e-08 0 1.46967e-08 0 1.46997e-08 0.0007 1.47027e-08 0 1.48767e-08 0 1.48797e-08 0.0007 1.48827e-08 0 1.50567e-08 0 1.50597e-08 0.0007 1.50627e-08 0 1.52367e-08 0 1.52397e-08 0.0007 1.52427e-08 0 1.54167e-08 0 1.54197e-08 0.0007 1.54227e-08 0 1.55967e-08 0 1.55997e-08 0.0007 1.56027e-08 0 1.57767e-08 0 1.57797e-08 0.0007 1.57827e-08 0 1.59567e-08 0 1.59597e-08 0.0007 1.59627e-08 0 1.61367e-08 0 1.61397e-08 0.0007 1.61427e-08 0 1.63167e-08 0 1.63197e-08 0.0007 1.63227e-08 0 1.64967e-08 0 1.64997e-08 0.0007 1.65027e-08 0 1.66767e-08 0 1.66797e-08 0.0007 1.66827e-08 0 1.68567e-08 0 1.68597e-08 0.0007 1.68627e-08 0 1.70367e-08 0 1.70397e-08 0.0007 1.70427e-08 0 1.72167e-08 0 1.72197e-08 0.0007 1.72227e-08 0 1.73967e-08 0 1.73997e-08 0.0007 1.74027e-08 0 1.75767e-08 0 1.75797e-08 0.0007 1.75827e-08 0 1.77567e-08 0 1.77597e-08 0.0007 1.77627e-08 0 1.79367e-08 0 1.79397e-08 0.0007 1.79427e-08 0 1.81167e-08 0 1.81197e-08 0.0007 1.81227e-08 0 1.82967e-08 0 1.82997e-08 0.0007 1.83027e-08 0 1.84767e-08 0 1.84797e-08 0.0007 1.84827e-08 0 1.86567e-08 0 1.86597e-08 0.0007 1.86627e-08 0 1.88367e-08 0 1.88397e-08 0.0007 1.88427e-08 0 1.90167e-08 0 1.90197e-08 0.0007 1.90227e-08 0 1.91967e-08 0 1.91997e-08 0.0007 1.92027e-08 0 1.93767e-08 0 1.93797e-08 0.0007 1.93827e-08 0 1.95567e-08 0 1.95597e-08 0.0007 1.95627e-08 0 1.97367e-08 0 1.97397e-08 0.0007 1.97427e-08 0 1.99167e-08 0 1.99197e-08 0.0007 1.99227e-08 0 2.00967e-08 0 2.00997e-08 0.0007 2.01027e-08 0 2.02767e-08 0 2.02797e-08 0.0007 2.02827e-08 0 2.04567e-08 0 2.04597e-08 0.0007 2.04627e-08 0 2.06367e-08 0 2.06397e-08 0.0007 2.06427e-08 0 2.08167e-08 0 2.08197e-08 0.0007 2.08227e-08 0 2.09967e-08 0 2.09997e-08 0.0007 2.10027e-08 0 2.11767e-08 0 2.11797e-08 0.0007 2.11827e-08 0 2.13567e-08 0 2.13597e-08 0.0007 2.13627e-08 0 2.15367e-08 0 2.15397e-08 0.0007 2.15427e-08 0 2.17167e-08 0 2.17197e-08 0.0007 2.17227e-08 0 2.18967e-08 0 2.18997e-08 0.0007 2.19027e-08 0 2.20767e-08 0 2.20797e-08 0.0007 2.20827e-08 0 2.22567e-08 0 2.22597e-08 0.0007 2.22627e-08 0 2.24367e-08 0 2.24397e-08 0.0007 2.24427e-08 0 2.26167e-08 0 2.26197e-08 0.0007 2.26227e-08 0 2.27967e-08 0 2.27997e-08 0.0007 2.28027e-08 0 2.29767e-08 0 2.29797e-08 0.0007 2.29827e-08 0 3.46767e-08 0 3.46797e-08 0.0007 3.46827e-08 0 3.48567e-08 0 3.48597e-08 0.0007 3.48627e-08 0 3.50367e-08 0 3.50397e-08 0.0007 3.50427e-08 0 3.52167e-08 0 3.52197e-08 0.0007 3.52227e-08 0 3.53967e-08 0 3.53997e-08 0.0007 3.54027e-08 0 3.55767e-08 0 3.55797e-08 0.0007 3.55827e-08 0 3.57567e-08 0 3.57597e-08 0.0007 3.57627e-08 0 3.59367e-08 0 3.59397e-08 0.0007 3.59427e-08 0 3.61167e-08 0 3.61197e-08 0.0007 3.61227e-08 0 3.62967e-08 0 3.62997e-08 0.0007 3.63027e-08 0 3.64767e-08 0 3.64797e-08 0.0007 3.64827e-08 0 3.66567e-08 0 3.66597e-08 0.0007 3.66627e-08 0 3.68367e-08 0 3.68397e-08 0.0007 3.68427e-08 0 3.70167e-08 0 3.70197e-08 0.0007 3.70227e-08 0 3.71967e-08 0 3.71997e-08 0.0007 3.72027e-08 0 3.73767e-08 0 3.73797e-08 0.0007 3.73827e-08 0 3.75567e-08 0 3.75597e-08 0.0007 3.75627e-08 0 3.77367e-08 0 3.77397e-08 0.0007 3.77427e-08 0 3.79167e-08 0 3.79197e-08 0.0007 3.79227e-08 0 3.80967e-08 0 3.80997e-08 0.0007 3.81027e-08 0 3.82767e-08 0 3.82797e-08 0.0007 3.82827e-08 0 3.84567e-08 0 3.84597e-08 0.0007 3.84627e-08 0 3.86367e-08 0 3.86397e-08 0.0007 3.86427e-08 0 3.88167e-08 0 3.88197e-08 0.0007 3.88227e-08 0 3.89967e-08 0 3.89997e-08 0.0007 3.90027e-08 0 3.91767e-08 0 3.91797e-08 0.0007 3.91827e-08 0 3.93567e-08 0 3.93597e-08 0.0007 3.93627e-08 0 3.95367e-08 0 3.95397e-08 0.0007 3.95427e-08 0 3.97167e-08 0 3.97197e-08 0.0007 3.97227e-08 0 3.98967e-08 0 3.98997e-08 0.0007 3.99027e-08 0 4.00767e-08 0 4.00797e-08 0.0007 4.00827e-08 0 4.02567e-08 0 4.02597e-08 0.0007 4.02627e-08 0 4.04367e-08 0 4.04397e-08 0.0007 4.04427e-08 0 4.06167e-08 0 4.06197e-08 0.0007 4.06227e-08 0 4.07967e-08 0 4.07997e-08 0.0007 4.08027e-08 0 4.09767e-08 0 4.09797e-08 0.0007 4.09827e-08 0 4.11567e-08 0 4.11597e-08 0.0007 4.11627e-08 0 4.13367e-08 0 4.13397e-08 0.0007 4.13427e-08 0 4.15167e-08 0 4.15197e-08 0.0007 4.15227e-08 0 4.16967e-08 0 4.16997e-08 0.0007 4.17027e-08 0 4.18767e-08 0 4.18797e-08 0.0007 4.18827e-08 0 4.20567e-08 0 4.20597e-08 0.0007 4.20627e-08 0 4.22367e-08 0 4.22397e-08 0.0007 4.22427e-08 0 4.24167e-08 0 4.24197e-08 0.0007 4.24227e-08 0 4.25967e-08 0 4.25997e-08 0.0007 4.26027e-08 0 4.27767e-08 0 4.27797e-08 0.0007 4.27827e-08 0 4.29567e-08 0 4.29597e-08 0.0007 4.29627e-08 0 4.31367e-08 0 4.31397e-08 0.0007 4.31427e-08 0 4.33167e-08 0 4.33197e-08 0.0007 4.33227e-08 0 4.34967e-08 0 4.34997e-08 0.0007 4.35027e-08 0 4.36767e-08 0 4.36797e-08 0.0007 4.36827e-08 0 4.38567e-08 0 4.38597e-08 0.0007 4.38627e-08 0 4.40367e-08 0 4.40397e-08 0.0007 4.40427e-08 0 4.42167e-08 0 4.42197e-08 0.0007 4.42227e-08 0 4.43967e-08 0 4.43997e-08 0.0007 4.44027e-08 0 4.45767e-08 0 4.45797e-08 0.0007 4.45827e-08 0 4.47567e-08 0 4.47597e-08 0.0007 4.47627e-08 0 4.49367e-08 0 4.49397e-08 0.0007 4.49427e-08 0 4.51167e-08 0 4.51197e-08 0.0007 4.51227e-08 0 4.52967e-08 0 4.52997e-08 0.0007 4.53027e-08 0 4.54767e-08 0 4.54797e-08 0.0007 4.54827e-08 0 4.56567e-08 0 4.56597e-08 0.0007 4.56627e-08 0 4.58367e-08 0 4.58397e-08 0.0007 4.58427e-08 0 4.60167e-08 0 4.60197e-08 0.0007 4.60227e-08 0)
IB3|H 0 B3  PWL(0 0 2.31711e-08 0 2.31741e-08 0.0007 2.31771e-08 0 2.33511e-08 0 2.33541e-08 0.0007 2.33571e-08 0 2.35311e-08 0 2.35341e-08 0.0007 2.35371e-08 0 2.37111e-08 0 2.37141e-08 0.0007 2.37171e-08 0 2.38911e-08 0 2.38941e-08 0.0007 2.38971e-08 0 2.40711e-08 0 2.40741e-08 0.0007 2.40771e-08 0 2.42511e-08 0 2.42541e-08 0.0007 2.42571e-08 0 2.44311e-08 0 2.44341e-08 0.0007 2.44371e-08 0 2.46111e-08 0 2.46141e-08 0.0007 2.46171e-08 0 2.47911e-08 0 2.47941e-08 0.0007 2.47971e-08 0 2.49711e-08 0 2.49741e-08 0.0007 2.49771e-08 0 2.51511e-08 0 2.51541e-08 0.0007 2.51571e-08 0 2.53311e-08 0 2.53341e-08 0.0007 2.53371e-08 0 2.55111e-08 0 2.55141e-08 0.0007 2.55171e-08 0 2.56911e-08 0 2.56941e-08 0.0007 2.56971e-08 0 2.58711e-08 0 2.58741e-08 0.0007 2.58771e-08 0 2.60511e-08 0 2.60541e-08 0.0007 2.60571e-08 0 2.62311e-08 0 2.62341e-08 0.0007 2.62371e-08 0 2.64111e-08 0 2.64141e-08 0.0007 2.64171e-08 0 2.65911e-08 0 2.65941e-08 0.0007 2.65971e-08 0 2.67711e-08 0 2.67741e-08 0.0007 2.67771e-08 0 2.69511e-08 0 2.69541e-08 0.0007 2.69571e-08 0 2.71311e-08 0 2.71341e-08 0.0007 2.71371e-08 0 2.73111e-08 0 2.73141e-08 0.0007 2.73171e-08 0 2.74911e-08 0 2.74941e-08 0.0007 2.74971e-08 0 2.76711e-08 0 2.76741e-08 0.0007 2.76771e-08 0 2.78511e-08 0 2.78541e-08 0.0007 2.78571e-08 0 2.80311e-08 0 2.80341e-08 0.0007 2.80371e-08 0 2.82111e-08 0 2.82141e-08 0.0007 2.82171e-08 0 2.83911e-08 0 2.83941e-08 0.0007 2.83971e-08 0 2.85711e-08 0 2.85741e-08 0.0007 2.85771e-08 0 2.87511e-08 0 2.87541e-08 0.0007 2.87571e-08 0 2.89311e-08 0 2.89341e-08 0.0007 2.89371e-08 0 2.91111e-08 0 2.91141e-08 0.0007 2.91171e-08 0 2.92911e-08 0 2.92941e-08 0.0007 2.92971e-08 0 2.94711e-08 0 2.94741e-08 0.0007 2.94771e-08 0 2.96511e-08 0 2.96541e-08 0.0007 2.96571e-08 0 2.98311e-08 0 2.98341e-08 0.0007 2.98371e-08 0 3.00111e-08 0 3.00141e-08 0.0007 3.00171e-08 0 3.01911e-08 0 3.01941e-08 0.0007 3.01971e-08 0 3.03711e-08 0 3.03741e-08 0.0007 3.03771e-08 0 3.05511e-08 0 3.05541e-08 0.0007 3.05571e-08 0 3.07311e-08 0 3.07341e-08 0.0007 3.07371e-08 0 3.09111e-08 0 3.09141e-08 0.0007 3.09171e-08 0 3.10911e-08 0 3.10941e-08 0.0007 3.10971e-08 0 3.12711e-08 0 3.12741e-08 0.0007 3.12771e-08 0 3.14511e-08 0 3.14541e-08 0.0007 3.14571e-08 0 3.16311e-08 0 3.16341e-08 0.0007 3.16371e-08 0 3.18111e-08 0 3.18141e-08 0.0007 3.18171e-08 0 3.19911e-08 0 3.19941e-08 0.0007 3.19971e-08 0 3.21711e-08 0 3.21741e-08 0.0007 3.21771e-08 0 3.23511e-08 0 3.23541e-08 0.0007 3.23571e-08 0 3.25311e-08 0 3.25341e-08 0.0007 3.25371e-08 0 3.27111e-08 0 3.27141e-08 0.0007 3.27171e-08 0 3.28911e-08 0 3.28941e-08 0.0007 3.28971e-08 0 3.30711e-08 0 3.30741e-08 0.0007 3.30771e-08 0 3.32511e-08 0 3.32541e-08 0.0007 3.32571e-08 0 3.34311e-08 0 3.34341e-08 0.0007 3.34371e-08 0 3.36111e-08 0 3.36141e-08 0.0007 3.36171e-08 0 3.37911e-08 0 3.37941e-08 0.0007 3.37971e-08 0 3.39711e-08 0 3.39741e-08 0.0007 3.39771e-08 0 3.41511e-08 0 3.41541e-08 0.0007 3.41571e-08 0 3.43311e-08 0 3.43341e-08 0.0007 3.43371e-08 0 3.45111e-08 0 3.45141e-08 0.0007 3.45171e-08 0 3.46911e-08 0 3.46941e-08 0.0007 3.46971e-08 0 3.48711e-08 0 3.48741e-08 0.0007 3.48771e-08 0 3.50511e-08 0 3.50541e-08 0.0007 3.50571e-08 0 3.52311e-08 0 3.52341e-08 0.0007 3.52371e-08 0 3.54111e-08 0 3.54141e-08 0.0007 3.54171e-08 0 3.55911e-08 0 3.55941e-08 0.0007 3.55971e-08 0 3.57711e-08 0 3.57741e-08 0.0007 3.57771e-08 0 3.59511e-08 0 3.59541e-08 0.0007 3.59571e-08 0 3.61311e-08 0 3.61341e-08 0.0007 3.61371e-08 0 3.63111e-08 0 3.63141e-08 0.0007 3.63171e-08 0 3.64911e-08 0 3.64941e-08 0.0007 3.64971e-08 0 3.66711e-08 0 3.66741e-08 0.0007 3.66771e-08 0 3.68511e-08 0 3.68541e-08 0.0007 3.68571e-08 0 3.70311e-08 0 3.70341e-08 0.0007 3.70371e-08 0 3.72111e-08 0 3.72141e-08 0.0007 3.72171e-08 0 3.73911e-08 0 3.73941e-08 0.0007 3.73971e-08 0 3.75711e-08 0 3.75741e-08 0.0007 3.75771e-08 0 3.77511e-08 0 3.77541e-08 0.0007 3.77571e-08 0 3.79311e-08 0 3.79341e-08 0.0007 3.79371e-08 0 3.81111e-08 0 3.81141e-08 0.0007 3.81171e-08 0 3.82911e-08 0 3.82941e-08 0.0007 3.82971e-08 0 3.84711e-08 0 3.84741e-08 0.0007 3.84771e-08 0 3.86511e-08 0 3.86541e-08 0.0007 3.86571e-08 0 3.88311e-08 0 3.88341e-08 0.0007 3.88371e-08 0 3.90111e-08 0 3.90141e-08 0.0007 3.90171e-08 0 3.91911e-08 0 3.91941e-08 0.0007 3.91971e-08 0 3.93711e-08 0 3.93741e-08 0.0007 3.93771e-08 0 3.95511e-08 0 3.95541e-08 0.0007 3.95571e-08 0 3.97311e-08 0 3.97341e-08 0.0007 3.97371e-08 0 3.99111e-08 0 3.99141e-08 0.0007 3.99171e-08 0 4.00911e-08 0 4.00941e-08 0.0007 4.00971e-08 0 4.02711e-08 0 4.02741e-08 0.0007 4.02771e-08 0 4.04511e-08 0 4.04541e-08 0.0007 4.04571e-08 0 4.06311e-08 0 4.06341e-08 0.0007 4.06371e-08 0 4.08111e-08 0 4.08141e-08 0.0007 4.08171e-08 0 4.09911e-08 0 4.09941e-08 0.0007 4.09971e-08 0 4.11711e-08 0 4.11741e-08 0.0007 4.11771e-08 0 4.13511e-08 0 4.13541e-08 0.0007 4.13571e-08 0 4.15311e-08 0 4.15341e-08 0.0007 4.15371e-08 0 4.17111e-08 0 4.17141e-08 0.0007 4.17171e-08 0 4.18911e-08 0 4.18941e-08 0.0007 4.18971e-08 0 4.20711e-08 0 4.20741e-08 0.0007 4.20771e-08 0 4.22511e-08 0 4.22541e-08 0.0007 4.22571e-08 0 4.24311e-08 0 4.24341e-08 0.0007 4.24371e-08 0 4.26111e-08 0 4.26141e-08 0.0007 4.26171e-08 0 4.27911e-08 0 4.27941e-08 0.0007 4.27971e-08 0 4.29711e-08 0 4.29741e-08 0.0007 4.29771e-08 0 4.31511e-08 0 4.31541e-08 0.0007 4.31571e-08 0 4.33311e-08 0 4.33341e-08 0.0007 4.33371e-08 0 4.35111e-08 0 4.35141e-08 0.0007 4.35171e-08 0 4.36911e-08 0 4.36941e-08 0.0007 4.36971e-08 0 4.38711e-08 0 4.38741e-08 0.0007 4.38771e-08 0 4.40511e-08 0 4.40541e-08 0.0007 4.40571e-08 0 4.42311e-08 0 4.42341e-08 0.0007 4.42371e-08 0 4.44111e-08 0 4.44141e-08 0.0007 4.44171e-08 0 4.45911e-08 0 4.45941e-08 0.0007 4.45971e-08 0 4.47711e-08 0 4.47741e-08 0.0007 4.47771e-08 0 4.49511e-08 0 4.49541e-08 0.0007 4.49571e-08 0 4.51311e-08 0 4.51341e-08 0.0007 4.51371e-08 0 4.53111e-08 0 4.53141e-08 0.0007 4.53171e-08 0 4.54911e-08 0 4.54941e-08 0.0007 4.54971e-08 0 4.56711e-08 0 4.56741e-08 0.0007 4.56771e-08 0 4.58511e-08 0 4.58541e-08 0.0007 4.58571e-08 0 4.60311e-08 0 4.60341e-08 0.0007 4.60371e-08 0)
IT00|T 0 T00  PWL(0 0 1.5e-11 0 1.8e-11 0.0021 2.1e-11 0 1.95e-10 0 1.98e-10 0.0021 2.01e-10 0 3.75e-10 0 3.78e-10 0.0021 3.81e-10 0 5.55e-10 0 5.58e-10 0.0021 5.61e-10 0 7.35e-10 0 7.38e-10 0.0021 7.41e-10 0 9.15e-10 0 9.18e-10 0.0021 9.21e-10 0 1.095e-09 0 1.098e-09 0.0021 1.101e-09 0 1.275e-09 0 1.278e-09 0.0021 1.281e-09 0 1.455e-09 0 1.458e-09 0.0021 1.461e-09 0 1.635e-09 0 1.638e-09 0.0021 1.641e-09 0 1.815e-09 0 1.818e-09 0.0021 1.821e-09 0 1.995e-09 0 1.998e-09 0.0021 2.001e-09 0 2.175e-09 0 2.178e-09 0.0021 2.181e-09 0 2.355e-09 0 2.358e-09 0.0021 2.361e-09 0 2.535e-09 0 2.538e-09 0.0021 2.541e-09 0 2.715e-09 0 2.718e-09 0.0021 2.721e-09 0 2.895e-09 0 2.898e-09 0.0021 2.901e-09 0 3.075e-09 0 3.078e-09 0.0021 3.081e-09 0 3.255e-09 0 3.258e-09 0.0021 3.261e-09 0 3.435e-09 0 3.438e-09 0.0021 3.441e-09 0 3.615e-09 0 3.618e-09 0.0021 3.621e-09 0 3.795e-09 0 3.798e-09 0.0021 3.801e-09 0 3.975e-09 0 3.978e-09 0.0021 3.981e-09 0 4.155e-09 0 4.158e-09 0.0021 4.161e-09 0 4.335e-09 0 4.338e-09 0.0021 4.341e-09 0 4.515e-09 0 4.518e-09 0.0021 4.521e-09 0 4.695e-09 0 4.698e-09 0.0021 4.701e-09 0 4.875e-09 0 4.878e-09 0.0021 4.881e-09 0 5.055e-09 0 5.058e-09 0.0021 5.061e-09 0 5.235e-09 0 5.238e-09 0.0021 5.241e-09 0 5.415e-09 0 5.418e-09 0.0021 5.421e-09 0 5.595e-09 0 5.598e-09 0.0021 5.601e-09 0 5.775e-09 0 5.778e-09 0.0021 5.781e-09 0 5.955e-09 0 5.958e-09 0.0021 5.961e-09 0 6.135e-09 0 6.138e-09 0.0021 6.141e-09 0 6.315e-09 0 6.318e-09 0.0021 6.321e-09 0 6.495e-09 0 6.498e-09 0.0021 6.501e-09 0 6.675e-09 0 6.678e-09 0.0021 6.681e-09 0 6.855e-09 0 6.858e-09 0.0021 6.861e-09 0 7.035e-09 0 7.038e-09 0.0021 7.041e-09 0 7.215e-09 0 7.218e-09 0.0021 7.221e-09 0 7.395e-09 0 7.398e-09 0.0021 7.401e-09 0 7.575e-09 0 7.578e-09 0.0021 7.581e-09 0 7.755e-09 0 7.758e-09 0.0021 7.761e-09 0 7.935e-09 0 7.938e-09 0.0021 7.941e-09 0 8.115e-09 0 8.118e-09 0.0021 8.121e-09 0 8.295e-09 0 8.298e-09 0.0021 8.301e-09 0 8.475e-09 0 8.478e-09 0.0021 8.481e-09 0 8.655e-09 0 8.658e-09 0.0021 8.661e-09 0 8.835e-09 0 8.838e-09 0.0021 8.841e-09 0 9.015e-09 0 9.018e-09 0.0021 9.021e-09 0 9.195e-09 0 9.198e-09 0.0021 9.201e-09 0 9.375e-09 0 9.378e-09 0.0021 9.381e-09 0 9.555e-09 0 9.558e-09 0.0021 9.561e-09 0 9.735e-09 0 9.738e-09 0.0021 9.741e-09 0 9.915e-09 0 9.918e-09 0.0021 9.921e-09 0 1.0095e-08 0 1.0098e-08 0.0021 1.0101e-08 0 1.0275e-08 0 1.0278e-08 0.0021 1.0281e-08 0 1.0455e-08 0 1.0458e-08 0.0021 1.0461e-08 0 1.0635e-08 0 1.0638e-08 0.0021 1.0641e-08 0 1.0815e-08 0 1.0818e-08 0.0021 1.0821e-08 0 1.0995e-08 0 1.0998e-08 0.0021 1.1001e-08 0 1.1175e-08 0 1.1178e-08 0.0021 1.1181e-08 0 1.1355e-08 0 1.1358e-08 0.0021 1.1361e-08 0 1.1535e-08 0 1.1538e-08 0.0021 1.1541e-08 0 1.1715e-08 0 1.1718e-08 0.0021 1.1721e-08 0 1.1895e-08 0 1.1898e-08 0.0021 1.1901e-08 0 1.2075e-08 0 1.2078e-08 0.0021 1.2081e-08 0 1.2255e-08 0 1.2258e-08 0.0021 1.2261e-08 0 1.2435e-08 0 1.2438e-08 0.0021 1.2441e-08 0 1.2615e-08 0 1.2618e-08 0.0021 1.2621e-08 0 1.2795e-08 0 1.2798e-08 0.0021 1.2801e-08 0 1.2975e-08 0 1.2978e-08 0.0021 1.2981e-08 0 1.3155e-08 0 1.3158e-08 0.0021 1.3161e-08 0 1.3335e-08 0 1.3338e-08 0.0021 1.3341e-08 0 1.3515e-08 0 1.3518e-08 0.0021 1.3521e-08 0 1.3695e-08 0 1.3698e-08 0.0021 1.3701e-08 0 1.3875e-08 0 1.3878e-08 0.0021 1.3881e-08 0 1.4055e-08 0 1.4058e-08 0.0021 1.4061e-08 0 1.4235e-08 0 1.4238e-08 0.0021 1.4241e-08 0 1.4415e-08 0 1.4418e-08 0.0021 1.4421e-08 0 1.4595e-08 0 1.4598e-08 0.0021 1.4601e-08 0 1.4775e-08 0 1.4778e-08 0.0021 1.4781e-08 0 1.4955e-08 0 1.4958e-08 0.0021 1.4961e-08 0 1.5135e-08 0 1.5138e-08 0.0021 1.5141e-08 0 1.5315e-08 0 1.5318e-08 0.0021 1.5321e-08 0 1.5495e-08 0 1.5498e-08 0.0021 1.5501e-08 0 1.5675e-08 0 1.5678e-08 0.0021 1.5681e-08 0 1.5855e-08 0 1.5858e-08 0.0021 1.5861e-08 0 1.6035e-08 0 1.6038e-08 0.0021 1.6041e-08 0 1.6215e-08 0 1.6218e-08 0.0021 1.6221e-08 0 1.6395e-08 0 1.6398e-08 0.0021 1.6401e-08 0 1.6575e-08 0 1.6578e-08 0.0021 1.6581e-08 0 1.6755e-08 0 1.6758e-08 0.0021 1.6761e-08 0 1.6935e-08 0 1.6938e-08 0.0021 1.6941e-08 0 1.7115e-08 0 1.7118e-08 0.0021 1.7121e-08 0 1.7295e-08 0 1.7298e-08 0.0021 1.7301e-08 0 1.7475e-08 0 1.7478e-08 0.0021 1.7481e-08 0 1.7655e-08 0 1.7658e-08 0.0021 1.7661e-08 0 1.7835e-08 0 1.7838e-08 0.0021 1.7841e-08 0 1.8015e-08 0 1.8018e-08 0.0021 1.8021e-08 0 1.8195e-08 0 1.8198e-08 0.0021 1.8201e-08 0 1.8375e-08 0 1.8378e-08 0.0021 1.8381e-08 0 1.8555e-08 0 1.8558e-08 0.0021 1.8561e-08 0 1.8735e-08 0 1.8738e-08 0.0021 1.8741e-08 0 1.8915e-08 0 1.8918e-08 0.0021 1.8921e-08 0 1.9095e-08 0 1.9098e-08 0.0021 1.9101e-08 0 1.9275e-08 0 1.9278e-08 0.0021 1.9281e-08 0 1.9455e-08 0 1.9458e-08 0.0021 1.9461e-08 0 1.9635e-08 0 1.9638e-08 0.0021 1.9641e-08 0 1.9815e-08 0 1.9818e-08 0.0021 1.9821e-08 0 1.9995e-08 0 1.9998e-08 0.0021 2.0001e-08 0 2.0175e-08 0 2.0178e-08 0.0021 2.0181e-08 0 2.0355e-08 0 2.0358e-08 0.0021 2.0361e-08 0 2.0535e-08 0 2.0538e-08 0.0021 2.0541e-08 0 2.0715e-08 0 2.0718e-08 0.0021 2.0721e-08 0 2.0895e-08 0 2.0898e-08 0.0021 2.0901e-08 0 2.1075e-08 0 2.1078e-08 0.0021 2.1081e-08 0 2.1255e-08 0 2.1258e-08 0.0021 2.1261e-08 0 2.1435e-08 0 2.1438e-08 0.0021 2.1441e-08 0 2.1615e-08 0 2.1618e-08 0.0021 2.1621e-08 0 2.1795e-08 0 2.1798e-08 0.0021 2.1801e-08 0 2.1975e-08 0 2.1978e-08 0.0021 2.1981e-08 0 2.2155e-08 0 2.2158e-08 0.0021 2.2161e-08 0 2.2335e-08 0 2.2338e-08 0.0021 2.2341e-08 0 2.2515e-08 0 2.2518e-08 0.0021 2.2521e-08 0 2.2695e-08 0 2.2698e-08 0.0021 2.2701e-08 0 2.2875e-08 0 2.2878e-08 0.0021 2.2881e-08 0 2.3055e-08 0 2.3058e-08 0.0021 2.3061e-08 0 2.3235e-08 0 2.3238e-08 0.0021 2.3241e-08 0 2.3415e-08 0 2.3418e-08 0.0021 2.3421e-08 0 2.3595e-08 0 2.3598e-08 0.0021 2.3601e-08 0 2.3775e-08 0 2.3778e-08 0.0021 2.3781e-08 0 2.3955e-08 0 2.3958e-08 0.0021 2.3961e-08 0 2.4135e-08 0 2.4138e-08 0.0021 2.4141e-08 0 2.4315e-08 0 2.4318e-08 0.0021 2.4321e-08 0 2.4495e-08 0 2.4498e-08 0.0021 2.4501e-08 0 2.4675e-08 0 2.4678e-08 0.0021 2.4681e-08 0 2.4855e-08 0 2.4858e-08 0.0021 2.4861e-08 0 2.5035e-08 0 2.5038e-08 0.0021 2.5041e-08 0 2.5215e-08 0 2.5218e-08 0.0021 2.5221e-08 0 2.5395e-08 0 2.5398e-08 0.0021 2.5401e-08 0 2.5575e-08 0 2.5578e-08 0.0021 2.5581e-08 0 2.5755e-08 0 2.5758e-08 0.0021 2.5761e-08 0 2.5935e-08 0 2.5938e-08 0.0021 2.5941e-08 0 2.6115e-08 0 2.6118e-08 0.0021 2.6121e-08 0 2.6295e-08 0 2.6298e-08 0.0021 2.6301e-08 0 2.6475e-08 0 2.6478e-08 0.0021 2.6481e-08 0 2.6655e-08 0 2.6658e-08 0.0021 2.6661e-08 0 2.6835e-08 0 2.6838e-08 0.0021 2.6841e-08 0 2.7015e-08 0 2.7018e-08 0.0021 2.7021e-08 0 2.7195e-08 0 2.7198e-08 0.0021 2.7201e-08 0 2.7375e-08 0 2.7378e-08 0.0021 2.7381e-08 0 2.7555e-08 0 2.7558e-08 0.0021 2.7561e-08 0 2.7735e-08 0 2.7738e-08 0.0021 2.7741e-08 0 2.7915e-08 0 2.7918e-08 0.0021 2.7921e-08 0 2.8095e-08 0 2.8098e-08 0.0021 2.8101e-08 0 2.8275e-08 0 2.8278e-08 0.0021 2.8281e-08 0 2.8455e-08 0 2.8458e-08 0.0021 2.8461e-08 0 2.8635e-08 0 2.8638e-08 0.0021 2.8641e-08 0 2.8815e-08 0 2.8818e-08 0.0021 2.8821e-08 0 2.8995e-08 0 2.8998e-08 0.0021 2.9001e-08 0 2.9175e-08 0 2.9178e-08 0.0021 2.9181e-08 0 2.9355e-08 0 2.9358e-08 0.0021 2.9361e-08 0 2.9535e-08 0 2.9538e-08 0.0021 2.9541e-08 0 2.9715e-08 0 2.9718e-08 0.0021 2.9721e-08 0 2.9895e-08 0 2.9898e-08 0.0021 2.9901e-08 0 3.0075e-08 0 3.0078e-08 0.0021 3.0081e-08 0 3.0255e-08 0 3.0258e-08 0.0021 3.0261e-08 0 3.0435e-08 0 3.0438e-08 0.0021 3.0441e-08 0 3.0615e-08 0 3.0618e-08 0.0021 3.0621e-08 0 3.0795e-08 0 3.0798e-08 0.0021 3.0801e-08 0 3.0975e-08 0 3.0978e-08 0.0021 3.0981e-08 0 3.1155e-08 0 3.1158e-08 0.0021 3.1161e-08 0 3.1335e-08 0 3.1338e-08 0.0021 3.1341e-08 0 3.1515e-08 0 3.1518e-08 0.0021 3.1521e-08 0 3.1695e-08 0 3.1698e-08 0.0021 3.1701e-08 0 3.1875e-08 0 3.1878e-08 0.0021 3.1881e-08 0 3.2055e-08 0 3.2058e-08 0.0021 3.2061e-08 0 3.2235e-08 0 3.2238e-08 0.0021 3.2241e-08 0 3.2415e-08 0 3.2418e-08 0.0021 3.2421e-08 0 3.2595e-08 0 3.2598e-08 0.0021 3.2601e-08 0 3.2775e-08 0 3.2778e-08 0.0021 3.2781e-08 0 3.2955e-08 0 3.2958e-08 0.0021 3.2961e-08 0 3.3135e-08 0 3.3138e-08 0.0021 3.3141e-08 0 3.3315e-08 0 3.3318e-08 0.0021 3.3321e-08 0 3.3495e-08 0 3.3498e-08 0.0021 3.3501e-08 0 3.3675e-08 0 3.3678e-08 0.0021 3.3681e-08 0 3.3855e-08 0 3.3858e-08 0.0021 3.3861e-08 0 3.4035e-08 0 3.4038e-08 0.0021 3.4041e-08 0 3.4215e-08 0 3.4218e-08 0.0021 3.4221e-08 0 3.4395e-08 0 3.4398e-08 0.0021 3.4401e-08 0 3.4575e-08 0 3.4578e-08 0.0021 3.4581e-08 0 3.4755e-08 0 3.4758e-08 0.0021 3.4761e-08 0 3.4935e-08 0 3.4938e-08 0.0021 3.4941e-08 0 3.5115e-08 0 3.5118e-08 0.0021 3.5121e-08 0 3.5295e-08 0 3.5298e-08 0.0021 3.5301e-08 0 3.5475e-08 0 3.5478e-08 0.0021 3.5481e-08 0 3.5655e-08 0 3.5658e-08 0.0021 3.5661e-08 0 3.5835e-08 0 3.5838e-08 0.0021 3.5841e-08 0 3.6015e-08 0 3.6018e-08 0.0021 3.6021e-08 0 3.6195e-08 0 3.6198e-08 0.0021 3.6201e-08 0 3.6375e-08 0 3.6378e-08 0.0021 3.6381e-08 0 3.6555e-08 0 3.6558e-08 0.0021 3.6561e-08 0 3.6735e-08 0 3.6738e-08 0.0021 3.6741e-08 0 3.6915e-08 0 3.6918e-08 0.0021 3.6921e-08 0 3.7095e-08 0 3.7098e-08 0.0021 3.7101e-08 0 3.7275e-08 0 3.7278e-08 0.0021 3.7281e-08 0 3.7455e-08 0 3.7458e-08 0.0021 3.7461e-08 0 3.7635e-08 0 3.7638e-08 0.0021 3.7641e-08 0 3.7815e-08 0 3.7818e-08 0.0021 3.7821e-08 0 3.7995e-08 0 3.7998e-08 0.0021 3.8001e-08 0 3.8175e-08 0 3.8178e-08 0.0021 3.8181e-08 0 3.8355e-08 0 3.8358e-08 0.0021 3.8361e-08 0 3.8535e-08 0 3.8538e-08 0.0021 3.8541e-08 0 3.8715e-08 0 3.8718e-08 0.0021 3.8721e-08 0 3.8895e-08 0 3.8898e-08 0.0021 3.8901e-08 0 3.9075e-08 0 3.9078e-08 0.0021 3.9081e-08 0 3.9255e-08 0 3.9258e-08 0.0021 3.9261e-08 0 3.9435e-08 0 3.9438e-08 0.0021 3.9441e-08 0 3.9615e-08 0 3.9618e-08 0.0021 3.9621e-08 0 3.9795e-08 0 3.9798e-08 0.0021 3.9801e-08 0 3.9975e-08 0 3.9978e-08 0.0021 3.9981e-08 0 4.0155e-08 0 4.0158e-08 0.0021 4.0161e-08 0 4.0335e-08 0 4.0338e-08 0.0021 4.0341e-08 0 4.0515e-08 0 4.0518e-08 0.0021 4.0521e-08 0 4.0695e-08 0 4.0698e-08 0.0021 4.0701e-08 0 4.0875e-08 0 4.0878e-08 0.0021 4.0881e-08 0 4.1055e-08 0 4.1058e-08 0.0021 4.1061e-08 0 4.1235e-08 0 4.1238e-08 0.0021 4.1241e-08 0 4.1415e-08 0 4.1418e-08 0.0021 4.1421e-08 0 4.1595e-08 0 4.1598e-08 0.0021 4.1601e-08 0 4.1775e-08 0 4.1778e-08 0.0021 4.1781e-08 0 4.1955e-08 0 4.1958e-08 0.0021 4.1961e-08 0 4.2135e-08 0 4.2138e-08 0.0021 4.2141e-08 0 4.2315e-08 0 4.2318e-08 0.0021 4.2321e-08 0 4.2495e-08 0 4.2498e-08 0.0021 4.2501e-08 0 4.2675e-08 0 4.2678e-08 0.0021 4.2681e-08 0 4.2855e-08 0 4.2858e-08 0.0021 4.2861e-08 0 4.3035e-08 0 4.3038e-08 0.0021 4.3041e-08 0 4.3215e-08 0 4.3218e-08 0.0021 4.3221e-08 0 4.3395e-08 0 4.3398e-08 0.0021 4.3401e-08 0 4.3575e-08 0 4.3578e-08 0.0021 4.3581e-08 0 4.3755e-08 0 4.3758e-08 0.0021 4.3761e-08 0 4.3935e-08 0 4.3938e-08 0.0021 4.3941e-08 0 4.4115e-08 0 4.4118e-08 0.0021 4.4121e-08 0 4.4295e-08 0 4.4298e-08 0.0021 4.4301e-08 0 4.4475e-08 0 4.4478e-08 0.0021 4.4481e-08 0 4.4655e-08 0 4.4658e-08 0.0021 4.4661e-08 0 4.4835e-08 0 4.4838e-08 0.0021 4.4841e-08 0 4.5015e-08 0 4.5018e-08 0.0021 4.5021e-08 0 4.5195e-08 0 4.5198e-08 0.0021 4.5201e-08 0 4.5375e-08 0 4.5378e-08 0.0021 4.5381e-08 0 4.5555e-08 0 4.5558e-08 0.0021 4.5561e-08 0 4.5735e-08 0 4.5738e-08 0.0021 4.5741e-08 0 4.5915e-08 0 4.5918e-08 0.0021 4.5921e-08 0)
IT01|T 0 T01  PWL(0 0 1.5e-11 0 1.8e-11 0.0021 2.1e-11 0 1.95e-10 0 1.98e-10 0.0021 2.01e-10 0 3.75e-10 0 3.78e-10 0.0021 3.81e-10 0 5.55e-10 0 5.58e-10 0.0021 5.61e-10 0 7.35e-10 0 7.38e-10 0.0021 7.41e-10 0 9.15e-10 0 9.18e-10 0.0021 9.21e-10 0 1.095e-09 0 1.098e-09 0.0021 1.101e-09 0 1.275e-09 0 1.278e-09 0.0021 1.281e-09 0 1.455e-09 0 1.458e-09 0.0021 1.461e-09 0 1.635e-09 0 1.638e-09 0.0021 1.641e-09 0 1.815e-09 0 1.818e-09 0.0021 1.821e-09 0 1.995e-09 0 1.998e-09 0.0021 2.001e-09 0 2.175e-09 0 2.178e-09 0.0021 2.181e-09 0 2.355e-09 0 2.358e-09 0.0021 2.361e-09 0 2.535e-09 0 2.538e-09 0.0021 2.541e-09 0 2.715e-09 0 2.718e-09 0.0021 2.721e-09 0 2.895e-09 0 2.898e-09 0.0021 2.901e-09 0 3.075e-09 0 3.078e-09 0.0021 3.081e-09 0 3.255e-09 0 3.258e-09 0.0021 3.261e-09 0 3.435e-09 0 3.438e-09 0.0021 3.441e-09 0 3.615e-09 0 3.618e-09 0.0021 3.621e-09 0 3.795e-09 0 3.798e-09 0.0021 3.801e-09 0 3.975e-09 0 3.978e-09 0.0021 3.981e-09 0 4.155e-09 0 4.158e-09 0.0021 4.161e-09 0 4.335e-09 0 4.338e-09 0.0021 4.341e-09 0 4.515e-09 0 4.518e-09 0.0021 4.521e-09 0 4.695e-09 0 4.698e-09 0.0021 4.701e-09 0 4.875e-09 0 4.878e-09 0.0021 4.881e-09 0 5.055e-09 0 5.058e-09 0.0021 5.061e-09 0 5.235e-09 0 5.238e-09 0.0021 5.241e-09 0 5.415e-09 0 5.418e-09 0.0021 5.421e-09 0 5.595e-09 0 5.598e-09 0.0021 5.601e-09 0 5.775e-09 0 5.778e-09 0.0021 5.781e-09 0 5.955e-09 0 5.958e-09 0.0021 5.961e-09 0 6.135e-09 0 6.138e-09 0.0021 6.141e-09 0 6.315e-09 0 6.318e-09 0.0021 6.321e-09 0 6.495e-09 0 6.498e-09 0.0021 6.501e-09 0 6.675e-09 0 6.678e-09 0.0021 6.681e-09 0 6.855e-09 0 6.858e-09 0.0021 6.861e-09 0 7.035e-09 0 7.038e-09 0.0021 7.041e-09 0 7.215e-09 0 7.218e-09 0.0021 7.221e-09 0 7.395e-09 0 7.398e-09 0.0021 7.401e-09 0 7.575e-09 0 7.578e-09 0.0021 7.581e-09 0 7.755e-09 0 7.758e-09 0.0021 7.761e-09 0 7.935e-09 0 7.938e-09 0.0021 7.941e-09 0 8.115e-09 0 8.118e-09 0.0021 8.121e-09 0 8.295e-09 0 8.298e-09 0.0021 8.301e-09 0 8.475e-09 0 8.478e-09 0.0021 8.481e-09 0 8.655e-09 0 8.658e-09 0.0021 8.661e-09 0 8.835e-09 0 8.838e-09 0.0021 8.841e-09 0 9.015e-09 0 9.018e-09 0.0021 9.021e-09 0 9.195e-09 0 9.198e-09 0.0021 9.201e-09 0 9.375e-09 0 9.378e-09 0.0021 9.381e-09 0 9.555e-09 0 9.558e-09 0.0021 9.561e-09 0 9.735e-09 0 9.738e-09 0.0021 9.741e-09 0 9.915e-09 0 9.918e-09 0.0021 9.921e-09 0 1.0095e-08 0 1.0098e-08 0.0021 1.0101e-08 0 1.0275e-08 0 1.0278e-08 0.0021 1.0281e-08 0 1.0455e-08 0 1.0458e-08 0.0021 1.0461e-08 0 1.0635e-08 0 1.0638e-08 0.0021 1.0641e-08 0 1.0815e-08 0 1.0818e-08 0.0021 1.0821e-08 0 1.0995e-08 0 1.0998e-08 0.0021 1.1001e-08 0 1.1175e-08 0 1.1178e-08 0.0021 1.1181e-08 0 1.1355e-08 0 1.1358e-08 0.0021 1.1361e-08 0 1.1535e-08 0 1.1538e-08 0.0021 1.1541e-08 0 1.1715e-08 0 1.1718e-08 0.0021 1.1721e-08 0 1.1895e-08 0 1.1898e-08 0.0021 1.1901e-08 0 1.2075e-08 0 1.2078e-08 0.0021 1.2081e-08 0 1.2255e-08 0 1.2258e-08 0.0021 1.2261e-08 0 1.2435e-08 0 1.2438e-08 0.0021 1.2441e-08 0 1.2615e-08 0 1.2618e-08 0.0021 1.2621e-08 0 1.2795e-08 0 1.2798e-08 0.0021 1.2801e-08 0 1.2975e-08 0 1.2978e-08 0.0021 1.2981e-08 0 1.3155e-08 0 1.3158e-08 0.0021 1.3161e-08 0 1.3335e-08 0 1.3338e-08 0.0021 1.3341e-08 0 1.3515e-08 0 1.3518e-08 0.0021 1.3521e-08 0 1.3695e-08 0 1.3698e-08 0.0021 1.3701e-08 0 1.3875e-08 0 1.3878e-08 0.0021 1.3881e-08 0 1.4055e-08 0 1.4058e-08 0.0021 1.4061e-08 0 1.4235e-08 0 1.4238e-08 0.0021 1.4241e-08 0 1.4415e-08 0 1.4418e-08 0.0021 1.4421e-08 0 1.4595e-08 0 1.4598e-08 0.0021 1.4601e-08 0 1.4775e-08 0 1.4778e-08 0.0021 1.4781e-08 0 1.4955e-08 0 1.4958e-08 0.0021 1.4961e-08 0 1.5135e-08 0 1.5138e-08 0.0021 1.5141e-08 0 1.5315e-08 0 1.5318e-08 0.0021 1.5321e-08 0 1.5495e-08 0 1.5498e-08 0.0021 1.5501e-08 0 1.5675e-08 0 1.5678e-08 0.0021 1.5681e-08 0 1.5855e-08 0 1.5858e-08 0.0021 1.5861e-08 0 1.6035e-08 0 1.6038e-08 0.0021 1.6041e-08 0 1.6215e-08 0 1.6218e-08 0.0021 1.6221e-08 0 1.6395e-08 0 1.6398e-08 0.0021 1.6401e-08 0 1.6575e-08 0 1.6578e-08 0.0021 1.6581e-08 0 1.6755e-08 0 1.6758e-08 0.0021 1.6761e-08 0 1.6935e-08 0 1.6938e-08 0.0021 1.6941e-08 0 1.7115e-08 0 1.7118e-08 0.0021 1.7121e-08 0 1.7295e-08 0 1.7298e-08 0.0021 1.7301e-08 0 1.7475e-08 0 1.7478e-08 0.0021 1.7481e-08 0 1.7655e-08 0 1.7658e-08 0.0021 1.7661e-08 0 1.7835e-08 0 1.7838e-08 0.0021 1.7841e-08 0 1.8015e-08 0 1.8018e-08 0.0021 1.8021e-08 0 1.8195e-08 0 1.8198e-08 0.0021 1.8201e-08 0 1.8375e-08 0 1.8378e-08 0.0021 1.8381e-08 0 1.8555e-08 0 1.8558e-08 0.0021 1.8561e-08 0 1.8735e-08 0 1.8738e-08 0.0021 1.8741e-08 0 1.8915e-08 0 1.8918e-08 0.0021 1.8921e-08 0 1.9095e-08 0 1.9098e-08 0.0021 1.9101e-08 0 1.9275e-08 0 1.9278e-08 0.0021 1.9281e-08 0 1.9455e-08 0 1.9458e-08 0.0021 1.9461e-08 0 1.9635e-08 0 1.9638e-08 0.0021 1.9641e-08 0 1.9815e-08 0 1.9818e-08 0.0021 1.9821e-08 0 1.9995e-08 0 1.9998e-08 0.0021 2.0001e-08 0 2.0175e-08 0 2.0178e-08 0.0021 2.0181e-08 0 2.0355e-08 0 2.0358e-08 0.0021 2.0361e-08 0 2.0535e-08 0 2.0538e-08 0.0021 2.0541e-08 0 2.0715e-08 0 2.0718e-08 0.0021 2.0721e-08 0 2.0895e-08 0 2.0898e-08 0.0021 2.0901e-08 0 2.1075e-08 0 2.1078e-08 0.0021 2.1081e-08 0 2.1255e-08 0 2.1258e-08 0.0021 2.1261e-08 0 2.1435e-08 0 2.1438e-08 0.0021 2.1441e-08 0 2.1615e-08 0 2.1618e-08 0.0021 2.1621e-08 0 2.1795e-08 0 2.1798e-08 0.0021 2.1801e-08 0 2.1975e-08 0 2.1978e-08 0.0021 2.1981e-08 0 2.2155e-08 0 2.2158e-08 0.0021 2.2161e-08 0 2.2335e-08 0 2.2338e-08 0.0021 2.2341e-08 0 2.2515e-08 0 2.2518e-08 0.0021 2.2521e-08 0 2.2695e-08 0 2.2698e-08 0.0021 2.2701e-08 0 2.2875e-08 0 2.2878e-08 0.0021 2.2881e-08 0 2.3055e-08 0 2.3058e-08 0.0021 2.3061e-08 0 2.3235e-08 0 2.3238e-08 0.0021 2.3241e-08 0 2.3415e-08 0 2.3418e-08 0.0021 2.3421e-08 0 2.3595e-08 0 2.3598e-08 0.0021 2.3601e-08 0 2.3775e-08 0 2.3778e-08 0.0021 2.3781e-08 0 2.3955e-08 0 2.3958e-08 0.0021 2.3961e-08 0 2.4135e-08 0 2.4138e-08 0.0021 2.4141e-08 0 2.4315e-08 0 2.4318e-08 0.0021 2.4321e-08 0 2.4495e-08 0 2.4498e-08 0.0021 2.4501e-08 0 2.4675e-08 0 2.4678e-08 0.0021 2.4681e-08 0 2.4855e-08 0 2.4858e-08 0.0021 2.4861e-08 0 2.5035e-08 0 2.5038e-08 0.0021 2.5041e-08 0 2.5215e-08 0 2.5218e-08 0.0021 2.5221e-08 0 2.5395e-08 0 2.5398e-08 0.0021 2.5401e-08 0 2.5575e-08 0 2.5578e-08 0.0021 2.5581e-08 0 2.5755e-08 0 2.5758e-08 0.0021 2.5761e-08 0 2.5935e-08 0 2.5938e-08 0.0021 2.5941e-08 0 2.6115e-08 0 2.6118e-08 0.0021 2.6121e-08 0 2.6295e-08 0 2.6298e-08 0.0021 2.6301e-08 0 2.6475e-08 0 2.6478e-08 0.0021 2.6481e-08 0 2.6655e-08 0 2.6658e-08 0.0021 2.6661e-08 0 2.6835e-08 0 2.6838e-08 0.0021 2.6841e-08 0 2.7015e-08 0 2.7018e-08 0.0021 2.7021e-08 0 2.7195e-08 0 2.7198e-08 0.0021 2.7201e-08 0 2.7375e-08 0 2.7378e-08 0.0021 2.7381e-08 0 2.7555e-08 0 2.7558e-08 0.0021 2.7561e-08 0 2.7735e-08 0 2.7738e-08 0.0021 2.7741e-08 0 2.7915e-08 0 2.7918e-08 0.0021 2.7921e-08 0 2.8095e-08 0 2.8098e-08 0.0021 2.8101e-08 0 2.8275e-08 0 2.8278e-08 0.0021 2.8281e-08 0 2.8455e-08 0 2.8458e-08 0.0021 2.8461e-08 0 2.8635e-08 0 2.8638e-08 0.0021 2.8641e-08 0 2.8815e-08 0 2.8818e-08 0.0021 2.8821e-08 0 2.8995e-08 0 2.8998e-08 0.0021 2.9001e-08 0 2.9175e-08 0 2.9178e-08 0.0021 2.9181e-08 0 2.9355e-08 0 2.9358e-08 0.0021 2.9361e-08 0 2.9535e-08 0 2.9538e-08 0.0021 2.9541e-08 0 2.9715e-08 0 2.9718e-08 0.0021 2.9721e-08 0 2.9895e-08 0 2.9898e-08 0.0021 2.9901e-08 0 3.0075e-08 0 3.0078e-08 0.0021 3.0081e-08 0 3.0255e-08 0 3.0258e-08 0.0021 3.0261e-08 0 3.0435e-08 0 3.0438e-08 0.0021 3.0441e-08 0 3.0615e-08 0 3.0618e-08 0.0021 3.0621e-08 0 3.0795e-08 0 3.0798e-08 0.0021 3.0801e-08 0 3.0975e-08 0 3.0978e-08 0.0021 3.0981e-08 0 3.1155e-08 0 3.1158e-08 0.0021 3.1161e-08 0 3.1335e-08 0 3.1338e-08 0.0021 3.1341e-08 0 3.1515e-08 0 3.1518e-08 0.0021 3.1521e-08 0 3.1695e-08 0 3.1698e-08 0.0021 3.1701e-08 0 3.1875e-08 0 3.1878e-08 0.0021 3.1881e-08 0 3.2055e-08 0 3.2058e-08 0.0021 3.2061e-08 0 3.2235e-08 0 3.2238e-08 0.0021 3.2241e-08 0 3.2415e-08 0 3.2418e-08 0.0021 3.2421e-08 0 3.2595e-08 0 3.2598e-08 0.0021 3.2601e-08 0 3.2775e-08 0 3.2778e-08 0.0021 3.2781e-08 0 3.2955e-08 0 3.2958e-08 0.0021 3.2961e-08 0 3.3135e-08 0 3.3138e-08 0.0021 3.3141e-08 0 3.3315e-08 0 3.3318e-08 0.0021 3.3321e-08 0 3.3495e-08 0 3.3498e-08 0.0021 3.3501e-08 0 3.3675e-08 0 3.3678e-08 0.0021 3.3681e-08 0 3.3855e-08 0 3.3858e-08 0.0021 3.3861e-08 0 3.4035e-08 0 3.4038e-08 0.0021 3.4041e-08 0 3.4215e-08 0 3.4218e-08 0.0021 3.4221e-08 0 3.4395e-08 0 3.4398e-08 0.0021 3.4401e-08 0 3.4575e-08 0 3.4578e-08 0.0021 3.4581e-08 0 3.4755e-08 0 3.4758e-08 0.0021 3.4761e-08 0 3.4935e-08 0 3.4938e-08 0.0021 3.4941e-08 0 3.5115e-08 0 3.5118e-08 0.0021 3.5121e-08 0 3.5295e-08 0 3.5298e-08 0.0021 3.5301e-08 0 3.5475e-08 0 3.5478e-08 0.0021 3.5481e-08 0 3.5655e-08 0 3.5658e-08 0.0021 3.5661e-08 0 3.5835e-08 0 3.5838e-08 0.0021 3.5841e-08 0 3.6015e-08 0 3.6018e-08 0.0021 3.6021e-08 0 3.6195e-08 0 3.6198e-08 0.0021 3.6201e-08 0 3.6375e-08 0 3.6378e-08 0.0021 3.6381e-08 0 3.6555e-08 0 3.6558e-08 0.0021 3.6561e-08 0 3.6735e-08 0 3.6738e-08 0.0021 3.6741e-08 0 3.6915e-08 0 3.6918e-08 0.0021 3.6921e-08 0 3.7095e-08 0 3.7098e-08 0.0021 3.7101e-08 0 3.7275e-08 0 3.7278e-08 0.0021 3.7281e-08 0 3.7455e-08 0 3.7458e-08 0.0021 3.7461e-08 0 3.7635e-08 0 3.7638e-08 0.0021 3.7641e-08 0 3.7815e-08 0 3.7818e-08 0.0021 3.7821e-08 0 3.7995e-08 0 3.7998e-08 0.0021 3.8001e-08 0 3.8175e-08 0 3.8178e-08 0.0021 3.8181e-08 0 3.8355e-08 0 3.8358e-08 0.0021 3.8361e-08 0 3.8535e-08 0 3.8538e-08 0.0021 3.8541e-08 0 3.8715e-08 0 3.8718e-08 0.0021 3.8721e-08 0 3.8895e-08 0 3.8898e-08 0.0021 3.8901e-08 0 3.9075e-08 0 3.9078e-08 0.0021 3.9081e-08 0 3.9255e-08 0 3.9258e-08 0.0021 3.9261e-08 0 3.9435e-08 0 3.9438e-08 0.0021 3.9441e-08 0 3.9615e-08 0 3.9618e-08 0.0021 3.9621e-08 0 3.9795e-08 0 3.9798e-08 0.0021 3.9801e-08 0 3.9975e-08 0 3.9978e-08 0.0021 3.9981e-08 0 4.0155e-08 0 4.0158e-08 0.0021 4.0161e-08 0 4.0335e-08 0 4.0338e-08 0.0021 4.0341e-08 0 4.0515e-08 0 4.0518e-08 0.0021 4.0521e-08 0 4.0695e-08 0 4.0698e-08 0.0021 4.0701e-08 0 4.0875e-08 0 4.0878e-08 0.0021 4.0881e-08 0 4.1055e-08 0 4.1058e-08 0.0021 4.1061e-08 0 4.1235e-08 0 4.1238e-08 0.0021 4.1241e-08 0 4.1415e-08 0 4.1418e-08 0.0021 4.1421e-08 0 4.1595e-08 0 4.1598e-08 0.0021 4.1601e-08 0 4.1775e-08 0 4.1778e-08 0.0021 4.1781e-08 0 4.1955e-08 0 4.1958e-08 0.0021 4.1961e-08 0 4.2135e-08 0 4.2138e-08 0.0021 4.2141e-08 0 4.2315e-08 0 4.2318e-08 0.0021 4.2321e-08 0 4.2495e-08 0 4.2498e-08 0.0021 4.2501e-08 0 4.2675e-08 0 4.2678e-08 0.0021 4.2681e-08 0 4.2855e-08 0 4.2858e-08 0.0021 4.2861e-08 0 4.3035e-08 0 4.3038e-08 0.0021 4.3041e-08 0 4.3215e-08 0 4.3218e-08 0.0021 4.3221e-08 0 4.3395e-08 0 4.3398e-08 0.0021 4.3401e-08 0 4.3575e-08 0 4.3578e-08 0.0021 4.3581e-08 0 4.3755e-08 0 4.3758e-08 0.0021 4.3761e-08 0 4.3935e-08 0 4.3938e-08 0.0021 4.3941e-08 0 4.4115e-08 0 4.4118e-08 0.0021 4.4121e-08 0 4.4295e-08 0 4.4298e-08 0.0021 4.4301e-08 0 4.4475e-08 0 4.4478e-08 0.0021 4.4481e-08 0 4.4655e-08 0 4.4658e-08 0.0021 4.4661e-08 0 4.4835e-08 0 4.4838e-08 0.0021 4.4841e-08 0 4.5015e-08 0 4.5018e-08 0.0021 4.5021e-08 0 4.5195e-08 0 4.5198e-08 0.0021 4.5201e-08 0 4.5375e-08 0 4.5378e-08 0.0021 4.5381e-08 0 4.5555e-08 0 4.5558e-08 0.0021 4.5561e-08 0 4.5735e-08 0 4.5738e-08 0.0021 4.5741e-08 0 4.5915e-08 0 4.5918e-08 0.0021 4.5921e-08 0)
IT02|T 0 T02  PWL(0 0 1.5e-11 0 1.8e-11 0.0021 2.1e-11 0 1.95e-10 0 1.98e-10 0.0021 2.01e-10 0 3.75e-10 0 3.78e-10 0.0021 3.81e-10 0 5.55e-10 0 5.58e-10 0.0021 5.61e-10 0 7.35e-10 0 7.38e-10 0.0021 7.41e-10 0 9.15e-10 0 9.18e-10 0.0021 9.21e-10 0 1.095e-09 0 1.098e-09 0.0021 1.101e-09 0 1.275e-09 0 1.278e-09 0.0021 1.281e-09 0 1.455e-09 0 1.458e-09 0.0021 1.461e-09 0 1.635e-09 0 1.638e-09 0.0021 1.641e-09 0 1.815e-09 0 1.818e-09 0.0021 1.821e-09 0 1.995e-09 0 1.998e-09 0.0021 2.001e-09 0 2.175e-09 0 2.178e-09 0.0021 2.181e-09 0 2.355e-09 0 2.358e-09 0.0021 2.361e-09 0 2.535e-09 0 2.538e-09 0.0021 2.541e-09 0 2.715e-09 0 2.718e-09 0.0021 2.721e-09 0 2.895e-09 0 2.898e-09 0.0021 2.901e-09 0 3.075e-09 0 3.078e-09 0.0021 3.081e-09 0 3.255e-09 0 3.258e-09 0.0021 3.261e-09 0 3.435e-09 0 3.438e-09 0.0021 3.441e-09 0 3.615e-09 0 3.618e-09 0.0021 3.621e-09 0 3.795e-09 0 3.798e-09 0.0021 3.801e-09 0 3.975e-09 0 3.978e-09 0.0021 3.981e-09 0 4.155e-09 0 4.158e-09 0.0021 4.161e-09 0 4.335e-09 0 4.338e-09 0.0021 4.341e-09 0 4.515e-09 0 4.518e-09 0.0021 4.521e-09 0 4.695e-09 0 4.698e-09 0.0021 4.701e-09 0 4.875e-09 0 4.878e-09 0.0021 4.881e-09 0 5.055e-09 0 5.058e-09 0.0021 5.061e-09 0 5.235e-09 0 5.238e-09 0.0021 5.241e-09 0 5.415e-09 0 5.418e-09 0.0021 5.421e-09 0 5.595e-09 0 5.598e-09 0.0021 5.601e-09 0 5.775e-09 0 5.778e-09 0.0021 5.781e-09 0 5.955e-09 0 5.958e-09 0.0021 5.961e-09 0 6.135e-09 0 6.138e-09 0.0021 6.141e-09 0 6.315e-09 0 6.318e-09 0.0021 6.321e-09 0 6.495e-09 0 6.498e-09 0.0021 6.501e-09 0 6.675e-09 0 6.678e-09 0.0021 6.681e-09 0 6.855e-09 0 6.858e-09 0.0021 6.861e-09 0 7.035e-09 0 7.038e-09 0.0021 7.041e-09 0 7.215e-09 0 7.218e-09 0.0021 7.221e-09 0 7.395e-09 0 7.398e-09 0.0021 7.401e-09 0 7.575e-09 0 7.578e-09 0.0021 7.581e-09 0 7.755e-09 0 7.758e-09 0.0021 7.761e-09 0 7.935e-09 0 7.938e-09 0.0021 7.941e-09 0 8.115e-09 0 8.118e-09 0.0021 8.121e-09 0 8.295e-09 0 8.298e-09 0.0021 8.301e-09 0 8.475e-09 0 8.478e-09 0.0021 8.481e-09 0 8.655e-09 0 8.658e-09 0.0021 8.661e-09 0 8.835e-09 0 8.838e-09 0.0021 8.841e-09 0 9.015e-09 0 9.018e-09 0.0021 9.021e-09 0 9.195e-09 0 9.198e-09 0.0021 9.201e-09 0 9.375e-09 0 9.378e-09 0.0021 9.381e-09 0 9.555e-09 0 9.558e-09 0.0021 9.561e-09 0 9.735e-09 0 9.738e-09 0.0021 9.741e-09 0 9.915e-09 0 9.918e-09 0.0021 9.921e-09 0 1.0095e-08 0 1.0098e-08 0.0021 1.0101e-08 0 1.0275e-08 0 1.0278e-08 0.0021 1.0281e-08 0 1.0455e-08 0 1.0458e-08 0.0021 1.0461e-08 0 1.0635e-08 0 1.0638e-08 0.0021 1.0641e-08 0 1.0815e-08 0 1.0818e-08 0.0021 1.0821e-08 0 1.0995e-08 0 1.0998e-08 0.0021 1.1001e-08 0 1.1175e-08 0 1.1178e-08 0.0021 1.1181e-08 0 1.1355e-08 0 1.1358e-08 0.0021 1.1361e-08 0 1.1535e-08 0 1.1538e-08 0.0021 1.1541e-08 0 1.1715e-08 0 1.1718e-08 0.0021 1.1721e-08 0 1.1895e-08 0 1.1898e-08 0.0021 1.1901e-08 0 1.2075e-08 0 1.2078e-08 0.0021 1.2081e-08 0 1.2255e-08 0 1.2258e-08 0.0021 1.2261e-08 0 1.2435e-08 0 1.2438e-08 0.0021 1.2441e-08 0 1.2615e-08 0 1.2618e-08 0.0021 1.2621e-08 0 1.2795e-08 0 1.2798e-08 0.0021 1.2801e-08 0 1.2975e-08 0 1.2978e-08 0.0021 1.2981e-08 0 1.3155e-08 0 1.3158e-08 0.0021 1.3161e-08 0 1.3335e-08 0 1.3338e-08 0.0021 1.3341e-08 0 1.3515e-08 0 1.3518e-08 0.0021 1.3521e-08 0 1.3695e-08 0 1.3698e-08 0.0021 1.3701e-08 0 1.3875e-08 0 1.3878e-08 0.0021 1.3881e-08 0 1.4055e-08 0 1.4058e-08 0.0021 1.4061e-08 0 1.4235e-08 0 1.4238e-08 0.0021 1.4241e-08 0 1.4415e-08 0 1.4418e-08 0.0021 1.4421e-08 0 1.4595e-08 0 1.4598e-08 0.0021 1.4601e-08 0 1.4775e-08 0 1.4778e-08 0.0021 1.4781e-08 0 1.4955e-08 0 1.4958e-08 0.0021 1.4961e-08 0 1.5135e-08 0 1.5138e-08 0.0021 1.5141e-08 0 1.5315e-08 0 1.5318e-08 0.0021 1.5321e-08 0 1.5495e-08 0 1.5498e-08 0.0021 1.5501e-08 0 1.5675e-08 0 1.5678e-08 0.0021 1.5681e-08 0 1.5855e-08 0 1.5858e-08 0.0021 1.5861e-08 0 1.6035e-08 0 1.6038e-08 0.0021 1.6041e-08 0 1.6215e-08 0 1.6218e-08 0.0021 1.6221e-08 0 1.6395e-08 0 1.6398e-08 0.0021 1.6401e-08 0 1.6575e-08 0 1.6578e-08 0.0021 1.6581e-08 0 1.6755e-08 0 1.6758e-08 0.0021 1.6761e-08 0 1.6935e-08 0 1.6938e-08 0.0021 1.6941e-08 0 1.7115e-08 0 1.7118e-08 0.0021 1.7121e-08 0 1.7295e-08 0 1.7298e-08 0.0021 1.7301e-08 0 1.7475e-08 0 1.7478e-08 0.0021 1.7481e-08 0 1.7655e-08 0 1.7658e-08 0.0021 1.7661e-08 0 1.7835e-08 0 1.7838e-08 0.0021 1.7841e-08 0 1.8015e-08 0 1.8018e-08 0.0021 1.8021e-08 0 1.8195e-08 0 1.8198e-08 0.0021 1.8201e-08 0 1.8375e-08 0 1.8378e-08 0.0021 1.8381e-08 0 1.8555e-08 0 1.8558e-08 0.0021 1.8561e-08 0 1.8735e-08 0 1.8738e-08 0.0021 1.8741e-08 0 1.8915e-08 0 1.8918e-08 0.0021 1.8921e-08 0 1.9095e-08 0 1.9098e-08 0.0021 1.9101e-08 0 1.9275e-08 0 1.9278e-08 0.0021 1.9281e-08 0 1.9455e-08 0 1.9458e-08 0.0021 1.9461e-08 0 1.9635e-08 0 1.9638e-08 0.0021 1.9641e-08 0 1.9815e-08 0 1.9818e-08 0.0021 1.9821e-08 0 1.9995e-08 0 1.9998e-08 0.0021 2.0001e-08 0 2.0175e-08 0 2.0178e-08 0.0021 2.0181e-08 0 2.0355e-08 0 2.0358e-08 0.0021 2.0361e-08 0 2.0535e-08 0 2.0538e-08 0.0021 2.0541e-08 0 2.0715e-08 0 2.0718e-08 0.0021 2.0721e-08 0 2.0895e-08 0 2.0898e-08 0.0021 2.0901e-08 0 2.1075e-08 0 2.1078e-08 0.0021 2.1081e-08 0 2.1255e-08 0 2.1258e-08 0.0021 2.1261e-08 0 2.1435e-08 0 2.1438e-08 0.0021 2.1441e-08 0 2.1615e-08 0 2.1618e-08 0.0021 2.1621e-08 0 2.1795e-08 0 2.1798e-08 0.0021 2.1801e-08 0 2.1975e-08 0 2.1978e-08 0.0021 2.1981e-08 0 2.2155e-08 0 2.2158e-08 0.0021 2.2161e-08 0 2.2335e-08 0 2.2338e-08 0.0021 2.2341e-08 0 2.2515e-08 0 2.2518e-08 0.0021 2.2521e-08 0 2.2695e-08 0 2.2698e-08 0.0021 2.2701e-08 0 2.2875e-08 0 2.2878e-08 0.0021 2.2881e-08 0 2.3055e-08 0 2.3058e-08 0.0021 2.3061e-08 0 2.3235e-08 0 2.3238e-08 0.0021 2.3241e-08 0 2.3415e-08 0 2.3418e-08 0.0021 2.3421e-08 0 2.3595e-08 0 2.3598e-08 0.0021 2.3601e-08 0 2.3775e-08 0 2.3778e-08 0.0021 2.3781e-08 0 2.3955e-08 0 2.3958e-08 0.0021 2.3961e-08 0 2.4135e-08 0 2.4138e-08 0.0021 2.4141e-08 0 2.4315e-08 0 2.4318e-08 0.0021 2.4321e-08 0 2.4495e-08 0 2.4498e-08 0.0021 2.4501e-08 0 2.4675e-08 0 2.4678e-08 0.0021 2.4681e-08 0 2.4855e-08 0 2.4858e-08 0.0021 2.4861e-08 0 2.5035e-08 0 2.5038e-08 0.0021 2.5041e-08 0 2.5215e-08 0 2.5218e-08 0.0021 2.5221e-08 0 2.5395e-08 0 2.5398e-08 0.0021 2.5401e-08 0 2.5575e-08 0 2.5578e-08 0.0021 2.5581e-08 0 2.5755e-08 0 2.5758e-08 0.0021 2.5761e-08 0 2.5935e-08 0 2.5938e-08 0.0021 2.5941e-08 0 2.6115e-08 0 2.6118e-08 0.0021 2.6121e-08 0 2.6295e-08 0 2.6298e-08 0.0021 2.6301e-08 0 2.6475e-08 0 2.6478e-08 0.0021 2.6481e-08 0 2.6655e-08 0 2.6658e-08 0.0021 2.6661e-08 0 2.6835e-08 0 2.6838e-08 0.0021 2.6841e-08 0 2.7015e-08 0 2.7018e-08 0.0021 2.7021e-08 0 2.7195e-08 0 2.7198e-08 0.0021 2.7201e-08 0 2.7375e-08 0 2.7378e-08 0.0021 2.7381e-08 0 2.7555e-08 0 2.7558e-08 0.0021 2.7561e-08 0 2.7735e-08 0 2.7738e-08 0.0021 2.7741e-08 0 2.7915e-08 0 2.7918e-08 0.0021 2.7921e-08 0 2.8095e-08 0 2.8098e-08 0.0021 2.8101e-08 0 2.8275e-08 0 2.8278e-08 0.0021 2.8281e-08 0 2.8455e-08 0 2.8458e-08 0.0021 2.8461e-08 0 2.8635e-08 0 2.8638e-08 0.0021 2.8641e-08 0 2.8815e-08 0 2.8818e-08 0.0021 2.8821e-08 0 2.8995e-08 0 2.8998e-08 0.0021 2.9001e-08 0 2.9175e-08 0 2.9178e-08 0.0021 2.9181e-08 0 2.9355e-08 0 2.9358e-08 0.0021 2.9361e-08 0 2.9535e-08 0 2.9538e-08 0.0021 2.9541e-08 0 2.9715e-08 0 2.9718e-08 0.0021 2.9721e-08 0 2.9895e-08 0 2.9898e-08 0.0021 2.9901e-08 0 3.0075e-08 0 3.0078e-08 0.0021 3.0081e-08 0 3.0255e-08 0 3.0258e-08 0.0021 3.0261e-08 0 3.0435e-08 0 3.0438e-08 0.0021 3.0441e-08 0 3.0615e-08 0 3.0618e-08 0.0021 3.0621e-08 0 3.0795e-08 0 3.0798e-08 0.0021 3.0801e-08 0 3.0975e-08 0 3.0978e-08 0.0021 3.0981e-08 0 3.1155e-08 0 3.1158e-08 0.0021 3.1161e-08 0 3.1335e-08 0 3.1338e-08 0.0021 3.1341e-08 0 3.1515e-08 0 3.1518e-08 0.0021 3.1521e-08 0 3.1695e-08 0 3.1698e-08 0.0021 3.1701e-08 0 3.1875e-08 0 3.1878e-08 0.0021 3.1881e-08 0 3.2055e-08 0 3.2058e-08 0.0021 3.2061e-08 0 3.2235e-08 0 3.2238e-08 0.0021 3.2241e-08 0 3.2415e-08 0 3.2418e-08 0.0021 3.2421e-08 0 3.2595e-08 0 3.2598e-08 0.0021 3.2601e-08 0 3.2775e-08 0 3.2778e-08 0.0021 3.2781e-08 0 3.2955e-08 0 3.2958e-08 0.0021 3.2961e-08 0 3.3135e-08 0 3.3138e-08 0.0021 3.3141e-08 0 3.3315e-08 0 3.3318e-08 0.0021 3.3321e-08 0 3.3495e-08 0 3.3498e-08 0.0021 3.3501e-08 0 3.3675e-08 0 3.3678e-08 0.0021 3.3681e-08 0 3.3855e-08 0 3.3858e-08 0.0021 3.3861e-08 0 3.4035e-08 0 3.4038e-08 0.0021 3.4041e-08 0 3.4215e-08 0 3.4218e-08 0.0021 3.4221e-08 0 3.4395e-08 0 3.4398e-08 0.0021 3.4401e-08 0 3.4575e-08 0 3.4578e-08 0.0021 3.4581e-08 0 3.4755e-08 0 3.4758e-08 0.0021 3.4761e-08 0 3.4935e-08 0 3.4938e-08 0.0021 3.4941e-08 0 3.5115e-08 0 3.5118e-08 0.0021 3.5121e-08 0 3.5295e-08 0 3.5298e-08 0.0021 3.5301e-08 0 3.5475e-08 0 3.5478e-08 0.0021 3.5481e-08 0 3.5655e-08 0 3.5658e-08 0.0021 3.5661e-08 0 3.5835e-08 0 3.5838e-08 0.0021 3.5841e-08 0 3.6015e-08 0 3.6018e-08 0.0021 3.6021e-08 0 3.6195e-08 0 3.6198e-08 0.0021 3.6201e-08 0 3.6375e-08 0 3.6378e-08 0.0021 3.6381e-08 0 3.6555e-08 0 3.6558e-08 0.0021 3.6561e-08 0 3.6735e-08 0 3.6738e-08 0.0021 3.6741e-08 0 3.6915e-08 0 3.6918e-08 0.0021 3.6921e-08 0 3.7095e-08 0 3.7098e-08 0.0021 3.7101e-08 0 3.7275e-08 0 3.7278e-08 0.0021 3.7281e-08 0 3.7455e-08 0 3.7458e-08 0.0021 3.7461e-08 0 3.7635e-08 0 3.7638e-08 0.0021 3.7641e-08 0 3.7815e-08 0 3.7818e-08 0.0021 3.7821e-08 0 3.7995e-08 0 3.7998e-08 0.0021 3.8001e-08 0 3.8175e-08 0 3.8178e-08 0.0021 3.8181e-08 0 3.8355e-08 0 3.8358e-08 0.0021 3.8361e-08 0 3.8535e-08 0 3.8538e-08 0.0021 3.8541e-08 0 3.8715e-08 0 3.8718e-08 0.0021 3.8721e-08 0 3.8895e-08 0 3.8898e-08 0.0021 3.8901e-08 0 3.9075e-08 0 3.9078e-08 0.0021 3.9081e-08 0 3.9255e-08 0 3.9258e-08 0.0021 3.9261e-08 0 3.9435e-08 0 3.9438e-08 0.0021 3.9441e-08 0 3.9615e-08 0 3.9618e-08 0.0021 3.9621e-08 0 3.9795e-08 0 3.9798e-08 0.0021 3.9801e-08 0 3.9975e-08 0 3.9978e-08 0.0021 3.9981e-08 0 4.0155e-08 0 4.0158e-08 0.0021 4.0161e-08 0 4.0335e-08 0 4.0338e-08 0.0021 4.0341e-08 0 4.0515e-08 0 4.0518e-08 0.0021 4.0521e-08 0 4.0695e-08 0 4.0698e-08 0.0021 4.0701e-08 0 4.0875e-08 0 4.0878e-08 0.0021 4.0881e-08 0 4.1055e-08 0 4.1058e-08 0.0021 4.1061e-08 0 4.1235e-08 0 4.1238e-08 0.0021 4.1241e-08 0 4.1415e-08 0 4.1418e-08 0.0021 4.1421e-08 0 4.1595e-08 0 4.1598e-08 0.0021 4.1601e-08 0 4.1775e-08 0 4.1778e-08 0.0021 4.1781e-08 0 4.1955e-08 0 4.1958e-08 0.0021 4.1961e-08 0 4.2135e-08 0 4.2138e-08 0.0021 4.2141e-08 0 4.2315e-08 0 4.2318e-08 0.0021 4.2321e-08 0 4.2495e-08 0 4.2498e-08 0.0021 4.2501e-08 0 4.2675e-08 0 4.2678e-08 0.0021 4.2681e-08 0 4.2855e-08 0 4.2858e-08 0.0021 4.2861e-08 0 4.3035e-08 0 4.3038e-08 0.0021 4.3041e-08 0 4.3215e-08 0 4.3218e-08 0.0021 4.3221e-08 0 4.3395e-08 0 4.3398e-08 0.0021 4.3401e-08 0 4.3575e-08 0 4.3578e-08 0.0021 4.3581e-08 0 4.3755e-08 0 4.3758e-08 0.0021 4.3761e-08 0 4.3935e-08 0 4.3938e-08 0.0021 4.3941e-08 0 4.4115e-08 0 4.4118e-08 0.0021 4.4121e-08 0 4.4295e-08 0 4.4298e-08 0.0021 4.4301e-08 0 4.4475e-08 0 4.4478e-08 0.0021 4.4481e-08 0 4.4655e-08 0 4.4658e-08 0.0021 4.4661e-08 0 4.4835e-08 0 4.4838e-08 0.0021 4.4841e-08 0 4.5015e-08 0 4.5018e-08 0.0021 4.5021e-08 0 4.5195e-08 0 4.5198e-08 0.0021 4.5201e-08 0 4.5375e-08 0 4.5378e-08 0.0021 4.5381e-08 0 4.5555e-08 0 4.5558e-08 0.0021 4.5561e-08 0 4.5735e-08 0 4.5738e-08 0.0021 4.5741e-08 0 4.5915e-08 0 4.5918e-08 0.0021 4.5921e-08 0)
IT03|T 0 T03  PWL(0 0 1.5e-11 0 1.8e-11 0.0021 2.1e-11 0 1.95e-10 0 1.98e-10 0.0021 2.01e-10 0 3.75e-10 0 3.78e-10 0.0021 3.81e-10 0 5.55e-10 0 5.58e-10 0.0021 5.61e-10 0 7.35e-10 0 7.38e-10 0.0021 7.41e-10 0 9.15e-10 0 9.18e-10 0.0021 9.21e-10 0 1.095e-09 0 1.098e-09 0.0021 1.101e-09 0 1.275e-09 0 1.278e-09 0.0021 1.281e-09 0 1.455e-09 0 1.458e-09 0.0021 1.461e-09 0 1.635e-09 0 1.638e-09 0.0021 1.641e-09 0 1.815e-09 0 1.818e-09 0.0021 1.821e-09 0 1.995e-09 0 1.998e-09 0.0021 2.001e-09 0 2.175e-09 0 2.178e-09 0.0021 2.181e-09 0 2.355e-09 0 2.358e-09 0.0021 2.361e-09 0 2.535e-09 0 2.538e-09 0.0021 2.541e-09 0 2.715e-09 0 2.718e-09 0.0021 2.721e-09 0 2.895e-09 0 2.898e-09 0.0021 2.901e-09 0 3.075e-09 0 3.078e-09 0.0021 3.081e-09 0 3.255e-09 0 3.258e-09 0.0021 3.261e-09 0 3.435e-09 0 3.438e-09 0.0021 3.441e-09 0 3.615e-09 0 3.618e-09 0.0021 3.621e-09 0 3.795e-09 0 3.798e-09 0.0021 3.801e-09 0 3.975e-09 0 3.978e-09 0.0021 3.981e-09 0 4.155e-09 0 4.158e-09 0.0021 4.161e-09 0 4.335e-09 0 4.338e-09 0.0021 4.341e-09 0 4.515e-09 0 4.518e-09 0.0021 4.521e-09 0 4.695e-09 0 4.698e-09 0.0021 4.701e-09 0 4.875e-09 0 4.878e-09 0.0021 4.881e-09 0 5.055e-09 0 5.058e-09 0.0021 5.061e-09 0 5.235e-09 0 5.238e-09 0.0021 5.241e-09 0 5.415e-09 0 5.418e-09 0.0021 5.421e-09 0 5.595e-09 0 5.598e-09 0.0021 5.601e-09 0 5.775e-09 0 5.778e-09 0.0021 5.781e-09 0 5.955e-09 0 5.958e-09 0.0021 5.961e-09 0 6.135e-09 0 6.138e-09 0.0021 6.141e-09 0 6.315e-09 0 6.318e-09 0.0021 6.321e-09 0 6.495e-09 0 6.498e-09 0.0021 6.501e-09 0 6.675e-09 0 6.678e-09 0.0021 6.681e-09 0 6.855e-09 0 6.858e-09 0.0021 6.861e-09 0 7.035e-09 0 7.038e-09 0.0021 7.041e-09 0 7.215e-09 0 7.218e-09 0.0021 7.221e-09 0 7.395e-09 0 7.398e-09 0.0021 7.401e-09 0 7.575e-09 0 7.578e-09 0.0021 7.581e-09 0 7.755e-09 0 7.758e-09 0.0021 7.761e-09 0 7.935e-09 0 7.938e-09 0.0021 7.941e-09 0 8.115e-09 0 8.118e-09 0.0021 8.121e-09 0 8.295e-09 0 8.298e-09 0.0021 8.301e-09 0 8.475e-09 0 8.478e-09 0.0021 8.481e-09 0 8.655e-09 0 8.658e-09 0.0021 8.661e-09 0 8.835e-09 0 8.838e-09 0.0021 8.841e-09 0 9.015e-09 0 9.018e-09 0.0021 9.021e-09 0 9.195e-09 0 9.198e-09 0.0021 9.201e-09 0 9.375e-09 0 9.378e-09 0.0021 9.381e-09 0 9.555e-09 0 9.558e-09 0.0021 9.561e-09 0 9.735e-09 0 9.738e-09 0.0021 9.741e-09 0 9.915e-09 0 9.918e-09 0.0021 9.921e-09 0 1.0095e-08 0 1.0098e-08 0.0021 1.0101e-08 0 1.0275e-08 0 1.0278e-08 0.0021 1.0281e-08 0 1.0455e-08 0 1.0458e-08 0.0021 1.0461e-08 0 1.0635e-08 0 1.0638e-08 0.0021 1.0641e-08 0 1.0815e-08 0 1.0818e-08 0.0021 1.0821e-08 0 1.0995e-08 0 1.0998e-08 0.0021 1.1001e-08 0 1.1175e-08 0 1.1178e-08 0.0021 1.1181e-08 0 1.1355e-08 0 1.1358e-08 0.0021 1.1361e-08 0 1.1535e-08 0 1.1538e-08 0.0021 1.1541e-08 0 1.1715e-08 0 1.1718e-08 0.0021 1.1721e-08 0 1.1895e-08 0 1.1898e-08 0.0021 1.1901e-08 0 1.2075e-08 0 1.2078e-08 0.0021 1.2081e-08 0 1.2255e-08 0 1.2258e-08 0.0021 1.2261e-08 0 1.2435e-08 0 1.2438e-08 0.0021 1.2441e-08 0 1.2615e-08 0 1.2618e-08 0.0021 1.2621e-08 0 1.2795e-08 0 1.2798e-08 0.0021 1.2801e-08 0 1.2975e-08 0 1.2978e-08 0.0021 1.2981e-08 0 1.3155e-08 0 1.3158e-08 0.0021 1.3161e-08 0 1.3335e-08 0 1.3338e-08 0.0021 1.3341e-08 0 1.3515e-08 0 1.3518e-08 0.0021 1.3521e-08 0 1.3695e-08 0 1.3698e-08 0.0021 1.3701e-08 0 1.3875e-08 0 1.3878e-08 0.0021 1.3881e-08 0 1.4055e-08 0 1.4058e-08 0.0021 1.4061e-08 0 1.4235e-08 0 1.4238e-08 0.0021 1.4241e-08 0 1.4415e-08 0 1.4418e-08 0.0021 1.4421e-08 0 1.4595e-08 0 1.4598e-08 0.0021 1.4601e-08 0 1.4775e-08 0 1.4778e-08 0.0021 1.4781e-08 0 1.4955e-08 0 1.4958e-08 0.0021 1.4961e-08 0 1.5135e-08 0 1.5138e-08 0.0021 1.5141e-08 0 1.5315e-08 0 1.5318e-08 0.0021 1.5321e-08 0 1.5495e-08 0 1.5498e-08 0.0021 1.5501e-08 0 1.5675e-08 0 1.5678e-08 0.0021 1.5681e-08 0 1.5855e-08 0 1.5858e-08 0.0021 1.5861e-08 0 1.6035e-08 0 1.6038e-08 0.0021 1.6041e-08 0 1.6215e-08 0 1.6218e-08 0.0021 1.6221e-08 0 1.6395e-08 0 1.6398e-08 0.0021 1.6401e-08 0 1.6575e-08 0 1.6578e-08 0.0021 1.6581e-08 0 1.6755e-08 0 1.6758e-08 0.0021 1.6761e-08 0 1.6935e-08 0 1.6938e-08 0.0021 1.6941e-08 0 1.7115e-08 0 1.7118e-08 0.0021 1.7121e-08 0 1.7295e-08 0 1.7298e-08 0.0021 1.7301e-08 0 1.7475e-08 0 1.7478e-08 0.0021 1.7481e-08 0 1.7655e-08 0 1.7658e-08 0.0021 1.7661e-08 0 1.7835e-08 0 1.7838e-08 0.0021 1.7841e-08 0 1.8015e-08 0 1.8018e-08 0.0021 1.8021e-08 0 1.8195e-08 0 1.8198e-08 0.0021 1.8201e-08 0 1.8375e-08 0 1.8378e-08 0.0021 1.8381e-08 0 1.8555e-08 0 1.8558e-08 0.0021 1.8561e-08 0 1.8735e-08 0 1.8738e-08 0.0021 1.8741e-08 0 1.8915e-08 0 1.8918e-08 0.0021 1.8921e-08 0 1.9095e-08 0 1.9098e-08 0.0021 1.9101e-08 0 1.9275e-08 0 1.9278e-08 0.0021 1.9281e-08 0 1.9455e-08 0 1.9458e-08 0.0021 1.9461e-08 0 1.9635e-08 0 1.9638e-08 0.0021 1.9641e-08 0 1.9815e-08 0 1.9818e-08 0.0021 1.9821e-08 0 1.9995e-08 0 1.9998e-08 0.0021 2.0001e-08 0 2.0175e-08 0 2.0178e-08 0.0021 2.0181e-08 0 2.0355e-08 0 2.0358e-08 0.0021 2.0361e-08 0 2.0535e-08 0 2.0538e-08 0.0021 2.0541e-08 0 2.0715e-08 0 2.0718e-08 0.0021 2.0721e-08 0 2.0895e-08 0 2.0898e-08 0.0021 2.0901e-08 0 2.1075e-08 0 2.1078e-08 0.0021 2.1081e-08 0 2.1255e-08 0 2.1258e-08 0.0021 2.1261e-08 0 2.1435e-08 0 2.1438e-08 0.0021 2.1441e-08 0 2.1615e-08 0 2.1618e-08 0.0021 2.1621e-08 0 2.1795e-08 0 2.1798e-08 0.0021 2.1801e-08 0 2.1975e-08 0 2.1978e-08 0.0021 2.1981e-08 0 2.2155e-08 0 2.2158e-08 0.0021 2.2161e-08 0 2.2335e-08 0 2.2338e-08 0.0021 2.2341e-08 0 2.2515e-08 0 2.2518e-08 0.0021 2.2521e-08 0 2.2695e-08 0 2.2698e-08 0.0021 2.2701e-08 0 2.2875e-08 0 2.2878e-08 0.0021 2.2881e-08 0 2.3055e-08 0 2.3058e-08 0.0021 2.3061e-08 0 2.3235e-08 0 2.3238e-08 0.0021 2.3241e-08 0 2.3415e-08 0 2.3418e-08 0.0021 2.3421e-08 0 2.3595e-08 0 2.3598e-08 0.0021 2.3601e-08 0 2.3775e-08 0 2.3778e-08 0.0021 2.3781e-08 0 2.3955e-08 0 2.3958e-08 0.0021 2.3961e-08 0 2.4135e-08 0 2.4138e-08 0.0021 2.4141e-08 0 2.4315e-08 0 2.4318e-08 0.0021 2.4321e-08 0 2.4495e-08 0 2.4498e-08 0.0021 2.4501e-08 0 2.4675e-08 0 2.4678e-08 0.0021 2.4681e-08 0 2.4855e-08 0 2.4858e-08 0.0021 2.4861e-08 0 2.5035e-08 0 2.5038e-08 0.0021 2.5041e-08 0 2.5215e-08 0 2.5218e-08 0.0021 2.5221e-08 0 2.5395e-08 0 2.5398e-08 0.0021 2.5401e-08 0 2.5575e-08 0 2.5578e-08 0.0021 2.5581e-08 0 2.5755e-08 0 2.5758e-08 0.0021 2.5761e-08 0 2.5935e-08 0 2.5938e-08 0.0021 2.5941e-08 0 2.6115e-08 0 2.6118e-08 0.0021 2.6121e-08 0 2.6295e-08 0 2.6298e-08 0.0021 2.6301e-08 0 2.6475e-08 0 2.6478e-08 0.0021 2.6481e-08 0 2.6655e-08 0 2.6658e-08 0.0021 2.6661e-08 0 2.6835e-08 0 2.6838e-08 0.0021 2.6841e-08 0 2.7015e-08 0 2.7018e-08 0.0021 2.7021e-08 0 2.7195e-08 0 2.7198e-08 0.0021 2.7201e-08 0 2.7375e-08 0 2.7378e-08 0.0021 2.7381e-08 0 2.7555e-08 0 2.7558e-08 0.0021 2.7561e-08 0 2.7735e-08 0 2.7738e-08 0.0021 2.7741e-08 0 2.7915e-08 0 2.7918e-08 0.0021 2.7921e-08 0 2.8095e-08 0 2.8098e-08 0.0021 2.8101e-08 0 2.8275e-08 0 2.8278e-08 0.0021 2.8281e-08 0 2.8455e-08 0 2.8458e-08 0.0021 2.8461e-08 0 2.8635e-08 0 2.8638e-08 0.0021 2.8641e-08 0 2.8815e-08 0 2.8818e-08 0.0021 2.8821e-08 0 2.8995e-08 0 2.8998e-08 0.0021 2.9001e-08 0 2.9175e-08 0 2.9178e-08 0.0021 2.9181e-08 0 2.9355e-08 0 2.9358e-08 0.0021 2.9361e-08 0 2.9535e-08 0 2.9538e-08 0.0021 2.9541e-08 0 2.9715e-08 0 2.9718e-08 0.0021 2.9721e-08 0 2.9895e-08 0 2.9898e-08 0.0021 2.9901e-08 0 3.0075e-08 0 3.0078e-08 0.0021 3.0081e-08 0 3.0255e-08 0 3.0258e-08 0.0021 3.0261e-08 0 3.0435e-08 0 3.0438e-08 0.0021 3.0441e-08 0 3.0615e-08 0 3.0618e-08 0.0021 3.0621e-08 0 3.0795e-08 0 3.0798e-08 0.0021 3.0801e-08 0 3.0975e-08 0 3.0978e-08 0.0021 3.0981e-08 0 3.1155e-08 0 3.1158e-08 0.0021 3.1161e-08 0 3.1335e-08 0 3.1338e-08 0.0021 3.1341e-08 0 3.1515e-08 0 3.1518e-08 0.0021 3.1521e-08 0 3.1695e-08 0 3.1698e-08 0.0021 3.1701e-08 0 3.1875e-08 0 3.1878e-08 0.0021 3.1881e-08 0 3.2055e-08 0 3.2058e-08 0.0021 3.2061e-08 0 3.2235e-08 0 3.2238e-08 0.0021 3.2241e-08 0 3.2415e-08 0 3.2418e-08 0.0021 3.2421e-08 0 3.2595e-08 0 3.2598e-08 0.0021 3.2601e-08 0 3.2775e-08 0 3.2778e-08 0.0021 3.2781e-08 0 3.2955e-08 0 3.2958e-08 0.0021 3.2961e-08 0 3.3135e-08 0 3.3138e-08 0.0021 3.3141e-08 0 3.3315e-08 0 3.3318e-08 0.0021 3.3321e-08 0 3.3495e-08 0 3.3498e-08 0.0021 3.3501e-08 0 3.3675e-08 0 3.3678e-08 0.0021 3.3681e-08 0 3.3855e-08 0 3.3858e-08 0.0021 3.3861e-08 0 3.4035e-08 0 3.4038e-08 0.0021 3.4041e-08 0 3.4215e-08 0 3.4218e-08 0.0021 3.4221e-08 0 3.4395e-08 0 3.4398e-08 0.0021 3.4401e-08 0 3.4575e-08 0 3.4578e-08 0.0021 3.4581e-08 0 3.4755e-08 0 3.4758e-08 0.0021 3.4761e-08 0 3.4935e-08 0 3.4938e-08 0.0021 3.4941e-08 0 3.5115e-08 0 3.5118e-08 0.0021 3.5121e-08 0 3.5295e-08 0 3.5298e-08 0.0021 3.5301e-08 0 3.5475e-08 0 3.5478e-08 0.0021 3.5481e-08 0 3.5655e-08 0 3.5658e-08 0.0021 3.5661e-08 0 3.5835e-08 0 3.5838e-08 0.0021 3.5841e-08 0 3.6015e-08 0 3.6018e-08 0.0021 3.6021e-08 0 3.6195e-08 0 3.6198e-08 0.0021 3.6201e-08 0 3.6375e-08 0 3.6378e-08 0.0021 3.6381e-08 0 3.6555e-08 0 3.6558e-08 0.0021 3.6561e-08 0 3.6735e-08 0 3.6738e-08 0.0021 3.6741e-08 0 3.6915e-08 0 3.6918e-08 0.0021 3.6921e-08 0 3.7095e-08 0 3.7098e-08 0.0021 3.7101e-08 0 3.7275e-08 0 3.7278e-08 0.0021 3.7281e-08 0 3.7455e-08 0 3.7458e-08 0.0021 3.7461e-08 0 3.7635e-08 0 3.7638e-08 0.0021 3.7641e-08 0 3.7815e-08 0 3.7818e-08 0.0021 3.7821e-08 0 3.7995e-08 0 3.7998e-08 0.0021 3.8001e-08 0 3.8175e-08 0 3.8178e-08 0.0021 3.8181e-08 0 3.8355e-08 0 3.8358e-08 0.0021 3.8361e-08 0 3.8535e-08 0 3.8538e-08 0.0021 3.8541e-08 0 3.8715e-08 0 3.8718e-08 0.0021 3.8721e-08 0 3.8895e-08 0 3.8898e-08 0.0021 3.8901e-08 0 3.9075e-08 0 3.9078e-08 0.0021 3.9081e-08 0 3.9255e-08 0 3.9258e-08 0.0021 3.9261e-08 0 3.9435e-08 0 3.9438e-08 0.0021 3.9441e-08 0 3.9615e-08 0 3.9618e-08 0.0021 3.9621e-08 0 3.9795e-08 0 3.9798e-08 0.0021 3.9801e-08 0 3.9975e-08 0 3.9978e-08 0.0021 3.9981e-08 0 4.0155e-08 0 4.0158e-08 0.0021 4.0161e-08 0 4.0335e-08 0 4.0338e-08 0.0021 4.0341e-08 0 4.0515e-08 0 4.0518e-08 0.0021 4.0521e-08 0 4.0695e-08 0 4.0698e-08 0.0021 4.0701e-08 0 4.0875e-08 0 4.0878e-08 0.0021 4.0881e-08 0 4.1055e-08 0 4.1058e-08 0.0021 4.1061e-08 0 4.1235e-08 0 4.1238e-08 0.0021 4.1241e-08 0 4.1415e-08 0 4.1418e-08 0.0021 4.1421e-08 0 4.1595e-08 0 4.1598e-08 0.0021 4.1601e-08 0 4.1775e-08 0 4.1778e-08 0.0021 4.1781e-08 0 4.1955e-08 0 4.1958e-08 0.0021 4.1961e-08 0 4.2135e-08 0 4.2138e-08 0.0021 4.2141e-08 0 4.2315e-08 0 4.2318e-08 0.0021 4.2321e-08 0 4.2495e-08 0 4.2498e-08 0.0021 4.2501e-08 0 4.2675e-08 0 4.2678e-08 0.0021 4.2681e-08 0 4.2855e-08 0 4.2858e-08 0.0021 4.2861e-08 0 4.3035e-08 0 4.3038e-08 0.0021 4.3041e-08 0 4.3215e-08 0 4.3218e-08 0.0021 4.3221e-08 0 4.3395e-08 0 4.3398e-08 0.0021 4.3401e-08 0 4.3575e-08 0 4.3578e-08 0.0021 4.3581e-08 0 4.3755e-08 0 4.3758e-08 0.0021 4.3761e-08 0 4.3935e-08 0 4.3938e-08 0.0021 4.3941e-08 0 4.4115e-08 0 4.4118e-08 0.0021 4.4121e-08 0 4.4295e-08 0 4.4298e-08 0.0021 4.4301e-08 0 4.4475e-08 0 4.4478e-08 0.0021 4.4481e-08 0 4.4655e-08 0 4.4658e-08 0.0021 4.4661e-08 0 4.4835e-08 0 4.4838e-08 0.0021 4.4841e-08 0 4.5015e-08 0 4.5018e-08 0.0021 4.5021e-08 0 4.5195e-08 0 4.5198e-08 0.0021 4.5201e-08 0 4.5375e-08 0 4.5378e-08 0.0021 4.5381e-08 0 4.5555e-08 0 4.5558e-08 0.0021 4.5561e-08 0 4.5735e-08 0 4.5738e-08 0.0021 4.5741e-08 0 4.5915e-08 0 4.5918e-08 0.0021 4.5921e-08 0)
ISPL_IG0_0|B1 0 SPL_IG0_0|3  PWL(0 0 5e-12 0.000175)
ISPL_IG0_0|B2 0 SPL_IG0_0|6  PWL(0 0 5e-12 0.00028)
ISPL_IG0_0|B3 0 SPL_IG0_0|10  PWL(0 0 5e-12 0.000175)
ISPL_IG0_0|B4 0 SPL_IG0_0|13  PWL(0 0 5e-12 0.000175)
LSPL_IG0_0|B1 SPL_IG0_0|3 SPL_IG0_0|1  9.175e-13
LSPL_IG0_0|B2 SPL_IG0_0|6 SPL_IG0_0|4  7.666e-13
LSPL_IG0_0|B3 SPL_IG0_0|10 SPL_IG0_0|8  1.928e-12
LSPL_IG0_0|B4 SPL_IG0_0|13 SPL_IG0_0|11  8.786e-13
BSPL_IG0_0|1 SPL_IG0_0|1 SPL_IG0_0|2 JJMIT AREA=2.5
BSPL_IG0_0|2 SPL_IG0_0|4 SPL_IG0_0|5 JJMIT AREA=3.0
BSPL_IG0_0|3 SPL_IG0_0|8 SPL_IG0_0|9 JJMIT AREA=2.5
BSPL_IG0_0|4 SPL_IG0_0|11 SPL_IG0_0|12 JJMIT AREA=2.5
LSPL_IG0_0|1 IG0_0_RX SPL_IG0_0|1  2.063e-12
LSPL_IG0_0|2 SPL_IG0_0|1 SPL_IG0_0|4  3.637e-12
LSPL_IG0_0|3 SPL_IG0_0|4 SPL_IG0_0|7  1.278e-12
LSPL_IG0_0|4 SPL_IG0_0|7 SPL_IG0_0|8  1.305e-12
LSPL_IG0_0|5 SPL_IG0_0|8 IG0_0_TO0  2.05e-12
LSPL_IG0_0|6 SPL_IG0_0|7 SPL_IG0_0|11  1.315e-12
LSPL_IG0_0|7 SPL_IG0_0|11 IG0_0_TO1  2.06e-12
LSPL_IG0_0|P1 SPL_IG0_0|2 0  4.676e-13
LSPL_IG0_0|P2 SPL_IG0_0|5 0  4.498e-13
LSPL_IG0_0|P3 SPL_IG0_0|9 0  5.183e-13
LSPL_IG0_0|P4 SPL_IG0_0|12 0  4.639e-13
RSPL_IG0_0|B1 SPL_IG0_0|1 SPL_IG0_0|101  2.7439617672
LSPL_IG0_0|RB1 SPL_IG0_0|101 0  1.550338398468e-12
RSPL_IG0_0|B2 SPL_IG0_0|4 SPL_IG0_0|104  2.286634806
LSPL_IG0_0|RB2 SPL_IG0_0|104 0  1.29194866539e-12
RSPL_IG0_0|B3 SPL_IG0_0|8 SPL_IG0_0|108  2.7439617672
LSPL_IG0_0|RB3 SPL_IG0_0|108 0  1.550338398468e-12
RSPL_IG0_0|B4 SPL_IG0_0|11 SPL_IG0_0|111  2.7439617672
LSPL_IG0_0|RB4 SPL_IG0_0|111 0  1.550338398468e-12
ISPL_IP1_0|B1 0 SPL_IP1_0|3  PWL(0 0 5e-12 0.000175)
ISPL_IP1_0|B2 0 SPL_IP1_0|6  PWL(0 0 5e-12 0.00028)
ISPL_IP1_0|B3 0 SPL_IP1_0|10  PWL(0 0 5e-12 0.000175)
ISPL_IP1_0|B4 0 SPL_IP1_0|13  PWL(0 0 5e-12 0.000175)
LSPL_IP1_0|B1 SPL_IP1_0|3 SPL_IP1_0|1  9.175e-13
LSPL_IP1_0|B2 SPL_IP1_0|6 SPL_IP1_0|4  7.666e-13
LSPL_IP1_0|B3 SPL_IP1_0|10 SPL_IP1_0|8  1.928e-12
LSPL_IP1_0|B4 SPL_IP1_0|13 SPL_IP1_0|11  8.786e-13
BSPL_IP1_0|1 SPL_IP1_0|1 SPL_IP1_0|2 JJMIT AREA=2.5
BSPL_IP1_0|2 SPL_IP1_0|4 SPL_IP1_0|5 JJMIT AREA=3.0
BSPL_IP1_0|3 SPL_IP1_0|8 SPL_IP1_0|9 JJMIT AREA=2.5
BSPL_IP1_0|4 SPL_IP1_0|11 SPL_IP1_0|12 JJMIT AREA=2.5
LSPL_IP1_0|1 IP1_0_RX SPL_IP1_0|1  2.063e-12
LSPL_IP1_0|2 SPL_IP1_0|1 SPL_IP1_0|4  3.637e-12
LSPL_IP1_0|3 SPL_IP1_0|4 SPL_IP1_0|7  1.278e-12
LSPL_IP1_0|4 SPL_IP1_0|7 SPL_IP1_0|8  1.305e-12
LSPL_IP1_0|5 SPL_IP1_0|8 IP1_0_TO1  2.05e-12
LSPL_IP1_0|6 SPL_IP1_0|7 SPL_IP1_0|11  1.315e-12
LSPL_IP1_0|7 SPL_IP1_0|11 IP1_0_OUT  2.06e-12
LSPL_IP1_0|P1 SPL_IP1_0|2 0  4.676e-13
LSPL_IP1_0|P2 SPL_IP1_0|5 0  4.498e-13
LSPL_IP1_0|P3 SPL_IP1_0|9 0  5.183e-13
LSPL_IP1_0|P4 SPL_IP1_0|12 0  4.639e-13
RSPL_IP1_0|B1 SPL_IP1_0|1 SPL_IP1_0|101  2.7439617672
LSPL_IP1_0|RB1 SPL_IP1_0|101 0  1.550338398468e-12
RSPL_IP1_0|B2 SPL_IP1_0|4 SPL_IP1_0|104  2.286634806
LSPL_IP1_0|RB2 SPL_IP1_0|104 0  1.29194866539e-12
RSPL_IP1_0|B3 SPL_IP1_0|8 SPL_IP1_0|108  2.7439617672
LSPL_IP1_0|RB3 SPL_IP1_0|108 0  1.550338398468e-12
RSPL_IP1_0|B4 SPL_IP1_0|11 SPL_IP1_0|111  2.7439617672
LSPL_IP1_0|RB4 SPL_IP1_0|111 0  1.550338398468e-12
ISPL_IG2_0|B1 0 SPL_IG2_0|3  PWL(0 0 5e-12 0.000175)
ISPL_IG2_0|B2 0 SPL_IG2_0|6  PWL(0 0 5e-12 0.00028)
ISPL_IG2_0|B3 0 SPL_IG2_0|10  PWL(0 0 5e-12 0.000175)
ISPL_IG2_0|B4 0 SPL_IG2_0|13  PWL(0 0 5e-12 0.000175)
LSPL_IG2_0|B1 SPL_IG2_0|3 SPL_IG2_0|1  9.175e-13
LSPL_IG2_0|B2 SPL_IG2_0|6 SPL_IG2_0|4  7.666e-13
LSPL_IG2_0|B3 SPL_IG2_0|10 SPL_IG2_0|8  1.928e-12
LSPL_IG2_0|B4 SPL_IG2_0|13 SPL_IG2_0|11  8.786e-13
BSPL_IG2_0|1 SPL_IG2_0|1 SPL_IG2_0|2 JJMIT AREA=2.5
BSPL_IG2_0|2 SPL_IG2_0|4 SPL_IG2_0|5 JJMIT AREA=3.0
BSPL_IG2_0|3 SPL_IG2_0|8 SPL_IG2_0|9 JJMIT AREA=2.5
BSPL_IG2_0|4 SPL_IG2_0|11 SPL_IG2_0|12 JJMIT AREA=2.5
LSPL_IG2_0|1 IG2_0_RX SPL_IG2_0|1  2.063e-12
LSPL_IG2_0|2 SPL_IG2_0|1 SPL_IG2_0|4  3.637e-12
LSPL_IG2_0|3 SPL_IG2_0|4 SPL_IG2_0|7  1.278e-12
LSPL_IG2_0|4 SPL_IG2_0|7 SPL_IG2_0|8  1.305e-12
LSPL_IG2_0|5 SPL_IG2_0|8 IG2_0_TO2  2.05e-12
LSPL_IG2_0|6 SPL_IG2_0|7 SPL_IG2_0|11  1.315e-12
LSPL_IG2_0|7 SPL_IG2_0|11 IG2_0_TO3  2.06e-12
LSPL_IG2_0|P1 SPL_IG2_0|2 0  4.676e-13
LSPL_IG2_0|P2 SPL_IG2_0|5 0  4.498e-13
LSPL_IG2_0|P3 SPL_IG2_0|9 0  5.183e-13
LSPL_IG2_0|P4 SPL_IG2_0|12 0  4.639e-13
RSPL_IG2_0|B1 SPL_IG2_0|1 SPL_IG2_0|101  2.7439617672
LSPL_IG2_0|RB1 SPL_IG2_0|101 0  1.550338398468e-12
RSPL_IG2_0|B2 SPL_IG2_0|4 SPL_IG2_0|104  2.286634806
LSPL_IG2_0|RB2 SPL_IG2_0|104 0  1.29194866539e-12
RSPL_IG2_0|B3 SPL_IG2_0|8 SPL_IG2_0|108  2.7439617672
LSPL_IG2_0|RB3 SPL_IG2_0|108 0  1.550338398468e-12
RSPL_IG2_0|B4 SPL_IG2_0|11 SPL_IG2_0|111  2.7439617672
LSPL_IG2_0|RB4 SPL_IG2_0|111 0  1.550338398468e-12
ISPL_IP3_0|B1 0 SPL_IP3_0|3  PWL(0 0 5e-12 0.000175)
ISPL_IP3_0|B2 0 SPL_IP3_0|6  PWL(0 0 5e-12 0.00028)
ISPL_IP3_0|B3 0 SPL_IP3_0|10  PWL(0 0 5e-12 0.000175)
ISPL_IP3_0|B4 0 SPL_IP3_0|13  PWL(0 0 5e-12 0.000175)
LSPL_IP3_0|B1 SPL_IP3_0|3 SPL_IP3_0|1  9.175e-13
LSPL_IP3_0|B2 SPL_IP3_0|6 SPL_IP3_0|4  7.666e-13
LSPL_IP3_0|B3 SPL_IP3_0|10 SPL_IP3_0|8  1.928e-12
LSPL_IP3_0|B4 SPL_IP3_0|13 SPL_IP3_0|11  8.786e-13
BSPL_IP3_0|1 SPL_IP3_0|1 SPL_IP3_0|2 JJMIT AREA=2.5
BSPL_IP3_0|2 SPL_IP3_0|4 SPL_IP3_0|5 JJMIT AREA=3.0
BSPL_IP3_0|3 SPL_IP3_0|8 SPL_IP3_0|9 JJMIT AREA=2.5
BSPL_IP3_0|4 SPL_IP3_0|11 SPL_IP3_0|12 JJMIT AREA=2.5
LSPL_IP3_0|1 IP3_0_RX SPL_IP3_0|1  2.063e-12
LSPL_IP3_0|2 SPL_IP3_0|1 SPL_IP3_0|4  3.637e-12
LSPL_IP3_0|3 SPL_IP3_0|4 SPL_IP3_0|7  1.278e-12
LSPL_IP3_0|4 SPL_IP3_0|7 SPL_IP3_0|8  1.305e-12
LSPL_IP3_0|5 SPL_IP3_0|8 IP3_0_TO1  2.05e-12
LSPL_IP3_0|6 SPL_IP3_0|7 SPL_IP3_0|11  1.315e-12
LSPL_IP3_0|7 SPL_IP3_0|11 IP3_0_OUT  2.06e-12
LSPL_IP3_0|P1 SPL_IP3_0|2 0  4.676e-13
LSPL_IP3_0|P2 SPL_IP3_0|5 0  4.498e-13
LSPL_IP3_0|P3 SPL_IP3_0|9 0  5.183e-13
LSPL_IP3_0|P4 SPL_IP3_0|12 0  4.639e-13
RSPL_IP3_0|B1 SPL_IP3_0|1 SPL_IP3_0|101  2.7439617672
LSPL_IP3_0|RB1 SPL_IP3_0|101 0  1.550338398468e-12
RSPL_IP3_0|B2 SPL_IP3_0|4 SPL_IP3_0|104  2.286634806
LSPL_IP3_0|RB2 SPL_IP3_0|104 0  1.29194866539e-12
RSPL_IP3_0|B3 SPL_IP3_0|8 SPL_IP3_0|108  2.7439617672
LSPL_IP3_0|RB3 SPL_IP3_0|108 0  1.550338398468e-12
RSPL_IP3_0|B4 SPL_IP3_0|11 SPL_IP3_0|111  2.7439617672
LSPL_IP3_0|RB4 SPL_IP3_0|111 0  1.550338398468e-12
IT04|T 0 T04  PWL(0 0 1.05e-11 0 1.35e-11 0.0014 1.65e-11 0 1.905e-10 0 1.935e-10 0.0014 1.965e-10 0 3.705e-10 0 3.735e-10 0.0014 3.765e-10 0 5.505e-10 0 5.535e-10 0.0014 5.565e-10 0 7.305e-10 0 7.335e-10 0.0014 7.365e-10 0 9.105e-10 0 9.135e-10 0.0014 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0014 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0014 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0014 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0014 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0014 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0014 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0014 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0014 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0014 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0014 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0014 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0014 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0014 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0014 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0014 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0014 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0014 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0014 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0014 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0014 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0014 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0014 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0014 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0014 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0014 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0014 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0014 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0014 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0014 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0014 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0014 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0014 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0014 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0014 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0014 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0014 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0014 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0014 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0014 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0014 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0014 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0014 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0014 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0014 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0014 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0014 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0014 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0014 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0014 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0014 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0014 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0014 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0014 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0014 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0014 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0014 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0014 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0014 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0014 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0014 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0014 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0014 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0014 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0014 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0014 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0014 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0014 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0014 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0014 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0014 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0014 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0014 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0014 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0014 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0014 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0014 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0014 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0014 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0014 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0014 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0014 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0014 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0014 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0014 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0014 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0014 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0014 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0014 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0014 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0014 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0014 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0014 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0014 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0014 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0014 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0014 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0014 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0014 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0014 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0014 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0014 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0014 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0014 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0014 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0014 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0014 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0014 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0014 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0014 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0014 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0014 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0014 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0014 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0014 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0014 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0014 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0014 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0014 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0014 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0014 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0014 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0014 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0014 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0014 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0014 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0014 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0014 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0014 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0014 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0014 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0014 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0014 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0014 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0014 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0014 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0014 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0014 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0014 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0014 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0014 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0014 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0014 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0014 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0014 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0014 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0014 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0014 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0014 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0014 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0014 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0014 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0014 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0014 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0014 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0014 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0014 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0014 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0014 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0014 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0014 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0014 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0014 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0014 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0014 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0014 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0014 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0014 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0014 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0014 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0014 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0014 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0014 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0014 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0014 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0014 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0014 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0014 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0014 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0014 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0014 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0014 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0014 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0014 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0014 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0014 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0014 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0014 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0014 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0014 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0014 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0014 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0014 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0014 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0014 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0014 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0014 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0014 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0014 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0014 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0014 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0014 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0014 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0014 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0014 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0014 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0014 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0014 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0014 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0014 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0014 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0014 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0014 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0014 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0014 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0014 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0014 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0014 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0014 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0014 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0014 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0014 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0014 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0014 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0014 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0014 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0014 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0014 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0014 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0014 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0014 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0014 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0014 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0014 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0014 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0014 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0014 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0014 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0014 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0014 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0014 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0014 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0014 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0014 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0014 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0014 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0014 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0014 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0014 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0014 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0014 4.59165e-08 0)
IT05|T 0 T05  PWL(0 0 1.05e-11 0 1.35e-11 0.0014 1.65e-11 0 1.905e-10 0 1.935e-10 0.0014 1.965e-10 0 3.705e-10 0 3.735e-10 0.0014 3.765e-10 0 5.505e-10 0 5.535e-10 0.0014 5.565e-10 0 7.305e-10 0 7.335e-10 0.0014 7.365e-10 0 9.105e-10 0 9.135e-10 0.0014 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0014 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0014 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0014 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0014 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0014 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0014 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0014 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0014 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0014 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0014 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0014 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0014 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0014 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0014 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0014 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0014 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0014 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0014 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0014 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0014 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0014 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0014 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0014 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0014 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0014 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0014 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0014 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0014 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0014 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0014 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0014 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0014 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0014 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0014 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0014 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0014 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0014 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0014 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0014 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0014 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0014 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0014 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0014 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0014 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0014 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0014 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0014 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0014 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0014 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0014 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0014 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0014 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0014 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0014 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0014 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0014 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0014 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0014 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0014 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0014 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0014 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0014 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0014 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0014 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0014 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0014 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0014 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0014 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0014 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0014 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0014 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0014 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0014 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0014 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0014 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0014 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0014 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0014 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0014 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0014 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0014 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0014 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0014 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0014 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0014 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0014 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0014 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0014 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0014 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0014 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0014 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0014 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0014 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0014 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0014 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0014 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0014 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0014 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0014 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0014 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0014 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0014 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0014 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0014 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0014 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0014 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0014 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0014 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0014 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0014 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0014 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0014 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0014 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0014 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0014 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0014 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0014 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0014 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0014 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0014 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0014 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0014 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0014 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0014 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0014 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0014 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0014 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0014 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0014 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0014 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0014 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0014 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0014 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0014 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0014 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0014 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0014 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0014 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0014 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0014 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0014 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0014 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0014 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0014 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0014 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0014 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0014 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0014 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0014 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0014 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0014 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0014 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0014 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0014 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0014 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0014 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0014 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0014 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0014 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0014 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0014 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0014 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0014 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0014 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0014 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0014 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0014 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0014 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0014 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0014 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0014 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0014 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0014 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0014 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0014 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0014 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0014 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0014 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0014 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0014 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0014 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0014 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0014 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0014 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0014 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0014 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0014 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0014 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0014 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0014 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0014 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0014 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0014 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0014 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0014 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0014 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0014 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0014 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0014 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0014 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0014 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0014 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0014 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0014 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0014 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0014 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0014 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0014 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0014 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0014 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0014 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0014 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0014 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0014 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0014 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0014 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0014 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0014 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0014 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0014 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0014 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0014 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0014 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0014 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0014 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0014 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0014 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0014 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0014 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0014 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0014 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0014 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0014 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0014 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0014 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0014 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0014 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0014 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0014 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0014 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0014 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0014 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0014 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0014 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0014 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0014 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0014 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0014 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0014 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0014 4.59165e-08 0)
IT06|T 0 T06  PWL(0 0 1.05e-11 0 1.35e-11 0.0014 1.65e-11 0 1.905e-10 0 1.935e-10 0.0014 1.965e-10 0 3.705e-10 0 3.735e-10 0.0014 3.765e-10 0 5.505e-10 0 5.535e-10 0.0014 5.565e-10 0 7.305e-10 0 7.335e-10 0.0014 7.365e-10 0 9.105e-10 0 9.135e-10 0.0014 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0014 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0014 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0014 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0014 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0014 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0014 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0014 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0014 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0014 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0014 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0014 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0014 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0014 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0014 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0014 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0014 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0014 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0014 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0014 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0014 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0014 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0014 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0014 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0014 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0014 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0014 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0014 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0014 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0014 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0014 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0014 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0014 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0014 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0014 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0014 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0014 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0014 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0014 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0014 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0014 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0014 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0014 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0014 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0014 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0014 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0014 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0014 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0014 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0014 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0014 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0014 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0014 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0014 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0014 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0014 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0014 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0014 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0014 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0014 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0014 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0014 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0014 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0014 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0014 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0014 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0014 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0014 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0014 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0014 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0014 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0014 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0014 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0014 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0014 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0014 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0014 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0014 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0014 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0014 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0014 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0014 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0014 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0014 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0014 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0014 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0014 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0014 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0014 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0014 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0014 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0014 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0014 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0014 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0014 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0014 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0014 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0014 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0014 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0014 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0014 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0014 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0014 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0014 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0014 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0014 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0014 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0014 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0014 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0014 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0014 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0014 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0014 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0014 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0014 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0014 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0014 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0014 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0014 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0014 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0014 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0014 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0014 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0014 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0014 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0014 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0014 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0014 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0014 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0014 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0014 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0014 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0014 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0014 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0014 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0014 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0014 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0014 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0014 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0014 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0014 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0014 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0014 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0014 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0014 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0014 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0014 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0014 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0014 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0014 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0014 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0014 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0014 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0014 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0014 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0014 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0014 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0014 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0014 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0014 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0014 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0014 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0014 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0014 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0014 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0014 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0014 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0014 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0014 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0014 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0014 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0014 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0014 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0014 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0014 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0014 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0014 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0014 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0014 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0014 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0014 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0014 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0014 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0014 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0014 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0014 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0014 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0014 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0014 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0014 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0014 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0014 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0014 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0014 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0014 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0014 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0014 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0014 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0014 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0014 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0014 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0014 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0014 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0014 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0014 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0014 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0014 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0014 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0014 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0014 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0014 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0014 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0014 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0014 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0014 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0014 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0014 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0014 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0014 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0014 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0014 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0014 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0014 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0014 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0014 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0014 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0014 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0014 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0014 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0014 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0014 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0014 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0014 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0014 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0014 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0014 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0014 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0014 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0014 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0014 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0014 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0014 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0014 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0014 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0014 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0014 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0014 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0014 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0014 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0014 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0014 4.59165e-08 0)
IT07|T 0 T07  PWL(0 0 1.05e-11 0 1.35e-11 0.0028 1.65e-11 0 1.905e-10 0 1.935e-10 0.0028 1.965e-10 0 3.705e-10 0 3.735e-10 0.0028 3.765e-10 0 5.505e-10 0 5.535e-10 0.0028 5.565e-10 0 7.305e-10 0 7.335e-10 0.0028 7.365e-10 0 9.105e-10 0 9.135e-10 0.0028 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0028 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0028 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0028 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0028 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0028 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0028 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0028 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0028 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0028 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0028 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0028 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0028 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0028 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0028 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0028 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0028 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0028 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0028 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0028 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0028 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0028 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0028 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0028 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0028 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0028 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0028 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0028 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0028 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0028 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0028 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0028 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0028 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0028 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0028 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0028 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0028 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0028 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0028 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0028 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0028 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0028 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0028 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0028 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0028 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0028 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0028 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0028 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0028 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0028 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0028 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0028 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0028 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0028 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0028 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0028 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0028 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0028 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0028 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0028 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0028 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0028 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0028 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0028 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0028 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0028 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0028 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0028 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0028 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0028 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0028 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0028 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0028 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0028 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0028 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0028 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0028 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0028 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0028 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0028 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0028 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0028 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0028 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0028 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0028 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0028 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0028 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0028 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0028 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0028 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0028 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0028 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0028 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0028 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0028 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0028 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0028 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0028 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0028 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0028 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0028 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0028 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0028 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0028 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0028 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0028 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0028 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0028 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0028 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0028 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0028 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0028 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0028 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0028 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0028 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0028 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0028 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0028 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0028 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0028 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0028 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0028 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0028 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0028 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0028 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0028 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0028 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0028 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0028 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0028 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0028 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0028 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0028 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0028 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0028 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0028 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0028 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0028 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0028 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0028 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0028 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0028 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0028 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0028 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0028 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0028 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0028 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0028 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0028 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0028 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0028 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0028 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0028 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0028 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0028 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0028 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0028 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0028 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0028 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0028 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0028 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0028 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0028 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0028 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0028 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0028 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0028 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0028 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0028 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0028 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0028 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0028 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0028 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0028 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0028 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0028 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0028 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0028 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0028 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0028 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0028 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0028 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0028 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0028 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0028 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0028 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0028 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0028 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0028 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0028 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0028 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0028 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0028 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0028 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0028 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0028 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0028 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0028 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0028 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0028 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0028 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0028 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0028 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0028 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0028 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0028 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0028 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0028 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0028 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0028 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0028 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0028 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0028 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0028 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0028 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0028 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0028 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0028 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0028 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0028 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0028 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0028 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0028 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0028 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0028 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0028 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0028 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0028 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0028 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0028 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0028 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0028 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0028 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0028 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0028 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0028 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0028 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0028 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0028 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0028 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0028 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0028 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0028 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0028 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0028 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0028 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0028 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0028 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0028 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0028 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0028 4.59165e-08 0)
ID01|T 0 D01  PWL(0 0 1.05e-11 0 1.35e-11 0.0007 1.65e-11 0 1.905e-10 0 1.935e-10 0.0007 1.965e-10 0 3.705e-10 0 3.735e-10 0.0007 3.765e-10 0 5.505e-10 0 5.535e-10 0.0007 5.565e-10 0 7.305e-10 0 7.335e-10 0.0007 7.365e-10 0 9.105e-10 0 9.135e-10 0.0007 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0007 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0007 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0007 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0007 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0007 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0007 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0007 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0007 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0007 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0007 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0007 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0007 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0007 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0007 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0007 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0007 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0007 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0007 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0007 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0007 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0007 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0007 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0007 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0007 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0007 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0007 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0007 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0007 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0007 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0007 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0007 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0007 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0007 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0007 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0007 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0007 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0007 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0007 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0007 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0007 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0007 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0007 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0007 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0007 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0007 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0007 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0007 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0007 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0007 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0007 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0007 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0007 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0007 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0007 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0007 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0007 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0007 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0007 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0007 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0007 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0007 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0007 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0007 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0007 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0007 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0007 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0007 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0007 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0007 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0007 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0007 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0007 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0007 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0007 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0007 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0007 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0007 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0007 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0007 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0007 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0007 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0007 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0007 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0007 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0007 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0007 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0007 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0007 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0007 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0007 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0007 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0007 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0007 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0007 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0007 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0007 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0007 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0007 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0007 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0007 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0007 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0007 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0007 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0007 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0007 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0007 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0007 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0007 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0007 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0007 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0007 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0007 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0007 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0007 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0007 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0007 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0007 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0007 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0007 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0007 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0007 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0007 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0007 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0007 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0007 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0007 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0007 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0007 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0007 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0007 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0007 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0007 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0007 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0007 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0007 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0007 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0007 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0007 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0007 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0007 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0007 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0007 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0007 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0007 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0007 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0007 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0007 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0007 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0007 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0007 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0007 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0007 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0007 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0007 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0007 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0007 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0007 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0007 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0007 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0007 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0007 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0007 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0007 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0007 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0007 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0007 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0007 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0007 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0007 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0007 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0007 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0007 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0007 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0007 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0007 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0007 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0007 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0007 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0007 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0007 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0007 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0007 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0007 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0007 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0007 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0007 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0007 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0007 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0007 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0007 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0007 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0007 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0007 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0007 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0007 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0007 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0007 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0007 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0007 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0007 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0007 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0007 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0007 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0007 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0007 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0007 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0007 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0007 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0007 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0007 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0007 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0007 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0007 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0007 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0007 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0007 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0007 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0007 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0007 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0007 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0007 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0007 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0007 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0007 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0007 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0007 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0007 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0007 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0007 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0007 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0007 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0007 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0007 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0007 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0007 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0007 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0007 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0007 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0007 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0007 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0007 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0007 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0007 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0007 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0007 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0007 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0007 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0007 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0007 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0007 4.59165e-08 0)
B_DFF_IP1_01|1 _DFF_IP1_01|1 _DFF_IP1_01|2 JJMIT AREA=2.5
B_DFF_IP1_01|2 _DFF_IP1_01|4 _DFF_IP1_01|5 JJMIT AREA=1.61
B_DFF_IP1_01|3 _DFF_IP1_01|5 _DFF_IP1_01|6 JJMIT AREA=1.54
B_DFF_IP1_01|4 _DFF_IP1_01|8 _DFF_IP1_01|9 JJMIT AREA=1.69
B_DFF_IP1_01|5 _DFF_IP1_01|10 _DFF_IP1_01|8 JJMIT AREA=1.38
B_DFF_IP1_01|6 _DFF_IP1_01|11 _DFF_IP1_01|12 JJMIT AREA=2.5
B_DFF_IP1_01|7 _DFF_IP1_01|14 _DFF_IP1_01|15 JJMIT AREA=2.5
I_DFF_IP1_01|B1 0 _DFF_IP1_01|3  PWL(0 0 5e-12 0.000175)
I_DFF_IP1_01|B2 0 _DFF_IP1_01|7  PWL(0 0 5e-12 0.000173)
I_DFF_IP1_01|B3 0 _DFF_IP1_01|13  PWL(0 0 5e-12 0.000175)
I_DFF_IP1_01|B4 0 _DFF_IP1_01|16  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|B1 _DFF_IP1_01|3 _DFF_IP1_01|1  2e-12
L_DFF_IP1_01|B2 _DFF_IP1_01|7 _DFF_IP1_01|5  2e-12
L_DFF_IP1_01|B3 _DFF_IP1_01|11 _DFF_IP1_01|13  2e-12
L_DFF_IP1_01|B4 _DFF_IP1_01|16 _DFF_IP1_01|14  2e-12
L_DFF_IP1_01|1 IP1_0_OUT _DFF_IP1_01|1  2.059e-12
L_DFF_IP1_01|2 _DFF_IP1_01|1 _DFF_IP1_01|4  4.123e-12
L_DFF_IP1_01|3 _DFF_IP1_01|5 _DFF_IP1_01|8  6.873e-12
L_DFF_IP1_01|4 _DFF_IP1_01|10 _DFF_IP1_01|11  5.195e-12
L_DFF_IP1_01|5 D01 _DFF_IP1_01|11  2.071e-12
L_DFF_IP1_01|6 _DFF_IP1_01|8 _DFF_IP1_01|14  3.287e-12
L_DFF_IP1_01|7 _DFF_IP1_01|14 IP1_1_OUT  2.066e-12
L_DFF_IP1_01|P1 _DFF_IP1_01|2 0  5.042e-13
L_DFF_IP1_01|P3 _DFF_IP1_01|6 0  5.799e-13
L_DFF_IP1_01|P4 _DFF_IP1_01|9 0  5.733e-13
L_DFF_IP1_01|P6 _DFF_IP1_01|12 0  4.605e-13
L_DFF_IP1_01|P7 _DFF_IP1_01|15 0  4.961e-13
R_DFF_IP1_01|B1 _DFF_IP1_01|1 _DFF_IP1_01|101  2.7439617672
L_DFF_IP1_01|RB1 _DFF_IP1_01|101 0  1.550338398468e-12
R_DFF_IP1_01|B2 _DFF_IP1_01|4 _DFF_IP1_01|104  4.260810197515528
L_DFF_IP1_01|RB2 _DFF_IP1_01|104 _DFF_IP1_01|5  2.407357761596273e-12
R_DFF_IP1_01|B3 _DFF_IP1_01|5 _DFF_IP1_01|105  4.454483388311688
L_DFF_IP1_01|RB3 _DFF_IP1_01|105 0  2.516783114396104e-12
R_DFF_IP1_01|B4 _DFF_IP1_01|8 _DFF_IP1_01|108  4.059115040236686
L_DFF_IP1_01|RB4 _DFF_IP1_01|108 0  2.2933999977337278e-12
R_DFF_IP1_01|B5 _DFF_IP1_01|10 _DFF_IP1_01|110  4.970945230434783
L_DFF_IP1_01|RB5 _DFF_IP1_01|110 _DFF_IP1_01|8  2.8085840551956523e-12
R_DFF_IP1_01|B6 _DFF_IP1_01|11 _DFF_IP1_01|111  2.7439617672
L_DFF_IP1_01|RB6 _DFF_IP1_01|111 0  1.550338398468e-12
R_DFF_IP1_01|B7 _DFF_IP1_01|14 _DFF_IP1_01|114  2.7439617672
L_DFF_IP1_01|RB7 _DFF_IP1_01|114 0  1.550338398468e-12
ID02|T 0 D02  PWL(0 0 1.05e-11 0 1.35e-11 0.0007 1.65e-11 0 1.905e-10 0 1.935e-10 0.0007 1.965e-10 0 3.705e-10 0 3.735e-10 0.0007 3.765e-10 0 5.505e-10 0 5.535e-10 0.0007 5.565e-10 0 7.305e-10 0 7.335e-10 0.0007 7.365e-10 0 9.105e-10 0 9.135e-10 0.0007 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0007 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0007 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0007 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0007 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0007 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0007 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0007 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0007 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0007 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0007 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0007 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0007 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0007 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0007 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0007 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0007 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0007 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0007 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0007 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0007 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0007 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0007 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0007 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0007 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0007 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0007 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0007 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0007 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0007 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0007 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0007 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0007 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0007 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0007 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0007 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0007 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0007 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0007 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0007 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0007 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0007 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0007 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0007 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0007 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0007 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0007 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0007 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0007 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0007 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0007 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0007 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0007 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0007 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0007 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0007 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0007 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0007 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0007 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0007 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0007 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0007 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0007 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0007 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0007 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0007 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0007 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0007 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0007 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0007 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0007 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0007 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0007 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0007 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0007 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0007 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0007 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0007 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0007 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0007 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0007 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0007 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0007 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0007 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0007 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0007 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0007 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0007 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0007 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0007 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0007 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0007 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0007 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0007 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0007 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0007 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0007 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0007 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0007 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0007 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0007 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0007 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0007 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0007 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0007 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0007 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0007 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0007 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0007 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0007 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0007 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0007 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0007 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0007 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0007 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0007 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0007 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0007 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0007 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0007 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0007 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0007 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0007 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0007 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0007 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0007 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0007 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0007 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0007 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0007 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0007 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0007 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0007 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0007 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0007 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0007 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0007 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0007 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0007 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0007 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0007 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0007 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0007 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0007 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0007 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0007 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0007 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0007 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0007 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0007 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0007 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0007 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0007 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0007 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0007 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0007 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0007 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0007 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0007 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0007 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0007 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0007 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0007 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0007 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0007 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0007 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0007 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0007 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0007 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0007 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0007 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0007 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0007 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0007 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0007 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0007 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0007 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0007 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0007 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0007 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0007 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0007 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0007 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0007 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0007 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0007 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0007 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0007 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0007 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0007 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0007 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0007 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0007 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0007 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0007 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0007 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0007 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0007 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0007 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0007 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0007 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0007 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0007 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0007 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0007 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0007 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0007 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0007 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0007 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0007 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0007 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0007 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0007 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0007 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0007 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0007 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0007 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0007 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0007 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0007 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0007 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0007 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0007 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0007 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0007 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0007 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0007 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0007 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0007 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0007 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0007 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0007 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0007 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0007 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0007 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0007 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0007 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0007 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0007 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0007 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0007 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0007 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0007 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0007 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0007 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0007 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0007 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0007 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0007 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0007 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0007 4.59165e-08 0)
B_DFF_IP2_01|1 _DFF_IP2_01|1 _DFF_IP2_01|2 JJMIT AREA=2.5
B_DFF_IP2_01|2 _DFF_IP2_01|4 _DFF_IP2_01|5 JJMIT AREA=1.61
B_DFF_IP2_01|3 _DFF_IP2_01|5 _DFF_IP2_01|6 JJMIT AREA=1.54
B_DFF_IP2_01|4 _DFF_IP2_01|8 _DFF_IP2_01|9 JJMIT AREA=1.69
B_DFF_IP2_01|5 _DFF_IP2_01|10 _DFF_IP2_01|8 JJMIT AREA=1.38
B_DFF_IP2_01|6 _DFF_IP2_01|11 _DFF_IP2_01|12 JJMIT AREA=2.5
B_DFF_IP2_01|7 _DFF_IP2_01|14 _DFF_IP2_01|15 JJMIT AREA=2.5
I_DFF_IP2_01|B1 0 _DFF_IP2_01|3  PWL(0 0 5e-12 0.000175)
I_DFF_IP2_01|B2 0 _DFF_IP2_01|7  PWL(0 0 5e-12 0.000173)
I_DFF_IP2_01|B3 0 _DFF_IP2_01|13  PWL(0 0 5e-12 0.000175)
I_DFF_IP2_01|B4 0 _DFF_IP2_01|16  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|B1 _DFF_IP2_01|3 _DFF_IP2_01|1  2e-12
L_DFF_IP2_01|B2 _DFF_IP2_01|7 _DFF_IP2_01|5  2e-12
L_DFF_IP2_01|B3 _DFF_IP2_01|11 _DFF_IP2_01|13  2e-12
L_DFF_IP2_01|B4 _DFF_IP2_01|16 _DFF_IP2_01|14  2e-12
L_DFF_IP2_01|1 IP2_0_OUT _DFF_IP2_01|1  2.059e-12
L_DFF_IP2_01|2 _DFF_IP2_01|1 _DFF_IP2_01|4  4.123e-12
L_DFF_IP2_01|3 _DFF_IP2_01|5 _DFF_IP2_01|8  6.873e-12
L_DFF_IP2_01|4 _DFF_IP2_01|10 _DFF_IP2_01|11  5.195e-12
L_DFF_IP2_01|5 D02 _DFF_IP2_01|11  2.071e-12
L_DFF_IP2_01|6 _DFF_IP2_01|8 _DFF_IP2_01|14  3.287e-12
L_DFF_IP2_01|7 _DFF_IP2_01|14 IP2_1_OUT  2.066e-12
L_DFF_IP2_01|P1 _DFF_IP2_01|2 0  5.042e-13
L_DFF_IP2_01|P3 _DFF_IP2_01|6 0  5.799e-13
L_DFF_IP2_01|P4 _DFF_IP2_01|9 0  5.733e-13
L_DFF_IP2_01|P6 _DFF_IP2_01|12 0  4.605e-13
L_DFF_IP2_01|P7 _DFF_IP2_01|15 0  4.961e-13
R_DFF_IP2_01|B1 _DFF_IP2_01|1 _DFF_IP2_01|101  2.7439617672
L_DFF_IP2_01|RB1 _DFF_IP2_01|101 0  1.550338398468e-12
R_DFF_IP2_01|B2 _DFF_IP2_01|4 _DFF_IP2_01|104  4.260810197515528
L_DFF_IP2_01|RB2 _DFF_IP2_01|104 _DFF_IP2_01|5  2.407357761596273e-12
R_DFF_IP2_01|B3 _DFF_IP2_01|5 _DFF_IP2_01|105  4.454483388311688
L_DFF_IP2_01|RB3 _DFF_IP2_01|105 0  2.516783114396104e-12
R_DFF_IP2_01|B4 _DFF_IP2_01|8 _DFF_IP2_01|108  4.059115040236686
L_DFF_IP2_01|RB4 _DFF_IP2_01|108 0  2.2933999977337278e-12
R_DFF_IP2_01|B5 _DFF_IP2_01|10 _DFF_IP2_01|110  4.970945230434783
L_DFF_IP2_01|RB5 _DFF_IP2_01|110 _DFF_IP2_01|8  2.8085840551956523e-12
R_DFF_IP2_01|B6 _DFF_IP2_01|11 _DFF_IP2_01|111  2.7439617672
L_DFF_IP2_01|RB6 _DFF_IP2_01|111 0  1.550338398468e-12
R_DFF_IP2_01|B7 _DFF_IP2_01|14 _DFF_IP2_01|114  2.7439617672
L_DFF_IP2_01|RB7 _DFF_IP2_01|114 0  1.550338398468e-12
ID03|T 0 D03  PWL(0 0 1.05e-11 0 1.35e-11 0.0007 1.65e-11 0 1.905e-10 0 1.935e-10 0.0007 1.965e-10 0 3.705e-10 0 3.735e-10 0.0007 3.765e-10 0 5.505e-10 0 5.535e-10 0.0007 5.565e-10 0 7.305e-10 0 7.335e-10 0.0007 7.365e-10 0 9.105e-10 0 9.135e-10 0.0007 9.165e-10 0 1.0905e-09 0 1.0935e-09 0.0007 1.0965e-09 0 1.2705e-09 0 1.2735e-09 0.0007 1.2765e-09 0 1.4505e-09 0 1.4535e-09 0.0007 1.4565e-09 0 1.6305e-09 0 1.6335e-09 0.0007 1.6365e-09 0 1.8105e-09 0 1.8135e-09 0.0007 1.8165e-09 0 1.9905e-09 0 1.9935e-09 0.0007 1.9965e-09 0 2.1705e-09 0 2.1735e-09 0.0007 2.1765e-09 0 2.3505e-09 0 2.3535e-09 0.0007 2.3565e-09 0 2.5305e-09 0 2.5335e-09 0.0007 2.5365e-09 0 2.7105e-09 0 2.7135e-09 0.0007 2.7165e-09 0 2.8905e-09 0 2.8935e-09 0.0007 2.8965e-09 0 3.0705e-09 0 3.0735e-09 0.0007 3.0765e-09 0 3.2505e-09 0 3.2535e-09 0.0007 3.2565e-09 0 3.4305e-09 0 3.4335e-09 0.0007 3.4365e-09 0 3.6105e-09 0 3.6135e-09 0.0007 3.6165e-09 0 3.7905e-09 0 3.7935e-09 0.0007 3.7965e-09 0 3.9705e-09 0 3.9735e-09 0.0007 3.9765e-09 0 4.1505e-09 0 4.1535e-09 0.0007 4.1565e-09 0 4.3305e-09 0 4.3335e-09 0.0007 4.3365e-09 0 4.5105e-09 0 4.5135e-09 0.0007 4.5165e-09 0 4.6905e-09 0 4.6935e-09 0.0007 4.6965e-09 0 4.8705e-09 0 4.8735e-09 0.0007 4.8765e-09 0 5.0505e-09 0 5.0535e-09 0.0007 5.0565e-09 0 5.2305e-09 0 5.2335e-09 0.0007 5.2365e-09 0 5.4105e-09 0 5.4135e-09 0.0007 5.4165e-09 0 5.5905e-09 0 5.5935e-09 0.0007 5.5965e-09 0 5.7705e-09 0 5.7735e-09 0.0007 5.7765e-09 0 5.9505e-09 0 5.9535e-09 0.0007 5.9565e-09 0 6.1305e-09 0 6.1335e-09 0.0007 6.1365e-09 0 6.3105e-09 0 6.3135e-09 0.0007 6.3165e-09 0 6.4905e-09 0 6.4935e-09 0.0007 6.4965e-09 0 6.6705e-09 0 6.6735e-09 0.0007 6.6765e-09 0 6.8505e-09 0 6.8535e-09 0.0007 6.8565e-09 0 7.0305e-09 0 7.0335e-09 0.0007 7.0365e-09 0 7.2105e-09 0 7.2135e-09 0.0007 7.2165e-09 0 7.3905e-09 0 7.3935e-09 0.0007 7.3965e-09 0 7.5705e-09 0 7.5735e-09 0.0007 7.5765e-09 0 7.7505e-09 0 7.7535e-09 0.0007 7.7565e-09 0 7.9305e-09 0 7.9335e-09 0.0007 7.9365e-09 0 8.1105e-09 0 8.1135e-09 0.0007 8.1165e-09 0 8.2905e-09 0 8.2935e-09 0.0007 8.2965e-09 0 8.4705e-09 0 8.4735e-09 0.0007 8.4765e-09 0 8.6505e-09 0 8.6535e-09 0.0007 8.6565e-09 0 8.8305e-09 0 8.8335e-09 0.0007 8.8365e-09 0 9.0105e-09 0 9.0135e-09 0.0007 9.0165e-09 0 9.1905e-09 0 9.1935e-09 0.0007 9.1965e-09 0 9.3705e-09 0 9.3735e-09 0.0007 9.3765e-09 0 9.5505e-09 0 9.5535e-09 0.0007 9.5565e-09 0 9.7305e-09 0 9.7335e-09 0.0007 9.7365e-09 0 9.9105e-09 0 9.9135e-09 0.0007 9.9165e-09 0 1.00905e-08 0 1.00935e-08 0.0007 1.00965e-08 0 1.02705e-08 0 1.02735e-08 0.0007 1.02765e-08 0 1.04505e-08 0 1.04535e-08 0.0007 1.04565e-08 0 1.06305e-08 0 1.06335e-08 0.0007 1.06365e-08 0 1.08105e-08 0 1.08135e-08 0.0007 1.08165e-08 0 1.09905e-08 0 1.09935e-08 0.0007 1.09965e-08 0 1.11705e-08 0 1.11735e-08 0.0007 1.11765e-08 0 1.13505e-08 0 1.13535e-08 0.0007 1.13565e-08 0 1.15305e-08 0 1.15335e-08 0.0007 1.15365e-08 0 1.17105e-08 0 1.17135e-08 0.0007 1.17165e-08 0 1.18905e-08 0 1.18935e-08 0.0007 1.18965e-08 0 1.20705e-08 0 1.20735e-08 0.0007 1.20765e-08 0 1.22505e-08 0 1.22535e-08 0.0007 1.22565e-08 0 1.24305e-08 0 1.24335e-08 0.0007 1.24365e-08 0 1.26105e-08 0 1.26135e-08 0.0007 1.26165e-08 0 1.27905e-08 0 1.27935e-08 0.0007 1.27965e-08 0 1.29705e-08 0 1.29735e-08 0.0007 1.29765e-08 0 1.31505e-08 0 1.31535e-08 0.0007 1.31565e-08 0 1.33305e-08 0 1.33335e-08 0.0007 1.33365e-08 0 1.35105e-08 0 1.35135e-08 0.0007 1.35165e-08 0 1.36905e-08 0 1.36935e-08 0.0007 1.36965e-08 0 1.38705e-08 0 1.38735e-08 0.0007 1.38765e-08 0 1.40505e-08 0 1.40535e-08 0.0007 1.40565e-08 0 1.42305e-08 0 1.42335e-08 0.0007 1.42365e-08 0 1.44105e-08 0 1.44135e-08 0.0007 1.44165e-08 0 1.45905e-08 0 1.45935e-08 0.0007 1.45965e-08 0 1.47705e-08 0 1.47735e-08 0.0007 1.47765e-08 0 1.49505e-08 0 1.49535e-08 0.0007 1.49565e-08 0 1.51305e-08 0 1.51335e-08 0.0007 1.51365e-08 0 1.53105e-08 0 1.53135e-08 0.0007 1.53165e-08 0 1.54905e-08 0 1.54935e-08 0.0007 1.54965e-08 0 1.56705e-08 0 1.56735e-08 0.0007 1.56765e-08 0 1.58505e-08 0 1.58535e-08 0.0007 1.58565e-08 0 1.60305e-08 0 1.60335e-08 0.0007 1.60365e-08 0 1.62105e-08 0 1.62135e-08 0.0007 1.62165e-08 0 1.63905e-08 0 1.63935e-08 0.0007 1.63965e-08 0 1.65705e-08 0 1.65735e-08 0.0007 1.65765e-08 0 1.67505e-08 0 1.67535e-08 0.0007 1.67565e-08 0 1.69305e-08 0 1.69335e-08 0.0007 1.69365e-08 0 1.71105e-08 0 1.71135e-08 0.0007 1.71165e-08 0 1.72905e-08 0 1.72935e-08 0.0007 1.72965e-08 0 1.74705e-08 0 1.74735e-08 0.0007 1.74765e-08 0 1.76505e-08 0 1.76535e-08 0.0007 1.76565e-08 0 1.78305e-08 0 1.78335e-08 0.0007 1.78365e-08 0 1.80105e-08 0 1.80135e-08 0.0007 1.80165e-08 0 1.81905e-08 0 1.81935e-08 0.0007 1.81965e-08 0 1.83705e-08 0 1.83735e-08 0.0007 1.83765e-08 0 1.85505e-08 0 1.85535e-08 0.0007 1.85565e-08 0 1.87305e-08 0 1.87335e-08 0.0007 1.87365e-08 0 1.89105e-08 0 1.89135e-08 0.0007 1.89165e-08 0 1.90905e-08 0 1.90935e-08 0.0007 1.90965e-08 0 1.92705e-08 0 1.92735e-08 0.0007 1.92765e-08 0 1.94505e-08 0 1.94535e-08 0.0007 1.94565e-08 0 1.96305e-08 0 1.96335e-08 0.0007 1.96365e-08 0 1.98105e-08 0 1.98135e-08 0.0007 1.98165e-08 0 1.99905e-08 0 1.99935e-08 0.0007 1.99965e-08 0 2.01705e-08 0 2.01735e-08 0.0007 2.01765e-08 0 2.03505e-08 0 2.03535e-08 0.0007 2.03565e-08 0 2.05305e-08 0 2.05335e-08 0.0007 2.05365e-08 0 2.07105e-08 0 2.07135e-08 0.0007 2.07165e-08 0 2.08905e-08 0 2.08935e-08 0.0007 2.08965e-08 0 2.10705e-08 0 2.10735e-08 0.0007 2.10765e-08 0 2.12505e-08 0 2.12535e-08 0.0007 2.12565e-08 0 2.14305e-08 0 2.14335e-08 0.0007 2.14365e-08 0 2.16105e-08 0 2.16135e-08 0.0007 2.16165e-08 0 2.17905e-08 0 2.17935e-08 0.0007 2.17965e-08 0 2.19705e-08 0 2.19735e-08 0.0007 2.19765e-08 0 2.21505e-08 0 2.21535e-08 0.0007 2.21565e-08 0 2.23305e-08 0 2.23335e-08 0.0007 2.23365e-08 0 2.25105e-08 0 2.25135e-08 0.0007 2.25165e-08 0 2.26905e-08 0 2.26935e-08 0.0007 2.26965e-08 0 2.28705e-08 0 2.28735e-08 0.0007 2.28765e-08 0 2.30505e-08 0 2.30535e-08 0.0007 2.30565e-08 0 2.32305e-08 0 2.32335e-08 0.0007 2.32365e-08 0 2.34105e-08 0 2.34135e-08 0.0007 2.34165e-08 0 2.35905e-08 0 2.35935e-08 0.0007 2.35965e-08 0 2.37705e-08 0 2.37735e-08 0.0007 2.37765e-08 0 2.39505e-08 0 2.39535e-08 0.0007 2.39565e-08 0 2.41305e-08 0 2.41335e-08 0.0007 2.41365e-08 0 2.43105e-08 0 2.43135e-08 0.0007 2.43165e-08 0 2.44905e-08 0 2.44935e-08 0.0007 2.44965e-08 0 2.46705e-08 0 2.46735e-08 0.0007 2.46765e-08 0 2.48505e-08 0 2.48535e-08 0.0007 2.48565e-08 0 2.50305e-08 0 2.50335e-08 0.0007 2.50365e-08 0 2.52105e-08 0 2.52135e-08 0.0007 2.52165e-08 0 2.53905e-08 0 2.53935e-08 0.0007 2.53965e-08 0 2.55705e-08 0 2.55735e-08 0.0007 2.55765e-08 0 2.57505e-08 0 2.57535e-08 0.0007 2.57565e-08 0 2.59305e-08 0 2.59335e-08 0.0007 2.59365e-08 0 2.61105e-08 0 2.61135e-08 0.0007 2.61165e-08 0 2.62905e-08 0 2.62935e-08 0.0007 2.62965e-08 0 2.64705e-08 0 2.64735e-08 0.0007 2.64765e-08 0 2.66505e-08 0 2.66535e-08 0.0007 2.66565e-08 0 2.68305e-08 0 2.68335e-08 0.0007 2.68365e-08 0 2.70105e-08 0 2.70135e-08 0.0007 2.70165e-08 0 2.71905e-08 0 2.71935e-08 0.0007 2.71965e-08 0 2.73705e-08 0 2.73735e-08 0.0007 2.73765e-08 0 2.75505e-08 0 2.75535e-08 0.0007 2.75565e-08 0 2.77305e-08 0 2.77335e-08 0.0007 2.77365e-08 0 2.79105e-08 0 2.79135e-08 0.0007 2.79165e-08 0 2.80905e-08 0 2.80935e-08 0.0007 2.80965e-08 0 2.82705e-08 0 2.82735e-08 0.0007 2.82765e-08 0 2.84505e-08 0 2.84535e-08 0.0007 2.84565e-08 0 2.86305e-08 0 2.86335e-08 0.0007 2.86365e-08 0 2.88105e-08 0 2.88135e-08 0.0007 2.88165e-08 0 2.89905e-08 0 2.89935e-08 0.0007 2.89965e-08 0 2.91705e-08 0 2.91735e-08 0.0007 2.91765e-08 0 2.93505e-08 0 2.93535e-08 0.0007 2.93565e-08 0 2.95305e-08 0 2.95335e-08 0.0007 2.95365e-08 0 2.97105e-08 0 2.97135e-08 0.0007 2.97165e-08 0 2.98905e-08 0 2.98935e-08 0.0007 2.98965e-08 0 3.00705e-08 0 3.00735e-08 0.0007 3.00765e-08 0 3.02505e-08 0 3.02535e-08 0.0007 3.02565e-08 0 3.04305e-08 0 3.04335e-08 0.0007 3.04365e-08 0 3.06105e-08 0 3.06135e-08 0.0007 3.06165e-08 0 3.07905e-08 0 3.07935e-08 0.0007 3.07965e-08 0 3.09705e-08 0 3.09735e-08 0.0007 3.09765e-08 0 3.11505e-08 0 3.11535e-08 0.0007 3.11565e-08 0 3.13305e-08 0 3.13335e-08 0.0007 3.13365e-08 0 3.15105e-08 0 3.15135e-08 0.0007 3.15165e-08 0 3.16905e-08 0 3.16935e-08 0.0007 3.16965e-08 0 3.18705e-08 0 3.18735e-08 0.0007 3.18765e-08 0 3.20505e-08 0 3.20535e-08 0.0007 3.20565e-08 0 3.22305e-08 0 3.22335e-08 0.0007 3.22365e-08 0 3.24105e-08 0 3.24135e-08 0.0007 3.24165e-08 0 3.25905e-08 0 3.25935e-08 0.0007 3.25965e-08 0 3.27705e-08 0 3.27735e-08 0.0007 3.27765e-08 0 3.29505e-08 0 3.29535e-08 0.0007 3.29565e-08 0 3.31305e-08 0 3.31335e-08 0.0007 3.31365e-08 0 3.33105e-08 0 3.33135e-08 0.0007 3.33165e-08 0 3.34905e-08 0 3.34935e-08 0.0007 3.34965e-08 0 3.36705e-08 0 3.36735e-08 0.0007 3.36765e-08 0 3.38505e-08 0 3.38535e-08 0.0007 3.38565e-08 0 3.40305e-08 0 3.40335e-08 0.0007 3.40365e-08 0 3.42105e-08 0 3.42135e-08 0.0007 3.42165e-08 0 3.43905e-08 0 3.43935e-08 0.0007 3.43965e-08 0 3.45705e-08 0 3.45735e-08 0.0007 3.45765e-08 0 3.47505e-08 0 3.47535e-08 0.0007 3.47565e-08 0 3.49305e-08 0 3.49335e-08 0.0007 3.49365e-08 0 3.51105e-08 0 3.51135e-08 0.0007 3.51165e-08 0 3.52905e-08 0 3.52935e-08 0.0007 3.52965e-08 0 3.54705e-08 0 3.54735e-08 0.0007 3.54765e-08 0 3.56505e-08 0 3.56535e-08 0.0007 3.56565e-08 0 3.58305e-08 0 3.58335e-08 0.0007 3.58365e-08 0 3.60105e-08 0 3.60135e-08 0.0007 3.60165e-08 0 3.61905e-08 0 3.61935e-08 0.0007 3.61965e-08 0 3.63705e-08 0 3.63735e-08 0.0007 3.63765e-08 0 3.65505e-08 0 3.65535e-08 0.0007 3.65565e-08 0 3.67305e-08 0 3.67335e-08 0.0007 3.67365e-08 0 3.69105e-08 0 3.69135e-08 0.0007 3.69165e-08 0 3.70905e-08 0 3.70935e-08 0.0007 3.70965e-08 0 3.72705e-08 0 3.72735e-08 0.0007 3.72765e-08 0 3.74505e-08 0 3.74535e-08 0.0007 3.74565e-08 0 3.76305e-08 0 3.76335e-08 0.0007 3.76365e-08 0 3.78105e-08 0 3.78135e-08 0.0007 3.78165e-08 0 3.79905e-08 0 3.79935e-08 0.0007 3.79965e-08 0 3.81705e-08 0 3.81735e-08 0.0007 3.81765e-08 0 3.83505e-08 0 3.83535e-08 0.0007 3.83565e-08 0 3.85305e-08 0 3.85335e-08 0.0007 3.85365e-08 0 3.87105e-08 0 3.87135e-08 0.0007 3.87165e-08 0 3.88905e-08 0 3.88935e-08 0.0007 3.88965e-08 0 3.90705e-08 0 3.90735e-08 0.0007 3.90765e-08 0 3.92505e-08 0 3.92535e-08 0.0007 3.92565e-08 0 3.94305e-08 0 3.94335e-08 0.0007 3.94365e-08 0 3.96105e-08 0 3.96135e-08 0.0007 3.96165e-08 0 3.97905e-08 0 3.97935e-08 0.0007 3.97965e-08 0 3.99705e-08 0 3.99735e-08 0.0007 3.99765e-08 0 4.01505e-08 0 4.01535e-08 0.0007 4.01565e-08 0 4.03305e-08 0 4.03335e-08 0.0007 4.03365e-08 0 4.05105e-08 0 4.05135e-08 0.0007 4.05165e-08 0 4.06905e-08 0 4.06935e-08 0.0007 4.06965e-08 0 4.08705e-08 0 4.08735e-08 0.0007 4.08765e-08 0 4.10505e-08 0 4.10535e-08 0.0007 4.10565e-08 0 4.12305e-08 0 4.12335e-08 0.0007 4.12365e-08 0 4.14105e-08 0 4.14135e-08 0.0007 4.14165e-08 0 4.15905e-08 0 4.15935e-08 0.0007 4.15965e-08 0 4.17705e-08 0 4.17735e-08 0.0007 4.17765e-08 0 4.19505e-08 0 4.19535e-08 0.0007 4.19565e-08 0 4.21305e-08 0 4.21335e-08 0.0007 4.21365e-08 0 4.23105e-08 0 4.23135e-08 0.0007 4.23165e-08 0 4.24905e-08 0 4.24935e-08 0.0007 4.24965e-08 0 4.26705e-08 0 4.26735e-08 0.0007 4.26765e-08 0 4.28505e-08 0 4.28535e-08 0.0007 4.28565e-08 0 4.30305e-08 0 4.30335e-08 0.0007 4.30365e-08 0 4.32105e-08 0 4.32135e-08 0.0007 4.32165e-08 0 4.33905e-08 0 4.33935e-08 0.0007 4.33965e-08 0 4.35705e-08 0 4.35735e-08 0.0007 4.35765e-08 0 4.37505e-08 0 4.37535e-08 0.0007 4.37565e-08 0 4.39305e-08 0 4.39335e-08 0.0007 4.39365e-08 0 4.41105e-08 0 4.41135e-08 0.0007 4.41165e-08 0 4.42905e-08 0 4.42935e-08 0.0007 4.42965e-08 0 4.44705e-08 0 4.44735e-08 0.0007 4.44765e-08 0 4.46505e-08 0 4.46535e-08 0.0007 4.46565e-08 0 4.48305e-08 0 4.48335e-08 0.0007 4.48365e-08 0 4.50105e-08 0 4.50135e-08 0.0007 4.50165e-08 0 4.51905e-08 0 4.51935e-08 0.0007 4.51965e-08 0 4.53705e-08 0 4.53735e-08 0.0007 4.53765e-08 0 4.55505e-08 0 4.55535e-08 0.0007 4.55565e-08 0 4.57305e-08 0 4.57335e-08 0.0007 4.57365e-08 0 4.59105e-08 0 4.59135e-08 0.0007 4.59165e-08 0)
B_DFF_IP3_01|1 _DFF_IP3_01|1 _DFF_IP3_01|2 JJMIT AREA=2.5
B_DFF_IP3_01|2 _DFF_IP3_01|4 _DFF_IP3_01|5 JJMIT AREA=1.61
B_DFF_IP3_01|3 _DFF_IP3_01|5 _DFF_IP3_01|6 JJMIT AREA=1.54
B_DFF_IP3_01|4 _DFF_IP3_01|8 _DFF_IP3_01|9 JJMIT AREA=1.69
B_DFF_IP3_01|5 _DFF_IP3_01|10 _DFF_IP3_01|8 JJMIT AREA=1.38
B_DFF_IP3_01|6 _DFF_IP3_01|11 _DFF_IP3_01|12 JJMIT AREA=2.5
B_DFF_IP3_01|7 _DFF_IP3_01|14 _DFF_IP3_01|15 JJMIT AREA=2.5
I_DFF_IP3_01|B1 0 _DFF_IP3_01|3  PWL(0 0 5e-12 0.000175)
I_DFF_IP3_01|B2 0 _DFF_IP3_01|7  PWL(0 0 5e-12 0.000173)
I_DFF_IP3_01|B3 0 _DFF_IP3_01|13  PWL(0 0 5e-12 0.000175)
I_DFF_IP3_01|B4 0 _DFF_IP3_01|16  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|B1 _DFF_IP3_01|3 _DFF_IP3_01|1  2e-12
L_DFF_IP3_01|B2 _DFF_IP3_01|7 _DFF_IP3_01|5  2e-12
L_DFF_IP3_01|B3 _DFF_IP3_01|11 _DFF_IP3_01|13  2e-12
L_DFF_IP3_01|B4 _DFF_IP3_01|16 _DFF_IP3_01|14  2e-12
L_DFF_IP3_01|1 IP3_0_OUT _DFF_IP3_01|1  2.059e-12
L_DFF_IP3_01|2 _DFF_IP3_01|1 _DFF_IP3_01|4  4.123e-12
L_DFF_IP3_01|3 _DFF_IP3_01|5 _DFF_IP3_01|8  6.873e-12
L_DFF_IP3_01|4 _DFF_IP3_01|10 _DFF_IP3_01|11  5.195e-12
L_DFF_IP3_01|5 D03 _DFF_IP3_01|11  2.071e-12
L_DFF_IP3_01|6 _DFF_IP3_01|8 _DFF_IP3_01|14  3.287e-12
L_DFF_IP3_01|7 _DFF_IP3_01|14 IP3_1_OUT  2.066e-12
L_DFF_IP3_01|P1 _DFF_IP3_01|2 0  5.042e-13
L_DFF_IP3_01|P3 _DFF_IP3_01|6 0  5.799e-13
L_DFF_IP3_01|P4 _DFF_IP3_01|9 0  5.733e-13
L_DFF_IP3_01|P6 _DFF_IP3_01|12 0  4.605e-13
L_DFF_IP3_01|P7 _DFF_IP3_01|15 0  4.961e-13
R_DFF_IP3_01|B1 _DFF_IP3_01|1 _DFF_IP3_01|101  2.7439617672
L_DFF_IP3_01|RB1 _DFF_IP3_01|101 0  1.550338398468e-12
R_DFF_IP3_01|B2 _DFF_IP3_01|4 _DFF_IP3_01|104  4.260810197515528
L_DFF_IP3_01|RB2 _DFF_IP3_01|104 _DFF_IP3_01|5  2.407357761596273e-12
R_DFF_IP3_01|B3 _DFF_IP3_01|5 _DFF_IP3_01|105  4.454483388311688
L_DFF_IP3_01|RB3 _DFF_IP3_01|105 0  2.516783114396104e-12
R_DFF_IP3_01|B4 _DFF_IP3_01|8 _DFF_IP3_01|108  4.059115040236686
L_DFF_IP3_01|RB4 _DFF_IP3_01|108 0  2.2933999977337278e-12
R_DFF_IP3_01|B5 _DFF_IP3_01|10 _DFF_IP3_01|110  4.970945230434783
L_DFF_IP3_01|RB5 _DFF_IP3_01|110 _DFF_IP3_01|8  2.8085840551956523e-12
R_DFF_IP3_01|B6 _DFF_IP3_01|11 _DFF_IP3_01|111  2.7439617672
L_DFF_IP3_01|RB6 _DFF_IP3_01|111 0  1.550338398468e-12
R_DFF_IP3_01|B7 _DFF_IP3_01|14 _DFF_IP3_01|114  2.7439617672
L_DFF_IP3_01|RB7 _DFF_IP3_01|114 0  1.550338398468e-12
IT08|T 0 T08  PWL(0 0 6e-12 0 9e-12 0.0014 1.2e-11 0 1.86e-10 0 1.89e-10 0.0014 1.92e-10 0 3.66e-10 0 3.69e-10 0.0014 3.72e-10 0 5.46e-10 0 5.49e-10 0.0014 5.52e-10 0 7.26e-10 0 7.29e-10 0.0014 7.32e-10 0 9.06e-10 0 9.09e-10 0.0014 9.12e-10 0 1.086e-09 0 1.089e-09 0.0014 1.092e-09 0 1.266e-09 0 1.269e-09 0.0014 1.272e-09 0 1.446e-09 0 1.449e-09 0.0014 1.452e-09 0 1.626e-09 0 1.629e-09 0.0014 1.632e-09 0 1.806e-09 0 1.809e-09 0.0014 1.812e-09 0 1.986e-09 0 1.989e-09 0.0014 1.992e-09 0 2.166e-09 0 2.169e-09 0.0014 2.172e-09 0 2.346e-09 0 2.349e-09 0.0014 2.352e-09 0 2.526e-09 0 2.529e-09 0.0014 2.532e-09 0 2.706e-09 0 2.709e-09 0.0014 2.712e-09 0 2.886e-09 0 2.889e-09 0.0014 2.892e-09 0 3.066e-09 0 3.069e-09 0.0014 3.072e-09 0 3.246e-09 0 3.249e-09 0.0014 3.252e-09 0 3.426e-09 0 3.429e-09 0.0014 3.432e-09 0 3.606e-09 0 3.609e-09 0.0014 3.612e-09 0 3.786e-09 0 3.789e-09 0.0014 3.792e-09 0 3.966e-09 0 3.969e-09 0.0014 3.972e-09 0 4.146e-09 0 4.149e-09 0.0014 4.152e-09 0 4.326e-09 0 4.329e-09 0.0014 4.332e-09 0 4.506e-09 0 4.509e-09 0.0014 4.512e-09 0 4.686e-09 0 4.689e-09 0.0014 4.692e-09 0 4.866e-09 0 4.869e-09 0.0014 4.872e-09 0 5.046e-09 0 5.049e-09 0.0014 5.052e-09 0 5.226e-09 0 5.229e-09 0.0014 5.232e-09 0 5.406e-09 0 5.409e-09 0.0014 5.412e-09 0 5.586e-09 0 5.589e-09 0.0014 5.592e-09 0 5.766e-09 0 5.769e-09 0.0014 5.772e-09 0 5.946e-09 0 5.949e-09 0.0014 5.952e-09 0 6.126e-09 0 6.129e-09 0.0014 6.132e-09 0 6.306e-09 0 6.309e-09 0.0014 6.312e-09 0 6.486e-09 0 6.489e-09 0.0014 6.492e-09 0 6.666e-09 0 6.669e-09 0.0014 6.672e-09 0 6.846e-09 0 6.849e-09 0.0014 6.852e-09 0 7.026e-09 0 7.029e-09 0.0014 7.032e-09 0 7.206e-09 0 7.209e-09 0.0014 7.212e-09 0 7.386e-09 0 7.389e-09 0.0014 7.392e-09 0 7.566e-09 0 7.569e-09 0.0014 7.572e-09 0 7.746e-09 0 7.749e-09 0.0014 7.752e-09 0 7.926e-09 0 7.929e-09 0.0014 7.932e-09 0 8.106e-09 0 8.109e-09 0.0014 8.112e-09 0 8.286e-09 0 8.289e-09 0.0014 8.292e-09 0 8.466e-09 0 8.469e-09 0.0014 8.472e-09 0 8.646e-09 0 8.649e-09 0.0014 8.652e-09 0 8.826e-09 0 8.829e-09 0.0014 8.832e-09 0 9.006e-09 0 9.009e-09 0.0014 9.012e-09 0 9.186e-09 0 9.189e-09 0.0014 9.192e-09 0 9.366e-09 0 9.369e-09 0.0014 9.372e-09 0 9.546e-09 0 9.549e-09 0.0014 9.552e-09 0 9.726e-09 0 9.729e-09 0.0014 9.732e-09 0 9.906e-09 0 9.909e-09 0.0014 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0014 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0014 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0014 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0014 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0014 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0014 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0014 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0014 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0014 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0014 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0014 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0014 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0014 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0014 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0014 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0014 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0014 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0014 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0014 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0014 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0014 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0014 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0014 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0014 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0014 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0014 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0014 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0014 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0014 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0014 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0014 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0014 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0014 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0014 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0014 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0014 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0014 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0014 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0014 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0014 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0014 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0014 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0014 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0014 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0014 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0014 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0014 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0014 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0014 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0014 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0014 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0014 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0014 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0014 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0014 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0014 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0014 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0014 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0014 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0014 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0014 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0014 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0014 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0014 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0014 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0014 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0014 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0014 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0014 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0014 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0014 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0014 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0014 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0014 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0014 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0014 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0014 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0014 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0014 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0014 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0014 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0014 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0014 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0014 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0014 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0014 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0014 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0014 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0014 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0014 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0014 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0014 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0014 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0014 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0014 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0014 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0014 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0014 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0014 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0014 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0014 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0014 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0014 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0014 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0014 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0014 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0014 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0014 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0014 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0014 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0014 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0014 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0014 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0014 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0014 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0014 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0014 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0014 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0014 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0014 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0014 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0014 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0014 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0014 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0014 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0014 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0014 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0014 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0014 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0014 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0014 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0014 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0014 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0014 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0014 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0014 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0014 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0014 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0014 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0014 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0014 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0014 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0014 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0014 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0014 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0014 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0014 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0014 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0014 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0014 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0014 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0014 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0014 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0014 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0014 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0014 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0014 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0014 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0014 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0014 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0014 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0014 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0014 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0014 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0014 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0014 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0014 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0014 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0014 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0014 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0014 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0014 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0014 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0014 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0014 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0014 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0014 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0014 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0014 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0014 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0014 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0014 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0014 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0014 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0014 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0014 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0014 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0014 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0014 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0014 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0014 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0014 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0014 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0014 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0014 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0014 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0014 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0014 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0014 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0014 4.5912e-08 0)
IT09|T 0 T09  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0007 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0007 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0007 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0007 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0007 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0007 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0007 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0007 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0007 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0007 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0007 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0007 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0007 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0007 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0007 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0007 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0007 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0007 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0007 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0007 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0007 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0007 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0007 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0007 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0007 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0007 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0007 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0007 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0007 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0007 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0007 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0007 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0007 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0007 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0007 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0007 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0007 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0007 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0007 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0007 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0007 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0007 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0007 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0007 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0007 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0007 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0007 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0007 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0007 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0007 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0007 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0007 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0007 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0007 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0007 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0007 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0007 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0007 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0007 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0007 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0007 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0007 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0007 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0007 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0007 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0007 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0007 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0007 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0007 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0007 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0007 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0007 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0007 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0007 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0007 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0007 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0007 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0007 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0007 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0007 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0007 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0007 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0007 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0007 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0007 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0007 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0007 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0007 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0007 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0007 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0007 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0007 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0007 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0007 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0007 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0007 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0007 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0007 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0007 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0007 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0007 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0007 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0007 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0007 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0007 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0007 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0007 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0007 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0007 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0007 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0007 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0007 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0007 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0007 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0007 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0007 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0007 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0007 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0007 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0007 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0007 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0007 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0007 4.5912e-08 0)
B_PG1_12|1 _PG1_12|1 _PG1_12|2 JJMIT AREA=2.5
B_PG1_12|2 _PG1_12|4 _PG1_12|5 JJMIT AREA=1.61
B_PG1_12|3 _PG1_12|5 _PG1_12|6 JJMIT AREA=1.54
B_PG1_12|4 _PG1_12|8 _PG1_12|9 JJMIT AREA=1.69
B_PG1_12|5 _PG1_12|10 _PG1_12|8 JJMIT AREA=1.38
B_PG1_12|6 _PG1_12|11 _PG1_12|12 JJMIT AREA=2.5
B_PG1_12|7 _PG1_12|14 _PG1_12|15 JJMIT AREA=2.5
I_PG1_12|B1 0 _PG1_12|3  PWL(0 0 5e-12 0.000175)
I_PG1_12|B2 0 _PG1_12|7  PWL(0 0 5e-12 0.000173)
I_PG1_12|B3 0 _PG1_12|13  PWL(0 0 5e-12 0.000175)
I_PG1_12|B4 0 _PG1_12|16  PWL(0 0 5e-12 0.000175)
L_PG1_12|B1 _PG1_12|3 _PG1_12|1  2e-12
L_PG1_12|B2 _PG1_12|7 _PG1_12|5  2e-12
L_PG1_12|B3 _PG1_12|11 _PG1_12|13  2e-12
L_PG1_12|B4 _PG1_12|16 _PG1_12|14  2e-12
L_PG1_12|1 G1_1_TO1 _PG1_12|1  2.059e-12
L_PG1_12|2 _PG1_12|1 _PG1_12|4  4.123e-12
L_PG1_12|3 _PG1_12|5 _PG1_12|8  6.873e-12
L_PG1_12|4 _PG1_12|10 _PG1_12|11  5.195e-12
L_PG1_12|5 T09 _PG1_12|11  2.071e-12
L_PG1_12|6 _PG1_12|8 _PG1_12|14  3.287e-12
L_PG1_12|7 _PG1_12|14 G1_2  2.066e-12
L_PG1_12|P1 _PG1_12|2 0  5.042e-13
L_PG1_12|P3 _PG1_12|6 0  5.799e-13
L_PG1_12|P4 _PG1_12|9 0  5.733e-13
L_PG1_12|P6 _PG1_12|12 0  4.605e-13
L_PG1_12|P7 _PG1_12|15 0  4.961e-13
R_PG1_12|B1 _PG1_12|1 _PG1_12|101  2.7439617672
L_PG1_12|RB1 _PG1_12|101 0  1.550338398468e-12
R_PG1_12|B2 _PG1_12|4 _PG1_12|104  4.260810197515528
L_PG1_12|RB2 _PG1_12|104 _PG1_12|5  2.407357761596273e-12
R_PG1_12|B3 _PG1_12|5 _PG1_12|105  4.454483388311688
L_PG1_12|RB3 _PG1_12|105 0  2.516783114396104e-12
R_PG1_12|B4 _PG1_12|8 _PG1_12|108  4.059115040236686
L_PG1_12|RB4 _PG1_12|108 0  2.2933999977337278e-12
R_PG1_12|B5 _PG1_12|10 _PG1_12|110  4.970945230434783
L_PG1_12|RB5 _PG1_12|110 _PG1_12|8  2.8085840551956523e-12
R_PG1_12|B6 _PG1_12|11 _PG1_12|111  2.7439617672
L_PG1_12|RB6 _PG1_12|111 0  1.550338398468e-12
R_PG1_12|B7 _PG1_12|14 _PG1_12|114  2.7439617672
L_PG1_12|RB7 _PG1_12|114 0  1.550338398468e-12
IT10|T 0 T10  PWL(0 0 6e-12 0 9e-12 0.0014 1.2e-11 0 1.86e-10 0 1.89e-10 0.0014 1.92e-10 0 3.66e-10 0 3.69e-10 0.0014 3.72e-10 0 5.46e-10 0 5.49e-10 0.0014 5.52e-10 0 7.26e-10 0 7.29e-10 0.0014 7.32e-10 0 9.06e-10 0 9.09e-10 0.0014 9.12e-10 0 1.086e-09 0 1.089e-09 0.0014 1.092e-09 0 1.266e-09 0 1.269e-09 0.0014 1.272e-09 0 1.446e-09 0 1.449e-09 0.0014 1.452e-09 0 1.626e-09 0 1.629e-09 0.0014 1.632e-09 0 1.806e-09 0 1.809e-09 0.0014 1.812e-09 0 1.986e-09 0 1.989e-09 0.0014 1.992e-09 0 2.166e-09 0 2.169e-09 0.0014 2.172e-09 0 2.346e-09 0 2.349e-09 0.0014 2.352e-09 0 2.526e-09 0 2.529e-09 0.0014 2.532e-09 0 2.706e-09 0 2.709e-09 0.0014 2.712e-09 0 2.886e-09 0 2.889e-09 0.0014 2.892e-09 0 3.066e-09 0 3.069e-09 0.0014 3.072e-09 0 3.246e-09 0 3.249e-09 0.0014 3.252e-09 0 3.426e-09 0 3.429e-09 0.0014 3.432e-09 0 3.606e-09 0 3.609e-09 0.0014 3.612e-09 0 3.786e-09 0 3.789e-09 0.0014 3.792e-09 0 3.966e-09 0 3.969e-09 0.0014 3.972e-09 0 4.146e-09 0 4.149e-09 0.0014 4.152e-09 0 4.326e-09 0 4.329e-09 0.0014 4.332e-09 0 4.506e-09 0 4.509e-09 0.0014 4.512e-09 0 4.686e-09 0 4.689e-09 0.0014 4.692e-09 0 4.866e-09 0 4.869e-09 0.0014 4.872e-09 0 5.046e-09 0 5.049e-09 0.0014 5.052e-09 0 5.226e-09 0 5.229e-09 0.0014 5.232e-09 0 5.406e-09 0 5.409e-09 0.0014 5.412e-09 0 5.586e-09 0 5.589e-09 0.0014 5.592e-09 0 5.766e-09 0 5.769e-09 0.0014 5.772e-09 0 5.946e-09 0 5.949e-09 0.0014 5.952e-09 0 6.126e-09 0 6.129e-09 0.0014 6.132e-09 0 6.306e-09 0 6.309e-09 0.0014 6.312e-09 0 6.486e-09 0 6.489e-09 0.0014 6.492e-09 0 6.666e-09 0 6.669e-09 0.0014 6.672e-09 0 6.846e-09 0 6.849e-09 0.0014 6.852e-09 0 7.026e-09 0 7.029e-09 0.0014 7.032e-09 0 7.206e-09 0 7.209e-09 0.0014 7.212e-09 0 7.386e-09 0 7.389e-09 0.0014 7.392e-09 0 7.566e-09 0 7.569e-09 0.0014 7.572e-09 0 7.746e-09 0 7.749e-09 0.0014 7.752e-09 0 7.926e-09 0 7.929e-09 0.0014 7.932e-09 0 8.106e-09 0 8.109e-09 0.0014 8.112e-09 0 8.286e-09 0 8.289e-09 0.0014 8.292e-09 0 8.466e-09 0 8.469e-09 0.0014 8.472e-09 0 8.646e-09 0 8.649e-09 0.0014 8.652e-09 0 8.826e-09 0 8.829e-09 0.0014 8.832e-09 0 9.006e-09 0 9.009e-09 0.0014 9.012e-09 0 9.186e-09 0 9.189e-09 0.0014 9.192e-09 0 9.366e-09 0 9.369e-09 0.0014 9.372e-09 0 9.546e-09 0 9.549e-09 0.0014 9.552e-09 0 9.726e-09 0 9.729e-09 0.0014 9.732e-09 0 9.906e-09 0 9.909e-09 0.0014 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0014 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0014 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0014 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0014 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0014 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0014 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0014 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0014 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0014 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0014 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0014 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0014 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0014 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0014 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0014 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0014 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0014 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0014 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0014 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0014 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0014 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0014 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0014 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0014 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0014 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0014 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0014 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0014 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0014 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0014 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0014 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0014 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0014 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0014 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0014 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0014 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0014 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0014 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0014 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0014 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0014 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0014 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0014 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0014 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0014 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0014 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0014 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0014 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0014 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0014 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0014 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0014 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0014 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0014 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0014 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0014 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0014 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0014 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0014 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0014 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0014 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0014 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0014 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0014 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0014 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0014 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0014 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0014 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0014 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0014 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0014 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0014 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0014 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0014 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0014 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0014 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0014 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0014 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0014 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0014 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0014 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0014 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0014 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0014 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0014 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0014 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0014 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0014 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0014 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0014 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0014 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0014 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0014 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0014 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0014 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0014 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0014 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0014 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0014 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0014 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0014 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0014 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0014 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0014 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0014 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0014 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0014 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0014 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0014 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0014 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0014 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0014 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0014 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0014 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0014 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0014 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0014 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0014 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0014 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0014 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0014 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0014 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0014 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0014 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0014 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0014 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0014 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0014 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0014 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0014 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0014 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0014 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0014 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0014 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0014 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0014 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0014 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0014 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0014 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0014 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0014 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0014 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0014 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0014 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0014 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0014 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0014 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0014 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0014 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0014 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0014 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0014 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0014 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0014 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0014 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0014 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0014 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0014 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0014 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0014 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0014 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0014 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0014 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0014 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0014 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0014 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0014 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0014 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0014 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0014 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0014 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0014 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0014 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0014 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0014 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0014 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0014 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0014 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0014 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0014 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0014 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0014 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0014 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0014 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0014 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0014 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0014 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0014 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0014 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0014 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0014 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0014 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0014 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0014 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0014 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0014 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0014 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0014 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0014 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0014 4.5912e-08 0)
IT11|T 0 T11  PWL(0 0 6e-12 0 9e-12 0.0014 1.2e-11 0 1.86e-10 0 1.89e-10 0.0014 1.92e-10 0 3.66e-10 0 3.69e-10 0.0014 3.72e-10 0 5.46e-10 0 5.49e-10 0.0014 5.52e-10 0 7.26e-10 0 7.29e-10 0.0014 7.32e-10 0 9.06e-10 0 9.09e-10 0.0014 9.12e-10 0 1.086e-09 0 1.089e-09 0.0014 1.092e-09 0 1.266e-09 0 1.269e-09 0.0014 1.272e-09 0 1.446e-09 0 1.449e-09 0.0014 1.452e-09 0 1.626e-09 0 1.629e-09 0.0014 1.632e-09 0 1.806e-09 0 1.809e-09 0.0014 1.812e-09 0 1.986e-09 0 1.989e-09 0.0014 1.992e-09 0 2.166e-09 0 2.169e-09 0.0014 2.172e-09 0 2.346e-09 0 2.349e-09 0.0014 2.352e-09 0 2.526e-09 0 2.529e-09 0.0014 2.532e-09 0 2.706e-09 0 2.709e-09 0.0014 2.712e-09 0 2.886e-09 0 2.889e-09 0.0014 2.892e-09 0 3.066e-09 0 3.069e-09 0.0014 3.072e-09 0 3.246e-09 0 3.249e-09 0.0014 3.252e-09 0 3.426e-09 0 3.429e-09 0.0014 3.432e-09 0 3.606e-09 0 3.609e-09 0.0014 3.612e-09 0 3.786e-09 0 3.789e-09 0.0014 3.792e-09 0 3.966e-09 0 3.969e-09 0.0014 3.972e-09 0 4.146e-09 0 4.149e-09 0.0014 4.152e-09 0 4.326e-09 0 4.329e-09 0.0014 4.332e-09 0 4.506e-09 0 4.509e-09 0.0014 4.512e-09 0 4.686e-09 0 4.689e-09 0.0014 4.692e-09 0 4.866e-09 0 4.869e-09 0.0014 4.872e-09 0 5.046e-09 0 5.049e-09 0.0014 5.052e-09 0 5.226e-09 0 5.229e-09 0.0014 5.232e-09 0 5.406e-09 0 5.409e-09 0.0014 5.412e-09 0 5.586e-09 0 5.589e-09 0.0014 5.592e-09 0 5.766e-09 0 5.769e-09 0.0014 5.772e-09 0 5.946e-09 0 5.949e-09 0.0014 5.952e-09 0 6.126e-09 0 6.129e-09 0.0014 6.132e-09 0 6.306e-09 0 6.309e-09 0.0014 6.312e-09 0 6.486e-09 0 6.489e-09 0.0014 6.492e-09 0 6.666e-09 0 6.669e-09 0.0014 6.672e-09 0 6.846e-09 0 6.849e-09 0.0014 6.852e-09 0 7.026e-09 0 7.029e-09 0.0014 7.032e-09 0 7.206e-09 0 7.209e-09 0.0014 7.212e-09 0 7.386e-09 0 7.389e-09 0.0014 7.392e-09 0 7.566e-09 0 7.569e-09 0.0014 7.572e-09 0 7.746e-09 0 7.749e-09 0.0014 7.752e-09 0 7.926e-09 0 7.929e-09 0.0014 7.932e-09 0 8.106e-09 0 8.109e-09 0.0014 8.112e-09 0 8.286e-09 0 8.289e-09 0.0014 8.292e-09 0 8.466e-09 0 8.469e-09 0.0014 8.472e-09 0 8.646e-09 0 8.649e-09 0.0014 8.652e-09 0 8.826e-09 0 8.829e-09 0.0014 8.832e-09 0 9.006e-09 0 9.009e-09 0.0014 9.012e-09 0 9.186e-09 0 9.189e-09 0.0014 9.192e-09 0 9.366e-09 0 9.369e-09 0.0014 9.372e-09 0 9.546e-09 0 9.549e-09 0.0014 9.552e-09 0 9.726e-09 0 9.729e-09 0.0014 9.732e-09 0 9.906e-09 0 9.909e-09 0.0014 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0014 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0014 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0014 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0014 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0014 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0014 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0014 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0014 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0014 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0014 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0014 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0014 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0014 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0014 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0014 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0014 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0014 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0014 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0014 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0014 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0014 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0014 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0014 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0014 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0014 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0014 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0014 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0014 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0014 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0014 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0014 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0014 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0014 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0014 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0014 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0014 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0014 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0014 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0014 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0014 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0014 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0014 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0014 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0014 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0014 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0014 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0014 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0014 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0014 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0014 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0014 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0014 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0014 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0014 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0014 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0014 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0014 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0014 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0014 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0014 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0014 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0014 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0014 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0014 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0014 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0014 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0014 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0014 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0014 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0014 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0014 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0014 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0014 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0014 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0014 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0014 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0014 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0014 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0014 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0014 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0014 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0014 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0014 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0014 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0014 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0014 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0014 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0014 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0014 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0014 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0014 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0014 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0014 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0014 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0014 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0014 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0014 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0014 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0014 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0014 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0014 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0014 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0014 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0014 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0014 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0014 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0014 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0014 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0014 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0014 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0014 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0014 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0014 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0014 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0014 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0014 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0014 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0014 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0014 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0014 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0014 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0014 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0014 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0014 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0014 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0014 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0014 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0014 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0014 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0014 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0014 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0014 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0014 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0014 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0014 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0014 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0014 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0014 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0014 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0014 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0014 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0014 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0014 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0014 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0014 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0014 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0014 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0014 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0014 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0014 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0014 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0014 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0014 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0014 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0014 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0014 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0014 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0014 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0014 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0014 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0014 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0014 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0014 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0014 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0014 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0014 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0014 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0014 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0014 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0014 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0014 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0014 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0014 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0014 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0014 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0014 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0014 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0014 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0014 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0014 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0014 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0014 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0014 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0014 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0014 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0014 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0014 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0014 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0014 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0014 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0014 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0014 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0014 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0014 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0014 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0014 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0014 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0014 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0014 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0014 4.5912e-08 0)
ID11|T 0 D11  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0007 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0007 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0007 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0007 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0007 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0007 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0007 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0007 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0007 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0007 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0007 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0007 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0007 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0007 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0007 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0007 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0007 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0007 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0007 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0007 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0007 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0007 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0007 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0007 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0007 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0007 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0007 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0007 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0007 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0007 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0007 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0007 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0007 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0007 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0007 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0007 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0007 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0007 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0007 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0007 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0007 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0007 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0007 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0007 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0007 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0007 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0007 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0007 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0007 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0007 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0007 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0007 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0007 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0007 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0007 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0007 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0007 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0007 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0007 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0007 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0007 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0007 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0007 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0007 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0007 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0007 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0007 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0007 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0007 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0007 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0007 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0007 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0007 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0007 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0007 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0007 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0007 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0007 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0007 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0007 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0007 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0007 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0007 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0007 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0007 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0007 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0007 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0007 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0007 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0007 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0007 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0007 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0007 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0007 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0007 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0007 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0007 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0007 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0007 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0007 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0007 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0007 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0007 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0007 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0007 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0007 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0007 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0007 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0007 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0007 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0007 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0007 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0007 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0007 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0007 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0007 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0007 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0007 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0007 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0007 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0007 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0007 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0007 4.5912e-08 0)
B_DFF_IP1_12|1 _DFF_IP1_12|1 _DFF_IP1_12|2 JJMIT AREA=2.5
B_DFF_IP1_12|2 _DFF_IP1_12|4 _DFF_IP1_12|5 JJMIT AREA=1.61
B_DFF_IP1_12|3 _DFF_IP1_12|5 _DFF_IP1_12|6 JJMIT AREA=1.54
B_DFF_IP1_12|4 _DFF_IP1_12|8 _DFF_IP1_12|9 JJMIT AREA=1.69
B_DFF_IP1_12|5 _DFF_IP1_12|10 _DFF_IP1_12|8 JJMIT AREA=1.38
B_DFF_IP1_12|6 _DFF_IP1_12|11 _DFF_IP1_12|12 JJMIT AREA=2.5
B_DFF_IP1_12|7 _DFF_IP1_12|14 _DFF_IP1_12|15 JJMIT AREA=2.5
I_DFF_IP1_12|B1 0 _DFF_IP1_12|3  PWL(0 0 5e-12 0.000175)
I_DFF_IP1_12|B2 0 _DFF_IP1_12|7  PWL(0 0 5e-12 0.000173)
I_DFF_IP1_12|B3 0 _DFF_IP1_12|13  PWL(0 0 5e-12 0.000175)
I_DFF_IP1_12|B4 0 _DFF_IP1_12|16  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|B1 _DFF_IP1_12|3 _DFF_IP1_12|1  2e-12
L_DFF_IP1_12|B2 _DFF_IP1_12|7 _DFF_IP1_12|5  2e-12
L_DFF_IP1_12|B3 _DFF_IP1_12|11 _DFF_IP1_12|13  2e-12
L_DFF_IP1_12|B4 _DFF_IP1_12|16 _DFF_IP1_12|14  2e-12
L_DFF_IP1_12|1 IP1_1_OUT_RX _DFF_IP1_12|1  2.059e-12
L_DFF_IP1_12|2 _DFF_IP1_12|1 _DFF_IP1_12|4  4.123e-12
L_DFF_IP1_12|3 _DFF_IP1_12|5 _DFF_IP1_12|8  6.873e-12
L_DFF_IP1_12|4 _DFF_IP1_12|10 _DFF_IP1_12|11  5.195e-12
L_DFF_IP1_12|5 D11 _DFF_IP1_12|11  2.071e-12
L_DFF_IP1_12|6 _DFF_IP1_12|8 _DFF_IP1_12|14  3.287e-12
L_DFF_IP1_12|7 _DFF_IP1_12|14 IP1_2_OUT  2.066e-12
L_DFF_IP1_12|P1 _DFF_IP1_12|2 0  5.042e-13
L_DFF_IP1_12|P3 _DFF_IP1_12|6 0  5.799e-13
L_DFF_IP1_12|P4 _DFF_IP1_12|9 0  5.733e-13
L_DFF_IP1_12|P6 _DFF_IP1_12|12 0  4.605e-13
L_DFF_IP1_12|P7 _DFF_IP1_12|15 0  4.961e-13
R_DFF_IP1_12|B1 _DFF_IP1_12|1 _DFF_IP1_12|101  2.7439617672
L_DFF_IP1_12|RB1 _DFF_IP1_12|101 0  1.550338398468e-12
R_DFF_IP1_12|B2 _DFF_IP1_12|4 _DFF_IP1_12|104  4.260810197515528
L_DFF_IP1_12|RB2 _DFF_IP1_12|104 _DFF_IP1_12|5  2.407357761596273e-12
R_DFF_IP1_12|B3 _DFF_IP1_12|5 _DFF_IP1_12|105  4.454483388311688
L_DFF_IP1_12|RB3 _DFF_IP1_12|105 0  2.516783114396104e-12
R_DFF_IP1_12|B4 _DFF_IP1_12|8 _DFF_IP1_12|108  4.059115040236686
L_DFF_IP1_12|RB4 _DFF_IP1_12|108 0  2.2933999977337278e-12
R_DFF_IP1_12|B5 _DFF_IP1_12|10 _DFF_IP1_12|110  4.970945230434783
L_DFF_IP1_12|RB5 _DFF_IP1_12|110 _DFF_IP1_12|8  2.8085840551956523e-12
R_DFF_IP1_12|B6 _DFF_IP1_12|11 _DFF_IP1_12|111  2.7439617672
L_DFF_IP1_12|RB6 _DFF_IP1_12|111 0  1.550338398468e-12
R_DFF_IP1_12|B7 _DFF_IP1_12|14 _DFF_IP1_12|114  2.7439617672
L_DFF_IP1_12|RB7 _DFF_IP1_12|114 0  1.550338398468e-12
ID12|T 0 D12  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0007 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0007 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0007 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0007 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0007 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0007 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0007 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0007 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0007 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0007 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0007 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0007 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0007 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0007 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0007 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0007 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0007 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0007 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0007 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0007 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0007 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0007 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0007 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0007 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0007 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0007 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0007 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0007 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0007 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0007 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0007 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0007 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0007 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0007 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0007 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0007 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0007 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0007 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0007 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0007 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0007 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0007 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0007 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0007 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0007 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0007 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0007 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0007 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0007 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0007 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0007 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0007 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0007 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0007 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0007 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0007 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0007 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0007 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0007 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0007 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0007 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0007 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0007 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0007 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0007 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0007 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0007 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0007 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0007 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0007 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0007 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0007 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0007 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0007 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0007 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0007 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0007 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0007 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0007 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0007 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0007 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0007 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0007 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0007 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0007 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0007 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0007 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0007 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0007 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0007 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0007 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0007 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0007 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0007 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0007 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0007 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0007 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0007 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0007 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0007 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0007 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0007 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0007 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0007 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0007 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0007 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0007 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0007 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0007 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0007 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0007 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0007 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0007 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0007 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0007 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0007 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0007 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0007 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0007 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0007 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0007 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0007 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0007 4.5912e-08 0)
B_DFF_IP2_12|1 _DFF_IP2_12|1 _DFF_IP2_12|2 JJMIT AREA=2.5
B_DFF_IP2_12|2 _DFF_IP2_12|4 _DFF_IP2_12|5 JJMIT AREA=1.61
B_DFF_IP2_12|3 _DFF_IP2_12|5 _DFF_IP2_12|6 JJMIT AREA=1.54
B_DFF_IP2_12|4 _DFF_IP2_12|8 _DFF_IP2_12|9 JJMIT AREA=1.69
B_DFF_IP2_12|5 _DFF_IP2_12|10 _DFF_IP2_12|8 JJMIT AREA=1.38
B_DFF_IP2_12|6 _DFF_IP2_12|11 _DFF_IP2_12|12 JJMIT AREA=2.5
B_DFF_IP2_12|7 _DFF_IP2_12|14 _DFF_IP2_12|15 JJMIT AREA=2.5
I_DFF_IP2_12|B1 0 _DFF_IP2_12|3  PWL(0 0 5e-12 0.000175)
I_DFF_IP2_12|B2 0 _DFF_IP2_12|7  PWL(0 0 5e-12 0.000173)
I_DFF_IP2_12|B3 0 _DFF_IP2_12|13  PWL(0 0 5e-12 0.000175)
I_DFF_IP2_12|B4 0 _DFF_IP2_12|16  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|B1 _DFF_IP2_12|3 _DFF_IP2_12|1  2e-12
L_DFF_IP2_12|B2 _DFF_IP2_12|7 _DFF_IP2_12|5  2e-12
L_DFF_IP2_12|B3 _DFF_IP2_12|11 _DFF_IP2_12|13  2e-12
L_DFF_IP2_12|B4 _DFF_IP2_12|16 _DFF_IP2_12|14  2e-12
L_DFF_IP2_12|1 IP2_1_OUT_RX _DFF_IP2_12|1  2.059e-12
L_DFF_IP2_12|2 _DFF_IP2_12|1 _DFF_IP2_12|4  4.123e-12
L_DFF_IP2_12|3 _DFF_IP2_12|5 _DFF_IP2_12|8  6.873e-12
L_DFF_IP2_12|4 _DFF_IP2_12|10 _DFF_IP2_12|11  5.195e-12
L_DFF_IP2_12|5 D12 _DFF_IP2_12|11  2.071e-12
L_DFF_IP2_12|6 _DFF_IP2_12|8 _DFF_IP2_12|14  3.287e-12
L_DFF_IP2_12|7 _DFF_IP2_12|14 IP2_2_OUT  2.066e-12
L_DFF_IP2_12|P1 _DFF_IP2_12|2 0  5.042e-13
L_DFF_IP2_12|P3 _DFF_IP2_12|6 0  5.799e-13
L_DFF_IP2_12|P4 _DFF_IP2_12|9 0  5.733e-13
L_DFF_IP2_12|P6 _DFF_IP2_12|12 0  4.605e-13
L_DFF_IP2_12|P7 _DFF_IP2_12|15 0  4.961e-13
R_DFF_IP2_12|B1 _DFF_IP2_12|1 _DFF_IP2_12|101  2.7439617672
L_DFF_IP2_12|RB1 _DFF_IP2_12|101 0  1.550338398468e-12
R_DFF_IP2_12|B2 _DFF_IP2_12|4 _DFF_IP2_12|104  4.260810197515528
L_DFF_IP2_12|RB2 _DFF_IP2_12|104 _DFF_IP2_12|5  2.407357761596273e-12
R_DFF_IP2_12|B3 _DFF_IP2_12|5 _DFF_IP2_12|105  4.454483388311688
L_DFF_IP2_12|RB3 _DFF_IP2_12|105 0  2.516783114396104e-12
R_DFF_IP2_12|B4 _DFF_IP2_12|8 _DFF_IP2_12|108  4.059115040236686
L_DFF_IP2_12|RB4 _DFF_IP2_12|108 0  2.2933999977337278e-12
R_DFF_IP2_12|B5 _DFF_IP2_12|10 _DFF_IP2_12|110  4.970945230434783
L_DFF_IP2_12|RB5 _DFF_IP2_12|110 _DFF_IP2_12|8  2.8085840551956523e-12
R_DFF_IP2_12|B6 _DFF_IP2_12|11 _DFF_IP2_12|111  2.7439617672
L_DFF_IP2_12|RB6 _DFF_IP2_12|111 0  1.550338398468e-12
R_DFF_IP2_12|B7 _DFF_IP2_12|14 _DFF_IP2_12|114  2.7439617672
L_DFF_IP2_12|RB7 _DFF_IP2_12|114 0  1.550338398468e-12
ID13|T 0 D13  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3946e-08 0 2.3949e-08 0.0007 2.3952e-08 0 2.4126e-08 0 2.4129e-08 0.0007 2.4132e-08 0 2.4306e-08 0 2.4309e-08 0.0007 2.4312e-08 0 2.4486e-08 0 2.4489e-08 0.0007 2.4492e-08 0 2.4666e-08 0 2.4669e-08 0.0007 2.4672e-08 0 2.4846e-08 0 2.4849e-08 0.0007 2.4852e-08 0 2.5026e-08 0 2.5029e-08 0.0007 2.5032e-08 0 2.5206e-08 0 2.5209e-08 0.0007 2.5212e-08 0 2.5386e-08 0 2.5389e-08 0.0007 2.5392e-08 0 2.5566e-08 0 2.5569e-08 0.0007 2.5572e-08 0 2.5746e-08 0 2.5749e-08 0.0007 2.5752e-08 0 2.5926e-08 0 2.5929e-08 0.0007 2.5932e-08 0 2.6106e-08 0 2.6109e-08 0.0007 2.6112e-08 0 2.6286e-08 0 2.6289e-08 0.0007 2.6292e-08 0 2.6466e-08 0 2.6469e-08 0.0007 2.6472e-08 0 2.6646e-08 0 2.6649e-08 0.0007 2.6652e-08 0 2.6826e-08 0 2.6829e-08 0.0007 2.6832e-08 0 2.7006e-08 0 2.7009e-08 0.0007 2.7012e-08 0 2.7186e-08 0 2.7189e-08 0.0007 2.7192e-08 0 2.7366e-08 0 2.7369e-08 0.0007 2.7372e-08 0 2.7546e-08 0 2.7549e-08 0.0007 2.7552e-08 0 2.7726e-08 0 2.7729e-08 0.0007 2.7732e-08 0 2.7906e-08 0 2.7909e-08 0.0007 2.7912e-08 0 2.8086e-08 0 2.8089e-08 0.0007 2.8092e-08 0 2.8266e-08 0 2.8269e-08 0.0007 2.8272e-08 0 2.8446e-08 0 2.8449e-08 0.0007 2.8452e-08 0 2.8626e-08 0 2.8629e-08 0.0007 2.8632e-08 0 2.8806e-08 0 2.8809e-08 0.0007 2.8812e-08 0 2.8986e-08 0 2.8989e-08 0.0007 2.8992e-08 0 2.9166e-08 0 2.9169e-08 0.0007 2.9172e-08 0 2.9346e-08 0 2.9349e-08 0.0007 2.9352e-08 0 2.9526e-08 0 2.9529e-08 0.0007 2.9532e-08 0 2.9706e-08 0 2.9709e-08 0.0007 2.9712e-08 0 2.9886e-08 0 2.9889e-08 0.0007 2.9892e-08 0 3.0066e-08 0 3.0069e-08 0.0007 3.0072e-08 0 3.0246e-08 0 3.0249e-08 0.0007 3.0252e-08 0 3.0426e-08 0 3.0429e-08 0.0007 3.0432e-08 0 3.0606e-08 0 3.0609e-08 0.0007 3.0612e-08 0 3.0786e-08 0 3.0789e-08 0.0007 3.0792e-08 0 3.0966e-08 0 3.0969e-08 0.0007 3.0972e-08 0 3.1146e-08 0 3.1149e-08 0.0007 3.1152e-08 0 3.1326e-08 0 3.1329e-08 0.0007 3.1332e-08 0 3.1506e-08 0 3.1509e-08 0.0007 3.1512e-08 0 3.1686e-08 0 3.1689e-08 0.0007 3.1692e-08 0 3.1866e-08 0 3.1869e-08 0.0007 3.1872e-08 0 3.2046e-08 0 3.2049e-08 0.0007 3.2052e-08 0 3.2226e-08 0 3.2229e-08 0.0007 3.2232e-08 0 3.2406e-08 0 3.2409e-08 0.0007 3.2412e-08 0 3.2586e-08 0 3.2589e-08 0.0007 3.2592e-08 0 3.2766e-08 0 3.2769e-08 0.0007 3.2772e-08 0 3.2946e-08 0 3.2949e-08 0.0007 3.2952e-08 0 3.3126e-08 0 3.3129e-08 0.0007 3.3132e-08 0 3.3306e-08 0 3.3309e-08 0.0007 3.3312e-08 0 3.3486e-08 0 3.3489e-08 0.0007 3.3492e-08 0 3.3666e-08 0 3.3669e-08 0.0007 3.3672e-08 0 3.3846e-08 0 3.3849e-08 0.0007 3.3852e-08 0 3.4026e-08 0 3.4029e-08 0.0007 3.4032e-08 0 3.4206e-08 0 3.4209e-08 0.0007 3.4212e-08 0 3.4386e-08 0 3.4389e-08 0.0007 3.4392e-08 0 3.4566e-08 0 3.4569e-08 0.0007 3.4572e-08 0 3.4746e-08 0 3.4749e-08 0.0007 3.4752e-08 0 3.4926e-08 0 3.4929e-08 0.0007 3.4932e-08 0 3.5106e-08 0 3.5109e-08 0.0007 3.5112e-08 0 3.5286e-08 0 3.5289e-08 0.0007 3.5292e-08 0 3.5466e-08 0 3.5469e-08 0.0007 3.5472e-08 0 3.5646e-08 0 3.5649e-08 0.0007 3.5652e-08 0 3.5826e-08 0 3.5829e-08 0.0007 3.5832e-08 0 3.6006e-08 0 3.6009e-08 0.0007 3.6012e-08 0 3.6186e-08 0 3.6189e-08 0.0007 3.6192e-08 0 3.6366e-08 0 3.6369e-08 0.0007 3.6372e-08 0 3.6546e-08 0 3.6549e-08 0.0007 3.6552e-08 0 3.6726e-08 0 3.6729e-08 0.0007 3.6732e-08 0 3.6906e-08 0 3.6909e-08 0.0007 3.6912e-08 0 3.7086e-08 0 3.7089e-08 0.0007 3.7092e-08 0 3.7266e-08 0 3.7269e-08 0.0007 3.7272e-08 0 3.7446e-08 0 3.7449e-08 0.0007 3.7452e-08 0 3.7626e-08 0 3.7629e-08 0.0007 3.7632e-08 0 3.7806e-08 0 3.7809e-08 0.0007 3.7812e-08 0 3.7986e-08 0 3.7989e-08 0.0007 3.7992e-08 0 3.8166e-08 0 3.8169e-08 0.0007 3.8172e-08 0 3.8346e-08 0 3.8349e-08 0.0007 3.8352e-08 0 3.8526e-08 0 3.8529e-08 0.0007 3.8532e-08 0 3.8706e-08 0 3.8709e-08 0.0007 3.8712e-08 0 3.8886e-08 0 3.8889e-08 0.0007 3.8892e-08 0 3.9066e-08 0 3.9069e-08 0.0007 3.9072e-08 0 3.9246e-08 0 3.9249e-08 0.0007 3.9252e-08 0 3.9426e-08 0 3.9429e-08 0.0007 3.9432e-08 0 3.9606e-08 0 3.9609e-08 0.0007 3.9612e-08 0 3.9786e-08 0 3.9789e-08 0.0007 3.9792e-08 0 3.9966e-08 0 3.9969e-08 0.0007 3.9972e-08 0 4.0146e-08 0 4.0149e-08 0.0007 4.0152e-08 0 4.0326e-08 0 4.0329e-08 0.0007 4.0332e-08 0 4.0506e-08 0 4.0509e-08 0.0007 4.0512e-08 0 4.0686e-08 0 4.0689e-08 0.0007 4.0692e-08 0 4.0866e-08 0 4.0869e-08 0.0007 4.0872e-08 0 4.1046e-08 0 4.1049e-08 0.0007 4.1052e-08 0 4.1226e-08 0 4.1229e-08 0.0007 4.1232e-08 0 4.1406e-08 0 4.1409e-08 0.0007 4.1412e-08 0 4.1586e-08 0 4.1589e-08 0.0007 4.1592e-08 0 4.1766e-08 0 4.1769e-08 0.0007 4.1772e-08 0 4.1946e-08 0 4.1949e-08 0.0007 4.1952e-08 0 4.2126e-08 0 4.2129e-08 0.0007 4.2132e-08 0 4.2306e-08 0 4.2309e-08 0.0007 4.2312e-08 0 4.2486e-08 0 4.2489e-08 0.0007 4.2492e-08 0 4.2666e-08 0 4.2669e-08 0.0007 4.2672e-08 0 4.2846e-08 0 4.2849e-08 0.0007 4.2852e-08 0 4.3026e-08 0 4.3029e-08 0.0007 4.3032e-08 0 4.3206e-08 0 4.3209e-08 0.0007 4.3212e-08 0 4.3386e-08 0 4.3389e-08 0.0007 4.3392e-08 0 4.3566e-08 0 4.3569e-08 0.0007 4.3572e-08 0 4.3746e-08 0 4.3749e-08 0.0007 4.3752e-08 0 4.3926e-08 0 4.3929e-08 0.0007 4.3932e-08 0 4.4106e-08 0 4.4109e-08 0.0007 4.4112e-08 0 4.4286e-08 0 4.4289e-08 0.0007 4.4292e-08 0 4.4466e-08 0 4.4469e-08 0.0007 4.4472e-08 0 4.4646e-08 0 4.4649e-08 0.0007 4.4652e-08 0 4.4826e-08 0 4.4829e-08 0.0007 4.4832e-08 0 4.5006e-08 0 4.5009e-08 0.0007 4.5012e-08 0 4.5186e-08 0 4.5189e-08 0.0007 4.5192e-08 0 4.5366e-08 0 4.5369e-08 0.0007 4.5372e-08 0 4.5546e-08 0 4.5549e-08 0.0007 4.5552e-08 0 4.5726e-08 0 4.5729e-08 0.0007 4.5732e-08 0 4.5906e-08 0 4.5909e-08 0.0007 4.5912e-08 0)
B_DFF_IP3_12|1 _DFF_IP3_12|1 _DFF_IP3_12|2 JJMIT AREA=2.5
B_DFF_IP3_12|2 _DFF_IP3_12|4 _DFF_IP3_12|5 JJMIT AREA=1.61
B_DFF_IP3_12|3 _DFF_IP3_12|5 _DFF_IP3_12|6 JJMIT AREA=1.54
B_DFF_IP3_12|4 _DFF_IP3_12|8 _DFF_IP3_12|9 JJMIT AREA=1.69
B_DFF_IP3_12|5 _DFF_IP3_12|10 _DFF_IP3_12|8 JJMIT AREA=1.38
B_DFF_IP3_12|6 _DFF_IP3_12|11 _DFF_IP3_12|12 JJMIT AREA=2.5
B_DFF_IP3_12|7 _DFF_IP3_12|14 _DFF_IP3_12|15 JJMIT AREA=2.5
I_DFF_IP3_12|B1 0 _DFF_IP3_12|3  PWL(0 0 5e-12 0.000175)
I_DFF_IP3_12|B2 0 _DFF_IP3_12|7  PWL(0 0 5e-12 0.000173)
I_DFF_IP3_12|B3 0 _DFF_IP3_12|13  PWL(0 0 5e-12 0.000175)
I_DFF_IP3_12|B4 0 _DFF_IP3_12|16  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|B1 _DFF_IP3_12|3 _DFF_IP3_12|1  2e-12
L_DFF_IP3_12|B2 _DFF_IP3_12|7 _DFF_IP3_12|5  2e-12
L_DFF_IP3_12|B3 _DFF_IP3_12|11 _DFF_IP3_12|13  2e-12
L_DFF_IP3_12|B4 _DFF_IP3_12|16 _DFF_IP3_12|14  2e-12
L_DFF_IP3_12|1 IP3_1_OUT_RX _DFF_IP3_12|1  2.059e-12
L_DFF_IP3_12|2 _DFF_IP3_12|1 _DFF_IP3_12|4  4.123e-12
L_DFF_IP3_12|3 _DFF_IP3_12|5 _DFF_IP3_12|8  6.873e-12
L_DFF_IP3_12|4 _DFF_IP3_12|10 _DFF_IP3_12|11  5.195e-12
L_DFF_IP3_12|5 D13 _DFF_IP3_12|11  2.071e-12
L_DFF_IP3_12|6 _DFF_IP3_12|8 _DFF_IP3_12|14  3.287e-12
L_DFF_IP3_12|7 _DFF_IP3_12|14 IP3_2_OUT  2.066e-12
L_DFF_IP3_12|P1 _DFF_IP3_12|2 0  5.042e-13
L_DFF_IP3_12|P3 _DFF_IP3_12|6 0  5.799e-13
L_DFF_IP3_12|P4 _DFF_IP3_12|9 0  5.733e-13
L_DFF_IP3_12|P6 _DFF_IP3_12|12 0  4.605e-13
L_DFF_IP3_12|P7 _DFF_IP3_12|15 0  4.961e-13
R_DFF_IP3_12|B1 _DFF_IP3_12|1 _DFF_IP3_12|101  2.7439617672
L_DFF_IP3_12|RB1 _DFF_IP3_12|101 0  1.550338398468e-12
R_DFF_IP3_12|B2 _DFF_IP3_12|4 _DFF_IP3_12|104  4.260810197515528
L_DFF_IP3_12|RB2 _DFF_IP3_12|104 _DFF_IP3_12|5  2.407357761596273e-12
R_DFF_IP3_12|B3 _DFF_IP3_12|5 _DFF_IP3_12|105  4.454483388311688
L_DFF_IP3_12|RB3 _DFF_IP3_12|105 0  2.516783114396104e-12
R_DFF_IP3_12|B4 _DFF_IP3_12|8 _DFF_IP3_12|108  4.059115040236686
L_DFF_IP3_12|RB4 _DFF_IP3_12|108 0  2.2933999977337278e-12
R_DFF_IP3_12|B5 _DFF_IP3_12|10 _DFF_IP3_12|110  4.970945230434783
L_DFF_IP3_12|RB5 _DFF_IP3_12|110 _DFF_IP3_12|8  2.8085840551956523e-12
R_DFF_IP3_12|B6 _DFF_IP3_12|11 _DFF_IP3_12|111  2.7439617672
L_DFF_IP3_12|RB6 _DFF_IP3_12|111 0  1.550338398468e-12
R_DFF_IP3_12|B7 _DFF_IP3_12|14 _DFF_IP3_12|114  2.7439617672
L_DFF_IP3_12|RB7 _DFF_IP3_12|114 0  1.550338398468e-12
IT12|T 0 T12  PWL(0 0 1.5e-12 0 4.5e-12 0.0007 7.5e-12 0 1.815e-10 0 1.845e-10 0.0007 1.875e-10 0 3.615e-10 0 3.645e-10 0.0007 3.675e-10 0 5.415e-10 0 5.445e-10 0.0007 5.475e-10 0 7.215e-10 0 7.245e-10 0.0007 7.275e-10 0 9.015e-10 0 9.045e-10 0.0007 9.075e-10 0 1.0815e-09 0 1.0845e-09 0.0007 1.0875e-09 0 1.2615e-09 0 1.2645e-09 0.0007 1.2675e-09 0 1.4415e-09 0 1.4445e-09 0.0007 1.4475e-09 0 1.6215e-09 0 1.6245e-09 0.0007 1.6275e-09 0 1.8015e-09 0 1.8045e-09 0.0007 1.8075e-09 0 1.9815e-09 0 1.9845e-09 0.0007 1.9875e-09 0 2.1615e-09 0 2.1645e-09 0.0007 2.1675e-09 0 2.3415e-09 0 2.3445e-09 0.0007 2.3475e-09 0 2.5215e-09 0 2.5245e-09 0.0007 2.5275e-09 0 2.7015e-09 0 2.7045e-09 0.0007 2.7075e-09 0 2.8815e-09 0 2.8845e-09 0.0007 2.8875e-09 0 3.0615e-09 0 3.0645e-09 0.0007 3.0675e-09 0 3.2415e-09 0 3.2445e-09 0.0007 3.2475e-09 0 3.4215e-09 0 3.4245e-09 0.0007 3.4275e-09 0 3.6015e-09 0 3.6045e-09 0.0007 3.6075e-09 0 3.7815e-09 0 3.7845e-09 0.0007 3.7875e-09 0 3.9615e-09 0 3.9645e-09 0.0007 3.9675e-09 0 4.1415e-09 0 4.1445e-09 0.0007 4.1475e-09 0 4.3215e-09 0 4.3245e-09 0.0007 4.3275e-09 0 4.5015e-09 0 4.5045e-09 0.0007 4.5075e-09 0 4.6815e-09 0 4.6845e-09 0.0007 4.6875e-09 0 4.8615e-09 0 4.8645e-09 0.0007 4.8675e-09 0 5.0415e-09 0 5.0445e-09 0.0007 5.0475e-09 0 5.2215e-09 0 5.2245e-09 0.0007 5.2275e-09 0 5.4015e-09 0 5.4045e-09 0.0007 5.4075e-09 0 5.5815e-09 0 5.5845e-09 0.0007 5.5875e-09 0 5.7615e-09 0 5.7645e-09 0.0007 5.7675e-09 0 5.9415e-09 0 5.9445e-09 0.0007 5.9475e-09 0 6.1215e-09 0 6.1245e-09 0.0007 6.1275e-09 0 6.3015e-09 0 6.3045e-09 0.0007 6.3075e-09 0 6.4815e-09 0 6.4845e-09 0.0007 6.4875e-09 0 6.6615e-09 0 6.6645e-09 0.0007 6.6675e-09 0 6.8415e-09 0 6.8445e-09 0.0007 6.8475e-09 0 7.0215e-09 0 7.0245e-09 0.0007 7.0275e-09 0 7.2015e-09 0 7.2045e-09 0.0007 7.2075e-09 0 7.3815e-09 0 7.3845e-09 0.0007 7.3875e-09 0 7.5615e-09 0 7.5645e-09 0.0007 7.5675e-09 0 7.7415e-09 0 7.7445e-09 0.0007 7.7475e-09 0 7.9215e-09 0 7.9245e-09 0.0007 7.9275e-09 0 8.1015e-09 0 8.1045e-09 0.0007 8.1075e-09 0 8.2815e-09 0 8.2845e-09 0.0007 8.2875e-09 0 8.4615e-09 0 8.4645e-09 0.0007 8.4675e-09 0 8.6415e-09 0 8.6445e-09 0.0007 8.6475e-09 0 8.8215e-09 0 8.8245e-09 0.0007 8.8275e-09 0 9.0015e-09 0 9.0045e-09 0.0007 9.0075e-09 0 9.1815e-09 0 9.1845e-09 0.0007 9.1875e-09 0 9.3615e-09 0 9.3645e-09 0.0007 9.3675e-09 0 9.5415e-09 0 9.5445e-09 0.0007 9.5475e-09 0 9.7215e-09 0 9.7245e-09 0.0007 9.7275e-09 0 9.9015e-09 0 9.9045e-09 0.0007 9.9075e-09 0 1.00815e-08 0 1.00845e-08 0.0007 1.00875e-08 0 1.02615e-08 0 1.02645e-08 0.0007 1.02675e-08 0 1.04415e-08 0 1.04445e-08 0.0007 1.04475e-08 0 1.06215e-08 0 1.06245e-08 0.0007 1.06275e-08 0 1.08015e-08 0 1.08045e-08 0.0007 1.08075e-08 0 1.09815e-08 0 1.09845e-08 0.0007 1.09875e-08 0 1.11615e-08 0 1.11645e-08 0.0007 1.11675e-08 0 1.13415e-08 0 1.13445e-08 0.0007 1.13475e-08 0 1.15215e-08 0 1.15245e-08 0.0007 1.15275e-08 0 1.17015e-08 0 1.17045e-08 0.0007 1.17075e-08 0 1.18815e-08 0 1.18845e-08 0.0007 1.18875e-08 0 1.20615e-08 0 1.20645e-08 0.0007 1.20675e-08 0 1.22415e-08 0 1.22445e-08 0.0007 1.22475e-08 0 1.24215e-08 0 1.24245e-08 0.0007 1.24275e-08 0 1.26015e-08 0 1.26045e-08 0.0007 1.26075e-08 0 1.27815e-08 0 1.27845e-08 0.0007 1.27875e-08 0 1.29615e-08 0 1.29645e-08 0.0007 1.29675e-08 0 1.31415e-08 0 1.31445e-08 0.0007 1.31475e-08 0 1.33215e-08 0 1.33245e-08 0.0007 1.33275e-08 0 1.35015e-08 0 1.35045e-08 0.0007 1.35075e-08 0 1.36815e-08 0 1.36845e-08 0.0007 1.36875e-08 0 1.38615e-08 0 1.38645e-08 0.0007 1.38675e-08 0 1.40415e-08 0 1.40445e-08 0.0007 1.40475e-08 0 1.42215e-08 0 1.42245e-08 0.0007 1.42275e-08 0 1.44015e-08 0 1.44045e-08 0.0007 1.44075e-08 0 1.45815e-08 0 1.45845e-08 0.0007 1.45875e-08 0 1.47615e-08 0 1.47645e-08 0.0007 1.47675e-08 0 1.49415e-08 0 1.49445e-08 0.0007 1.49475e-08 0 1.51215e-08 0 1.51245e-08 0.0007 1.51275e-08 0 1.53015e-08 0 1.53045e-08 0.0007 1.53075e-08 0 1.54815e-08 0 1.54845e-08 0.0007 1.54875e-08 0 1.56615e-08 0 1.56645e-08 0.0007 1.56675e-08 0 1.58415e-08 0 1.58445e-08 0.0007 1.58475e-08 0 1.60215e-08 0 1.60245e-08 0.0007 1.60275e-08 0 1.62015e-08 0 1.62045e-08 0.0007 1.62075e-08 0 1.63815e-08 0 1.63845e-08 0.0007 1.63875e-08 0 1.65615e-08 0 1.65645e-08 0.0007 1.65675e-08 0 1.67415e-08 0 1.67445e-08 0.0007 1.67475e-08 0 1.69215e-08 0 1.69245e-08 0.0007 1.69275e-08 0 1.71015e-08 0 1.71045e-08 0.0007 1.71075e-08 0 1.72815e-08 0 1.72845e-08 0.0007 1.72875e-08 0 1.74615e-08 0 1.74645e-08 0.0007 1.74675e-08 0 1.76415e-08 0 1.76445e-08 0.0007 1.76475e-08 0 1.78215e-08 0 1.78245e-08 0.0007 1.78275e-08 0 1.80015e-08 0 1.80045e-08 0.0007 1.80075e-08 0 1.81815e-08 0 1.81845e-08 0.0007 1.81875e-08 0 1.83615e-08 0 1.83645e-08 0.0007 1.83675e-08 0 1.85415e-08 0 1.85445e-08 0.0007 1.85475e-08 0 1.87215e-08 0 1.87245e-08 0.0007 1.87275e-08 0 1.89015e-08 0 1.89045e-08 0.0007 1.89075e-08 0 1.90815e-08 0 1.90845e-08 0.0007 1.90875e-08 0 1.92615e-08 0 1.92645e-08 0.0007 1.92675e-08 0 1.94415e-08 0 1.94445e-08 0.0007 1.94475e-08 0 1.96215e-08 0 1.96245e-08 0.0007 1.96275e-08 0 1.98015e-08 0 1.98045e-08 0.0007 1.98075e-08 0 1.99815e-08 0 1.99845e-08 0.0007 1.99875e-08 0 2.01615e-08 0 2.01645e-08 0.0007 2.01675e-08 0 2.03415e-08 0 2.03445e-08 0.0007 2.03475e-08 0 2.05215e-08 0 2.05245e-08 0.0007 2.05275e-08 0 2.07015e-08 0 2.07045e-08 0.0007 2.07075e-08 0 2.08815e-08 0 2.08845e-08 0.0007 2.08875e-08 0 2.10615e-08 0 2.10645e-08 0.0007 2.10675e-08 0 2.12415e-08 0 2.12445e-08 0.0007 2.12475e-08 0 2.14215e-08 0 2.14245e-08 0.0007 2.14275e-08 0 2.16015e-08 0 2.16045e-08 0.0007 2.16075e-08 0 2.17815e-08 0 2.17845e-08 0.0007 2.17875e-08 0 2.19615e-08 0 2.19645e-08 0.0007 2.19675e-08 0 2.21415e-08 0 2.21445e-08 0.0007 2.21475e-08 0 2.23215e-08 0 2.23245e-08 0.0007 2.23275e-08 0 2.25015e-08 0 2.25045e-08 0.0007 2.25075e-08 0 2.26815e-08 0 2.26845e-08 0.0007 2.26875e-08 0 2.28615e-08 0 2.28645e-08 0.0007 2.28675e-08 0 2.30415e-08 0 2.30445e-08 0.0007 2.30475e-08 0 2.32215e-08 0 2.32245e-08 0.0007 2.32275e-08 0 2.34015e-08 0 2.34045e-08 0.0007 2.34075e-08 0 2.35815e-08 0 2.35845e-08 0.0007 2.35875e-08 0 2.37615e-08 0 2.37645e-08 0.0007 2.37675e-08 0 2.39415e-08 0 2.39445e-08 0.0007 2.39475e-08 0 2.41215e-08 0 2.41245e-08 0.0007 2.41275e-08 0 2.43015e-08 0 2.43045e-08 0.0007 2.43075e-08 0 2.44815e-08 0 2.44845e-08 0.0007 2.44875e-08 0 2.46615e-08 0 2.46645e-08 0.0007 2.46675e-08 0 2.48415e-08 0 2.48445e-08 0.0007 2.48475e-08 0 2.50215e-08 0 2.50245e-08 0.0007 2.50275e-08 0 2.52015e-08 0 2.52045e-08 0.0007 2.52075e-08 0 2.53815e-08 0 2.53845e-08 0.0007 2.53875e-08 0 2.55615e-08 0 2.55645e-08 0.0007 2.55675e-08 0 2.57415e-08 0 2.57445e-08 0.0007 2.57475e-08 0 2.59215e-08 0 2.59245e-08 0.0007 2.59275e-08 0 2.61015e-08 0 2.61045e-08 0.0007 2.61075e-08 0 2.62815e-08 0 2.62845e-08 0.0007 2.62875e-08 0 2.64615e-08 0 2.64645e-08 0.0007 2.64675e-08 0 2.66415e-08 0 2.66445e-08 0.0007 2.66475e-08 0 2.68215e-08 0 2.68245e-08 0.0007 2.68275e-08 0 2.70015e-08 0 2.70045e-08 0.0007 2.70075e-08 0 2.71815e-08 0 2.71845e-08 0.0007 2.71875e-08 0 2.73615e-08 0 2.73645e-08 0.0007 2.73675e-08 0 2.75415e-08 0 2.75445e-08 0.0007 2.75475e-08 0 2.77215e-08 0 2.77245e-08 0.0007 2.77275e-08 0 2.79015e-08 0 2.79045e-08 0.0007 2.79075e-08 0 2.80815e-08 0 2.80845e-08 0.0007 2.80875e-08 0 2.82615e-08 0 2.82645e-08 0.0007 2.82675e-08 0 2.84415e-08 0 2.84445e-08 0.0007 2.84475e-08 0 2.86215e-08 0 2.86245e-08 0.0007 2.86275e-08 0 2.88015e-08 0 2.88045e-08 0.0007 2.88075e-08 0 2.89815e-08 0 2.89845e-08 0.0007 2.89875e-08 0 2.91615e-08 0 2.91645e-08 0.0007 2.91675e-08 0 2.93415e-08 0 2.93445e-08 0.0007 2.93475e-08 0 2.95215e-08 0 2.95245e-08 0.0007 2.95275e-08 0 2.97015e-08 0 2.97045e-08 0.0007 2.97075e-08 0 2.98815e-08 0 2.98845e-08 0.0007 2.98875e-08 0 3.00615e-08 0 3.00645e-08 0.0007 3.00675e-08 0 3.02415e-08 0 3.02445e-08 0.0007 3.02475e-08 0 3.04215e-08 0 3.04245e-08 0.0007 3.04275e-08 0 3.06015e-08 0 3.06045e-08 0.0007 3.06075e-08 0 3.07815e-08 0 3.07845e-08 0.0007 3.07875e-08 0 3.09615e-08 0 3.09645e-08 0.0007 3.09675e-08 0 3.11415e-08 0 3.11445e-08 0.0007 3.11475e-08 0 3.13215e-08 0 3.13245e-08 0.0007 3.13275e-08 0 3.15015e-08 0 3.15045e-08 0.0007 3.15075e-08 0 3.16815e-08 0 3.16845e-08 0.0007 3.16875e-08 0 3.18615e-08 0 3.18645e-08 0.0007 3.18675e-08 0 3.20415e-08 0 3.20445e-08 0.0007 3.20475e-08 0 3.22215e-08 0 3.22245e-08 0.0007 3.22275e-08 0 3.24015e-08 0 3.24045e-08 0.0007 3.24075e-08 0 3.25815e-08 0 3.25845e-08 0.0007 3.25875e-08 0 3.27615e-08 0 3.27645e-08 0.0007 3.27675e-08 0 3.29415e-08 0 3.29445e-08 0.0007 3.29475e-08 0 3.31215e-08 0 3.31245e-08 0.0007 3.31275e-08 0 3.33015e-08 0 3.33045e-08 0.0007 3.33075e-08 0 3.34815e-08 0 3.34845e-08 0.0007 3.34875e-08 0 3.36615e-08 0 3.36645e-08 0.0007 3.36675e-08 0 3.38415e-08 0 3.38445e-08 0.0007 3.38475e-08 0 3.40215e-08 0 3.40245e-08 0.0007 3.40275e-08 0 3.42015e-08 0 3.42045e-08 0.0007 3.42075e-08 0 3.43815e-08 0 3.43845e-08 0.0007 3.43875e-08 0 3.45615e-08 0 3.45645e-08 0.0007 3.45675e-08 0 3.47415e-08 0 3.47445e-08 0.0007 3.47475e-08 0 3.49215e-08 0 3.49245e-08 0.0007 3.49275e-08 0 3.51015e-08 0 3.51045e-08 0.0007 3.51075e-08 0 3.52815e-08 0 3.52845e-08 0.0007 3.52875e-08 0 3.54615e-08 0 3.54645e-08 0.0007 3.54675e-08 0 3.56415e-08 0 3.56445e-08 0.0007 3.56475e-08 0 3.58215e-08 0 3.58245e-08 0.0007 3.58275e-08 0 3.60015e-08 0 3.60045e-08 0.0007 3.60075e-08 0 3.61815e-08 0 3.61845e-08 0.0007 3.61875e-08 0 3.63615e-08 0 3.63645e-08 0.0007 3.63675e-08 0 3.65415e-08 0 3.65445e-08 0.0007 3.65475e-08 0 3.67215e-08 0 3.67245e-08 0.0007 3.67275e-08 0 3.69015e-08 0 3.69045e-08 0.0007 3.69075e-08 0 3.70815e-08 0 3.70845e-08 0.0007 3.70875e-08 0 3.72615e-08 0 3.72645e-08 0.0007 3.72675e-08 0 3.74415e-08 0 3.74445e-08 0.0007 3.74475e-08 0 3.76215e-08 0 3.76245e-08 0.0007 3.76275e-08 0 3.78015e-08 0 3.78045e-08 0.0007 3.78075e-08 0 3.79815e-08 0 3.79845e-08 0.0007 3.79875e-08 0 3.81615e-08 0 3.81645e-08 0.0007 3.81675e-08 0 3.83415e-08 0 3.83445e-08 0.0007 3.83475e-08 0 3.85215e-08 0 3.85245e-08 0.0007 3.85275e-08 0 3.87015e-08 0 3.87045e-08 0.0007 3.87075e-08 0 3.88815e-08 0 3.88845e-08 0.0007 3.88875e-08 0 3.90615e-08 0 3.90645e-08 0.0007 3.90675e-08 0 3.92415e-08 0 3.92445e-08 0.0007 3.92475e-08 0 3.94215e-08 0 3.94245e-08 0.0007 3.94275e-08 0 3.96015e-08 0 3.96045e-08 0.0007 3.96075e-08 0 3.97815e-08 0 3.97845e-08 0.0007 3.97875e-08 0 3.99615e-08 0 3.99645e-08 0.0007 3.99675e-08 0 4.01415e-08 0 4.01445e-08 0.0007 4.01475e-08 0 4.03215e-08 0 4.03245e-08 0.0007 4.03275e-08 0 4.05015e-08 0 4.05045e-08 0.0007 4.05075e-08 0 4.06815e-08 0 4.06845e-08 0.0007 4.06875e-08 0 4.08615e-08 0 4.08645e-08 0.0007 4.08675e-08 0 4.10415e-08 0 4.10445e-08 0.0007 4.10475e-08 0 4.12215e-08 0 4.12245e-08 0.0007 4.12275e-08 0 4.14015e-08 0 4.14045e-08 0.0007 4.14075e-08 0 4.15815e-08 0 4.15845e-08 0.0007 4.15875e-08 0 4.17615e-08 0 4.17645e-08 0.0007 4.17675e-08 0 4.19415e-08 0 4.19445e-08 0.0007 4.19475e-08 0 4.21215e-08 0 4.21245e-08 0.0007 4.21275e-08 0 4.23015e-08 0 4.23045e-08 0.0007 4.23075e-08 0 4.24815e-08 0 4.24845e-08 0.0007 4.24875e-08 0 4.26615e-08 0 4.26645e-08 0.0007 4.26675e-08 0 4.28415e-08 0 4.28445e-08 0.0007 4.28475e-08 0 4.30215e-08 0 4.30245e-08 0.0007 4.30275e-08 0 4.32015e-08 0 4.32045e-08 0.0007 4.32075e-08 0 4.33815e-08 0 4.33845e-08 0.0007 4.33875e-08 0 4.35615e-08 0 4.35645e-08 0.0007 4.35675e-08 0 4.37415e-08 0 4.37445e-08 0.0007 4.37475e-08 0 4.39215e-08 0 4.39245e-08 0.0007 4.39275e-08 0 4.41015e-08 0 4.41045e-08 0.0007 4.41075e-08 0 4.42815e-08 0 4.42845e-08 0.0007 4.42875e-08 0 4.44615e-08 0 4.44645e-08 0.0007 4.44675e-08 0 4.46415e-08 0 4.46445e-08 0.0007 4.46475e-08 0 4.48215e-08 0 4.48245e-08 0.0007 4.48275e-08 0 4.50015e-08 0 4.50045e-08 0.0007 4.50075e-08 0 4.51815e-08 0 4.51845e-08 0.0007 4.51875e-08 0 4.53615e-08 0 4.53645e-08 0.0007 4.53675e-08 0 4.55415e-08 0 4.55445e-08 0.0007 4.55475e-08 0 4.57215e-08 0 4.57245e-08 0.0007 4.57275e-08 0 4.59015e-08 0 4.59045e-08 0.0007 4.59075e-08 0)
B_S0|1 _S0|1 _S0|2 JJMIT AREA=2.5
B_S0|2 _S0|4 _S0|5 JJMIT AREA=1.61
B_S0|3 _S0|5 _S0|6 JJMIT AREA=1.54
B_S0|4 _S0|8 _S0|9 JJMIT AREA=1.69
B_S0|5 _S0|10 _S0|8 JJMIT AREA=1.38
B_S0|6 _S0|11 _S0|12 JJMIT AREA=2.5
B_S0|7 _S0|14 _S0|15 JJMIT AREA=2.5
I_S0|B1 0 _S0|3  PWL(0 0 5e-12 0.000175)
I_S0|B2 0 _S0|7  PWL(0 0 5e-12 0.000173)
I_S0|B3 0 _S0|13  PWL(0 0 5e-12 0.000175)
I_S0|B4 0 _S0|16  PWL(0 0 5e-12 0.000175)
L_S0|B1 _S0|3 _S0|1  2e-12
L_S0|B2 _S0|7 _S0|5  2e-12
L_S0|B3 _S0|11 _S0|13  2e-12
L_S0|B4 _S0|16 _S0|14  2e-12
L_S0|1 P0_2_RX _S0|1  2.059e-12
L_S0|2 _S0|1 _S0|4  4.123e-12
L_S0|3 _S0|5 _S0|8  6.873e-12
L_S0|4 _S0|10 _S0|11  5.195e-12
L_S0|5 T12 _S0|11  2.071e-12
L_S0|6 _S0|8 _S0|14  3.287e-12
L_S0|7 _S0|14 S0  2.066e-12
L_S0|P1 _S0|2 0  5.042e-13
L_S0|P3 _S0|6 0  5.799e-13
L_S0|P4 _S0|9 0  5.733e-13
L_S0|P6 _S0|12 0  4.605e-13
L_S0|P7 _S0|15 0  4.961e-13
R_S0|B1 _S0|1 _S0|101  2.7439617672
L_S0|RB1 _S0|101 0  1.550338398468e-12
R_S0|B2 _S0|4 _S0|104  4.260810197515528
L_S0|RB2 _S0|104 _S0|5  2.407357761596273e-12
R_S0|B3 _S0|5 _S0|105  4.454483388311688
L_S0|RB3 _S0|105 0  2.516783114396104e-12
R_S0|B4 _S0|8 _S0|108  4.059115040236686
L_S0|RB4 _S0|108 0  2.2933999977337278e-12
R_S0|B5 _S0|10 _S0|110  4.970945230434783
L_S0|RB5 _S0|110 _S0|8  2.8085840551956523e-12
R_S0|B6 _S0|11 _S0|111  2.7439617672
L_S0|RB6 _S0|111 0  1.550338398468e-12
R_S0|B7 _S0|14 _S0|114  2.7439617672
L_S0|RB7 _S0|114 0  1.550338398468e-12
IT13|T 0 T13  PWL(0 0 1.5e-12 0 4.5e-12 0.0007 7.5e-12 0 1.815e-10 0 1.845e-10 0.0007 1.875e-10 0 3.615e-10 0 3.645e-10 0.0007 3.675e-10 0 5.415e-10 0 5.445e-10 0.0007 5.475e-10 0 7.215e-10 0 7.245e-10 0.0007 7.275e-10 0 9.015e-10 0 9.045e-10 0.0007 9.075e-10 0 1.0815e-09 0 1.0845e-09 0.0007 1.0875e-09 0 1.2615e-09 0 1.2645e-09 0.0007 1.2675e-09 0 1.4415e-09 0 1.4445e-09 0.0007 1.4475e-09 0 1.6215e-09 0 1.6245e-09 0.0007 1.6275e-09 0 1.8015e-09 0 1.8045e-09 0.0007 1.8075e-09 0 1.9815e-09 0 1.9845e-09 0.0007 1.9875e-09 0 2.1615e-09 0 2.1645e-09 0.0007 2.1675e-09 0 2.3415e-09 0 2.3445e-09 0.0007 2.3475e-09 0 2.5215e-09 0 2.5245e-09 0.0007 2.5275e-09 0 2.7015e-09 0 2.7045e-09 0.0007 2.7075e-09 0 2.8815e-09 0 2.8845e-09 0.0007 2.8875e-09 0 3.0615e-09 0 3.0645e-09 0.0007 3.0675e-09 0 3.2415e-09 0 3.2445e-09 0.0007 3.2475e-09 0 3.4215e-09 0 3.4245e-09 0.0007 3.4275e-09 0 3.6015e-09 0 3.6045e-09 0.0007 3.6075e-09 0 3.7815e-09 0 3.7845e-09 0.0007 3.7875e-09 0 3.9615e-09 0 3.9645e-09 0.0007 3.9675e-09 0 4.1415e-09 0 4.1445e-09 0.0007 4.1475e-09 0 4.3215e-09 0 4.3245e-09 0.0007 4.3275e-09 0 4.5015e-09 0 4.5045e-09 0.0007 4.5075e-09 0 4.6815e-09 0 4.6845e-09 0.0007 4.6875e-09 0 4.8615e-09 0 4.8645e-09 0.0007 4.8675e-09 0 5.0415e-09 0 5.0445e-09 0.0007 5.0475e-09 0 5.2215e-09 0 5.2245e-09 0.0007 5.2275e-09 0 5.4015e-09 0 5.4045e-09 0.0007 5.4075e-09 0 5.5815e-09 0 5.5845e-09 0.0007 5.5875e-09 0 5.7615e-09 0 5.7645e-09 0.0007 5.7675e-09 0 5.9415e-09 0 5.9445e-09 0.0007 5.9475e-09 0 6.1215e-09 0 6.1245e-09 0.0007 6.1275e-09 0 6.3015e-09 0 6.3045e-09 0.0007 6.3075e-09 0 6.4815e-09 0 6.4845e-09 0.0007 6.4875e-09 0 6.6615e-09 0 6.6645e-09 0.0007 6.6675e-09 0 6.8415e-09 0 6.8445e-09 0.0007 6.8475e-09 0 7.0215e-09 0 7.0245e-09 0.0007 7.0275e-09 0 7.2015e-09 0 7.2045e-09 0.0007 7.2075e-09 0 7.3815e-09 0 7.3845e-09 0.0007 7.3875e-09 0 7.5615e-09 0 7.5645e-09 0.0007 7.5675e-09 0 7.7415e-09 0 7.7445e-09 0.0007 7.7475e-09 0 7.9215e-09 0 7.9245e-09 0.0007 7.9275e-09 0 8.1015e-09 0 8.1045e-09 0.0007 8.1075e-09 0 8.2815e-09 0 8.2845e-09 0.0007 8.2875e-09 0 8.4615e-09 0 8.4645e-09 0.0007 8.4675e-09 0 8.6415e-09 0 8.6445e-09 0.0007 8.6475e-09 0 8.8215e-09 0 8.8245e-09 0.0007 8.8275e-09 0 9.0015e-09 0 9.0045e-09 0.0007 9.0075e-09 0 9.1815e-09 0 9.1845e-09 0.0007 9.1875e-09 0 9.3615e-09 0 9.3645e-09 0.0007 9.3675e-09 0 9.5415e-09 0 9.5445e-09 0.0007 9.5475e-09 0 9.7215e-09 0 9.7245e-09 0.0007 9.7275e-09 0 9.9015e-09 0 9.9045e-09 0.0007 9.9075e-09 0 1.00815e-08 0 1.00845e-08 0.0007 1.00875e-08 0 1.02615e-08 0 1.02645e-08 0.0007 1.02675e-08 0 1.04415e-08 0 1.04445e-08 0.0007 1.04475e-08 0 1.06215e-08 0 1.06245e-08 0.0007 1.06275e-08 0 1.08015e-08 0 1.08045e-08 0.0007 1.08075e-08 0 1.09815e-08 0 1.09845e-08 0.0007 1.09875e-08 0 1.11615e-08 0 1.11645e-08 0.0007 1.11675e-08 0 1.13415e-08 0 1.13445e-08 0.0007 1.13475e-08 0 1.15215e-08 0 1.15245e-08 0.0007 1.15275e-08 0 1.17015e-08 0 1.17045e-08 0.0007 1.17075e-08 0 1.18815e-08 0 1.18845e-08 0.0007 1.18875e-08 0 1.20615e-08 0 1.20645e-08 0.0007 1.20675e-08 0 1.22415e-08 0 1.22445e-08 0.0007 1.22475e-08 0 1.24215e-08 0 1.24245e-08 0.0007 1.24275e-08 0 1.26015e-08 0 1.26045e-08 0.0007 1.26075e-08 0 1.27815e-08 0 1.27845e-08 0.0007 1.27875e-08 0 1.29615e-08 0 1.29645e-08 0.0007 1.29675e-08 0 1.31415e-08 0 1.31445e-08 0.0007 1.31475e-08 0 1.33215e-08 0 1.33245e-08 0.0007 1.33275e-08 0 1.35015e-08 0 1.35045e-08 0.0007 1.35075e-08 0 1.36815e-08 0 1.36845e-08 0.0007 1.36875e-08 0 1.38615e-08 0 1.38645e-08 0.0007 1.38675e-08 0 1.40415e-08 0 1.40445e-08 0.0007 1.40475e-08 0 1.42215e-08 0 1.42245e-08 0.0007 1.42275e-08 0 1.44015e-08 0 1.44045e-08 0.0007 1.44075e-08 0 1.45815e-08 0 1.45845e-08 0.0007 1.45875e-08 0 1.47615e-08 0 1.47645e-08 0.0007 1.47675e-08 0 1.49415e-08 0 1.49445e-08 0.0007 1.49475e-08 0 1.51215e-08 0 1.51245e-08 0.0007 1.51275e-08 0 1.53015e-08 0 1.53045e-08 0.0007 1.53075e-08 0 1.54815e-08 0 1.54845e-08 0.0007 1.54875e-08 0 1.56615e-08 0 1.56645e-08 0.0007 1.56675e-08 0 1.58415e-08 0 1.58445e-08 0.0007 1.58475e-08 0 1.60215e-08 0 1.60245e-08 0.0007 1.60275e-08 0 1.62015e-08 0 1.62045e-08 0.0007 1.62075e-08 0 1.63815e-08 0 1.63845e-08 0.0007 1.63875e-08 0 1.65615e-08 0 1.65645e-08 0.0007 1.65675e-08 0 1.67415e-08 0 1.67445e-08 0.0007 1.67475e-08 0 1.69215e-08 0 1.69245e-08 0.0007 1.69275e-08 0 1.71015e-08 0 1.71045e-08 0.0007 1.71075e-08 0 1.72815e-08 0 1.72845e-08 0.0007 1.72875e-08 0 1.74615e-08 0 1.74645e-08 0.0007 1.74675e-08 0 1.76415e-08 0 1.76445e-08 0.0007 1.76475e-08 0 1.78215e-08 0 1.78245e-08 0.0007 1.78275e-08 0 1.80015e-08 0 1.80045e-08 0.0007 1.80075e-08 0 1.81815e-08 0 1.81845e-08 0.0007 1.81875e-08 0 1.83615e-08 0 1.83645e-08 0.0007 1.83675e-08 0 1.85415e-08 0 1.85445e-08 0.0007 1.85475e-08 0 1.87215e-08 0 1.87245e-08 0.0007 1.87275e-08 0 1.89015e-08 0 1.89045e-08 0.0007 1.89075e-08 0 1.90815e-08 0 1.90845e-08 0.0007 1.90875e-08 0 1.92615e-08 0 1.92645e-08 0.0007 1.92675e-08 0 1.94415e-08 0 1.94445e-08 0.0007 1.94475e-08 0 1.96215e-08 0 1.96245e-08 0.0007 1.96275e-08 0 1.98015e-08 0 1.98045e-08 0.0007 1.98075e-08 0 1.99815e-08 0 1.99845e-08 0.0007 1.99875e-08 0 2.01615e-08 0 2.01645e-08 0.0007 2.01675e-08 0 2.03415e-08 0 2.03445e-08 0.0007 2.03475e-08 0 2.05215e-08 0 2.05245e-08 0.0007 2.05275e-08 0 2.07015e-08 0 2.07045e-08 0.0007 2.07075e-08 0 2.08815e-08 0 2.08845e-08 0.0007 2.08875e-08 0 2.10615e-08 0 2.10645e-08 0.0007 2.10675e-08 0 2.12415e-08 0 2.12445e-08 0.0007 2.12475e-08 0 2.14215e-08 0 2.14245e-08 0.0007 2.14275e-08 0 2.16015e-08 0 2.16045e-08 0.0007 2.16075e-08 0 2.17815e-08 0 2.17845e-08 0.0007 2.17875e-08 0 2.19615e-08 0 2.19645e-08 0.0007 2.19675e-08 0 2.21415e-08 0 2.21445e-08 0.0007 2.21475e-08 0 2.23215e-08 0 2.23245e-08 0.0007 2.23275e-08 0 2.25015e-08 0 2.25045e-08 0.0007 2.25075e-08 0 2.26815e-08 0 2.26845e-08 0.0007 2.26875e-08 0 2.28615e-08 0 2.28645e-08 0.0007 2.28675e-08 0 2.30415e-08 0 2.30445e-08 0.0007 2.30475e-08 0 2.32215e-08 0 2.32245e-08 0.0007 2.32275e-08 0 2.34015e-08 0 2.34045e-08 0.0007 2.34075e-08 0 2.35815e-08 0 2.35845e-08 0.0007 2.35875e-08 0 2.37615e-08 0 2.37645e-08 0.0007 2.37675e-08 0 2.39415e-08 0 2.39445e-08 0.0007 2.39475e-08 0 2.41215e-08 0 2.41245e-08 0.0007 2.41275e-08 0 2.43015e-08 0 2.43045e-08 0.0007 2.43075e-08 0 2.44815e-08 0 2.44845e-08 0.0007 2.44875e-08 0 2.46615e-08 0 2.46645e-08 0.0007 2.46675e-08 0 2.48415e-08 0 2.48445e-08 0.0007 2.48475e-08 0 2.50215e-08 0 2.50245e-08 0.0007 2.50275e-08 0 2.52015e-08 0 2.52045e-08 0.0007 2.52075e-08 0 2.53815e-08 0 2.53845e-08 0.0007 2.53875e-08 0 2.55615e-08 0 2.55645e-08 0.0007 2.55675e-08 0 2.57415e-08 0 2.57445e-08 0.0007 2.57475e-08 0 2.59215e-08 0 2.59245e-08 0.0007 2.59275e-08 0 2.61015e-08 0 2.61045e-08 0.0007 2.61075e-08 0 2.62815e-08 0 2.62845e-08 0.0007 2.62875e-08 0 2.64615e-08 0 2.64645e-08 0.0007 2.64675e-08 0 2.66415e-08 0 2.66445e-08 0.0007 2.66475e-08 0 2.68215e-08 0 2.68245e-08 0.0007 2.68275e-08 0 2.70015e-08 0 2.70045e-08 0.0007 2.70075e-08 0 2.71815e-08 0 2.71845e-08 0.0007 2.71875e-08 0 2.73615e-08 0 2.73645e-08 0.0007 2.73675e-08 0 2.75415e-08 0 2.75445e-08 0.0007 2.75475e-08 0 2.77215e-08 0 2.77245e-08 0.0007 2.77275e-08 0 2.79015e-08 0 2.79045e-08 0.0007 2.79075e-08 0 2.80815e-08 0 2.80845e-08 0.0007 2.80875e-08 0 2.82615e-08 0 2.82645e-08 0.0007 2.82675e-08 0 2.84415e-08 0 2.84445e-08 0.0007 2.84475e-08 0 2.86215e-08 0 2.86245e-08 0.0007 2.86275e-08 0 2.88015e-08 0 2.88045e-08 0.0007 2.88075e-08 0 2.89815e-08 0 2.89845e-08 0.0007 2.89875e-08 0 2.91615e-08 0 2.91645e-08 0.0007 2.91675e-08 0 2.93415e-08 0 2.93445e-08 0.0007 2.93475e-08 0 2.95215e-08 0 2.95245e-08 0.0007 2.95275e-08 0 2.97015e-08 0 2.97045e-08 0.0007 2.97075e-08 0 2.98815e-08 0 2.98845e-08 0.0007 2.98875e-08 0 3.00615e-08 0 3.00645e-08 0.0007 3.00675e-08 0 3.02415e-08 0 3.02445e-08 0.0007 3.02475e-08 0 3.04215e-08 0 3.04245e-08 0.0007 3.04275e-08 0 3.06015e-08 0 3.06045e-08 0.0007 3.06075e-08 0 3.07815e-08 0 3.07845e-08 0.0007 3.07875e-08 0 3.09615e-08 0 3.09645e-08 0.0007 3.09675e-08 0 3.11415e-08 0 3.11445e-08 0.0007 3.11475e-08 0 3.13215e-08 0 3.13245e-08 0.0007 3.13275e-08 0 3.15015e-08 0 3.15045e-08 0.0007 3.15075e-08 0 3.16815e-08 0 3.16845e-08 0.0007 3.16875e-08 0 3.18615e-08 0 3.18645e-08 0.0007 3.18675e-08 0 3.20415e-08 0 3.20445e-08 0.0007 3.20475e-08 0 3.22215e-08 0 3.22245e-08 0.0007 3.22275e-08 0 3.24015e-08 0 3.24045e-08 0.0007 3.24075e-08 0 3.25815e-08 0 3.25845e-08 0.0007 3.25875e-08 0 3.27615e-08 0 3.27645e-08 0.0007 3.27675e-08 0 3.29415e-08 0 3.29445e-08 0.0007 3.29475e-08 0 3.31215e-08 0 3.31245e-08 0.0007 3.31275e-08 0 3.33015e-08 0 3.33045e-08 0.0007 3.33075e-08 0 3.34815e-08 0 3.34845e-08 0.0007 3.34875e-08 0 3.36615e-08 0 3.36645e-08 0.0007 3.36675e-08 0 3.38415e-08 0 3.38445e-08 0.0007 3.38475e-08 0 3.40215e-08 0 3.40245e-08 0.0007 3.40275e-08 0 3.42015e-08 0 3.42045e-08 0.0007 3.42075e-08 0 3.43815e-08 0 3.43845e-08 0.0007 3.43875e-08 0 3.45615e-08 0 3.45645e-08 0.0007 3.45675e-08 0 3.47415e-08 0 3.47445e-08 0.0007 3.47475e-08 0 3.49215e-08 0 3.49245e-08 0.0007 3.49275e-08 0 3.51015e-08 0 3.51045e-08 0.0007 3.51075e-08 0 3.52815e-08 0 3.52845e-08 0.0007 3.52875e-08 0 3.54615e-08 0 3.54645e-08 0.0007 3.54675e-08 0 3.56415e-08 0 3.56445e-08 0.0007 3.56475e-08 0 3.58215e-08 0 3.58245e-08 0.0007 3.58275e-08 0 3.60015e-08 0 3.60045e-08 0.0007 3.60075e-08 0 3.61815e-08 0 3.61845e-08 0.0007 3.61875e-08 0 3.63615e-08 0 3.63645e-08 0.0007 3.63675e-08 0 3.65415e-08 0 3.65445e-08 0.0007 3.65475e-08 0 3.67215e-08 0 3.67245e-08 0.0007 3.67275e-08 0 3.69015e-08 0 3.69045e-08 0.0007 3.69075e-08 0 3.70815e-08 0 3.70845e-08 0.0007 3.70875e-08 0 3.72615e-08 0 3.72645e-08 0.0007 3.72675e-08 0 3.74415e-08 0 3.74445e-08 0.0007 3.74475e-08 0 3.76215e-08 0 3.76245e-08 0.0007 3.76275e-08 0 3.78015e-08 0 3.78045e-08 0.0007 3.78075e-08 0 3.79815e-08 0 3.79845e-08 0.0007 3.79875e-08 0 3.81615e-08 0 3.81645e-08 0.0007 3.81675e-08 0 3.83415e-08 0 3.83445e-08 0.0007 3.83475e-08 0 3.85215e-08 0 3.85245e-08 0.0007 3.85275e-08 0 3.87015e-08 0 3.87045e-08 0.0007 3.87075e-08 0 3.88815e-08 0 3.88845e-08 0.0007 3.88875e-08 0 3.90615e-08 0 3.90645e-08 0.0007 3.90675e-08 0 3.92415e-08 0 3.92445e-08 0.0007 3.92475e-08 0 3.94215e-08 0 3.94245e-08 0.0007 3.94275e-08 0 3.96015e-08 0 3.96045e-08 0.0007 3.96075e-08 0 3.97815e-08 0 3.97845e-08 0.0007 3.97875e-08 0 3.99615e-08 0 3.99645e-08 0.0007 3.99675e-08 0 4.01415e-08 0 4.01445e-08 0.0007 4.01475e-08 0 4.03215e-08 0 4.03245e-08 0.0007 4.03275e-08 0 4.05015e-08 0 4.05045e-08 0.0007 4.05075e-08 0 4.06815e-08 0 4.06845e-08 0.0007 4.06875e-08 0 4.08615e-08 0 4.08645e-08 0.0007 4.08675e-08 0 4.10415e-08 0 4.10445e-08 0.0007 4.10475e-08 0 4.12215e-08 0 4.12245e-08 0.0007 4.12275e-08 0 4.14015e-08 0 4.14045e-08 0.0007 4.14075e-08 0 4.15815e-08 0 4.15845e-08 0.0007 4.15875e-08 0 4.17615e-08 0 4.17645e-08 0.0007 4.17675e-08 0 4.19415e-08 0 4.19445e-08 0.0007 4.19475e-08 0 4.21215e-08 0 4.21245e-08 0.0007 4.21275e-08 0 4.23015e-08 0 4.23045e-08 0.0007 4.23075e-08 0 4.24815e-08 0 4.24845e-08 0.0007 4.24875e-08 0 4.26615e-08 0 4.26645e-08 0.0007 4.26675e-08 0 4.28415e-08 0 4.28445e-08 0.0007 4.28475e-08 0 4.30215e-08 0 4.30245e-08 0.0007 4.30275e-08 0 4.32015e-08 0 4.32045e-08 0.0007 4.32075e-08 0 4.33815e-08 0 4.33845e-08 0.0007 4.33875e-08 0 4.35615e-08 0 4.35645e-08 0.0007 4.35675e-08 0 4.37415e-08 0 4.37445e-08 0.0007 4.37475e-08 0 4.39215e-08 0 4.39245e-08 0.0007 4.39275e-08 0 4.41015e-08 0 4.41045e-08 0.0007 4.41075e-08 0 4.42815e-08 0 4.42845e-08 0.0007 4.42875e-08 0 4.44615e-08 0 4.44645e-08 0.0007 4.44675e-08 0 4.46415e-08 0 4.46445e-08 0.0007 4.46475e-08 0 4.48215e-08 0 4.48245e-08 0.0007 4.48275e-08 0 4.50015e-08 0 4.50045e-08 0.0007 4.50075e-08 0 4.51815e-08 0 4.51845e-08 0.0007 4.51875e-08 0 4.53615e-08 0 4.53645e-08 0.0007 4.53675e-08 0 4.55415e-08 0 4.55445e-08 0.0007 4.55475e-08 0 4.57215e-08 0 4.57245e-08 0.0007 4.57275e-08 0 4.59015e-08 0 4.59045e-08 0.0007 4.59075e-08 0)
B_S1|1 _S1|1 _S1|2 JJMIT AREA=2.5
B_S1|2 _S1|4 _S1|5 JJMIT AREA=2.09
B_S1|3 _S1|25 _S1|6 JJMIT AREA=1.71
B_S1|4 _S1|9 _S1|10 JJMIT AREA=2.5
B_S1|5 _S1|12 _S1|13 JJMIT AREA=2.09
B_S1|6 _S1|26 _S1|14 JJMIT AREA=1.71
B_S1|7 _S1|27 _S1|16 JJMIT AREA=1.62
B_S1|8 _S1|17 _S1|18 JJMIT AREA=2.5
B_S1|9 _S1|20 _S1|16 JJMIT AREA=1.45
B_S1|10 _S1|16 _S1|21 JJMIT AREA=0.89
B_S1|11 _S1|22 _S1|23 JJMIT AREA=2.5
I_S1|B1 0 _S1|3  PWL(0 0 5e-12 0.000175)
I_S1|B2 0 _S1|7  PWL(0 0 5e-12 0.000112)
I_S1|B3 0 _S1|11  PWL(0 0 5e-12 0.000175)
I_S1|B4 0 _S1|15  PWL(0 0 5e-12 0.000112)
I_S1|B5 0 _S1|19  PWL(0 0 5e-12 0.000175)
I_S1|B6 0 _S1|24  PWL(0 0 5e-12 0.000175)
L_S1|B1 _S1|3 _S1|1  2e-12
L_S1|B2 _S1|7 _S1|6  2e-12
L_S1|B3 _S1|11 _S1|9  2e-12
L_S1|B4 _S1|15 _S1|14  2e-12
L_S1|B5 _S1|19 _S1|17  2e-12
L_S1|B6 _S1|24 _S1|22  2e-12
L_S1|1 G0_2_RX _S1|1  2.06e-12
L_S1|2 _S1|1 _S1|4  3.233e-12
L_S1|3 _S1|4 _S1|25  1.419e-12
L_S1|4 _S1|6 _S1|8  6.051e-12
L_S1|5 IP1_2_OUT_RX _S1|9  2.092e-12
L_S1|6 _S1|9 _S1|12  3.221e-12
L_S1|7 _S1|12 _S1|26  1.384e-12
L_S1|8 _S1|14 _S1|8  6.059e-12
L_S1|9 _S1|8 _S1|27  1.301e-12
L_S1|10 T13 _S1|17  2.082e-12
L_S1|11 _S1|17 _S1|20  1.43e-12
L_S1|12 _S1|16 _S1|22  3.892e-12
L_S1|13 _S1|22 S1  2.077e-12
L_S1|P1 _S1|2 0  5.508e-13
L_S1|P2 _S1|5 0  4.769e-13
L_S1|P4 _S1|10 0  4.767e-13
L_S1|P5 _S1|13 0  4.812e-13
L_S1|P8 _S1|18 0  4.526e-13
L_S1|P10 _S1|21 0  5.69e-13
L_S1|P11 _S1|23 0  4.746e-13
R_S1|B1 _S1|1 _S1|101  2.7439617672
L_S1|RB1 _S1|101 0  2.050338398468e-12
R_S1|B2 _S1|4 _S1|104  3.2822509177033496
L_S1|RB2 _S1|104 0  2.3544717685023925e-12
R_S1|B3 _S1|4 _S1|106  4.011640010526316
L_S1|RB3 _S1|106 _S1|6  2.766576605947368e-12
R_S1|B4 _S1|9 _S1|109  2.7439617672
L_S1|RB4 _S1|109 0  2.050338398468e-12
R_S1|B5 _S1|12 _S1|112  3.2822509177033496
L_S1|RB5 _S1|112 0  2.3544717685023925e-12
R_S1|B6 _S1|12 _S1|114  4.011640010526316
L_S1|RB6 _S1|114 _S1|14  2.766576605947368e-12
R_S1|B7 _S1|8 _S1|108  4.2345089
L_S1|RB7 _S1|108 _S1|16  2.8924975284999997e-12
R_S1|B8 _S1|17 _S1|117  2.7439617672
L_S1|RB8 _S1|117 0  2.050338398468e-12
R_S1|B9 _S1|20 _S1|120  4.730968564137931
L_S1|RB9 _S1|120 _S1|16  3.172997238737931e-12
R_S1|B10 _S1|16 _S1|116  7.707757773033708
L_S1|RB10 _S1|116 0  4.854883141764045e-12
R_S1|B11 _S1|22 _S1|122  2.7439617672
L_S1|RB11 _S1|122 0  2.050338398468e-12
IT14|T 0 T14  PWL(0 0 1.5e-12 0 4.5e-12 0.0007 7.5e-12 0 1.815e-10 0 1.845e-10 0.0007 1.875e-10 0 3.615e-10 0 3.645e-10 0.0007 3.675e-10 0 5.415e-10 0 5.445e-10 0.0007 5.475e-10 0 7.215e-10 0 7.245e-10 0.0007 7.275e-10 0 9.015e-10 0 9.045e-10 0.0007 9.075e-10 0 1.0815e-09 0 1.0845e-09 0.0007 1.0875e-09 0 1.2615e-09 0 1.2645e-09 0.0007 1.2675e-09 0 1.4415e-09 0 1.4445e-09 0.0007 1.4475e-09 0 1.6215e-09 0 1.6245e-09 0.0007 1.6275e-09 0 1.8015e-09 0 1.8045e-09 0.0007 1.8075e-09 0 1.9815e-09 0 1.9845e-09 0.0007 1.9875e-09 0 2.1615e-09 0 2.1645e-09 0.0007 2.1675e-09 0 2.3415e-09 0 2.3445e-09 0.0007 2.3475e-09 0 2.5215e-09 0 2.5245e-09 0.0007 2.5275e-09 0 2.7015e-09 0 2.7045e-09 0.0007 2.7075e-09 0 2.8815e-09 0 2.8845e-09 0.0007 2.8875e-09 0 3.0615e-09 0 3.0645e-09 0.0007 3.0675e-09 0 3.2415e-09 0 3.2445e-09 0.0007 3.2475e-09 0 3.4215e-09 0 3.4245e-09 0.0007 3.4275e-09 0 3.6015e-09 0 3.6045e-09 0.0007 3.6075e-09 0 3.7815e-09 0 3.7845e-09 0.0007 3.7875e-09 0 3.9615e-09 0 3.9645e-09 0.0007 3.9675e-09 0 4.1415e-09 0 4.1445e-09 0.0007 4.1475e-09 0 4.3215e-09 0 4.3245e-09 0.0007 4.3275e-09 0 4.5015e-09 0 4.5045e-09 0.0007 4.5075e-09 0 4.6815e-09 0 4.6845e-09 0.0007 4.6875e-09 0 4.8615e-09 0 4.8645e-09 0.0007 4.8675e-09 0 5.0415e-09 0 5.0445e-09 0.0007 5.0475e-09 0 5.2215e-09 0 5.2245e-09 0.0007 5.2275e-09 0 5.4015e-09 0 5.4045e-09 0.0007 5.4075e-09 0 5.5815e-09 0 5.5845e-09 0.0007 5.5875e-09 0 5.7615e-09 0 5.7645e-09 0.0007 5.7675e-09 0 5.9415e-09 0 5.9445e-09 0.0007 5.9475e-09 0 6.1215e-09 0 6.1245e-09 0.0007 6.1275e-09 0 6.3015e-09 0 6.3045e-09 0.0007 6.3075e-09 0 6.4815e-09 0 6.4845e-09 0.0007 6.4875e-09 0 6.6615e-09 0 6.6645e-09 0.0007 6.6675e-09 0 6.8415e-09 0 6.8445e-09 0.0007 6.8475e-09 0 7.0215e-09 0 7.0245e-09 0.0007 7.0275e-09 0 7.2015e-09 0 7.2045e-09 0.0007 7.2075e-09 0 7.3815e-09 0 7.3845e-09 0.0007 7.3875e-09 0 7.5615e-09 0 7.5645e-09 0.0007 7.5675e-09 0 7.7415e-09 0 7.7445e-09 0.0007 7.7475e-09 0 7.9215e-09 0 7.9245e-09 0.0007 7.9275e-09 0 8.1015e-09 0 8.1045e-09 0.0007 8.1075e-09 0 8.2815e-09 0 8.2845e-09 0.0007 8.2875e-09 0 8.4615e-09 0 8.4645e-09 0.0007 8.4675e-09 0 8.6415e-09 0 8.6445e-09 0.0007 8.6475e-09 0 8.8215e-09 0 8.8245e-09 0.0007 8.8275e-09 0 9.0015e-09 0 9.0045e-09 0.0007 9.0075e-09 0 9.1815e-09 0 9.1845e-09 0.0007 9.1875e-09 0 9.3615e-09 0 9.3645e-09 0.0007 9.3675e-09 0 9.5415e-09 0 9.5445e-09 0.0007 9.5475e-09 0 9.7215e-09 0 9.7245e-09 0.0007 9.7275e-09 0 9.9015e-09 0 9.9045e-09 0.0007 9.9075e-09 0 1.00815e-08 0 1.00845e-08 0.0007 1.00875e-08 0 1.02615e-08 0 1.02645e-08 0.0007 1.02675e-08 0 1.04415e-08 0 1.04445e-08 0.0007 1.04475e-08 0 1.06215e-08 0 1.06245e-08 0.0007 1.06275e-08 0 1.08015e-08 0 1.08045e-08 0.0007 1.08075e-08 0 1.09815e-08 0 1.09845e-08 0.0007 1.09875e-08 0 1.11615e-08 0 1.11645e-08 0.0007 1.11675e-08 0 1.13415e-08 0 1.13445e-08 0.0007 1.13475e-08 0 1.15215e-08 0 1.15245e-08 0.0007 1.15275e-08 0 1.17015e-08 0 1.17045e-08 0.0007 1.17075e-08 0 1.18815e-08 0 1.18845e-08 0.0007 1.18875e-08 0 1.20615e-08 0 1.20645e-08 0.0007 1.20675e-08 0 1.22415e-08 0 1.22445e-08 0.0007 1.22475e-08 0 1.24215e-08 0 1.24245e-08 0.0007 1.24275e-08 0 1.26015e-08 0 1.26045e-08 0.0007 1.26075e-08 0 1.27815e-08 0 1.27845e-08 0.0007 1.27875e-08 0 1.29615e-08 0 1.29645e-08 0.0007 1.29675e-08 0 1.31415e-08 0 1.31445e-08 0.0007 1.31475e-08 0 1.33215e-08 0 1.33245e-08 0.0007 1.33275e-08 0 1.35015e-08 0 1.35045e-08 0.0007 1.35075e-08 0 1.36815e-08 0 1.36845e-08 0.0007 1.36875e-08 0 1.38615e-08 0 1.38645e-08 0.0007 1.38675e-08 0 1.40415e-08 0 1.40445e-08 0.0007 1.40475e-08 0 1.42215e-08 0 1.42245e-08 0.0007 1.42275e-08 0 1.44015e-08 0 1.44045e-08 0.0007 1.44075e-08 0 1.45815e-08 0 1.45845e-08 0.0007 1.45875e-08 0 1.47615e-08 0 1.47645e-08 0.0007 1.47675e-08 0 1.49415e-08 0 1.49445e-08 0.0007 1.49475e-08 0 1.51215e-08 0 1.51245e-08 0.0007 1.51275e-08 0 1.53015e-08 0 1.53045e-08 0.0007 1.53075e-08 0 1.54815e-08 0 1.54845e-08 0.0007 1.54875e-08 0 1.56615e-08 0 1.56645e-08 0.0007 1.56675e-08 0 1.58415e-08 0 1.58445e-08 0.0007 1.58475e-08 0 1.60215e-08 0 1.60245e-08 0.0007 1.60275e-08 0 1.62015e-08 0 1.62045e-08 0.0007 1.62075e-08 0 1.63815e-08 0 1.63845e-08 0.0007 1.63875e-08 0 1.65615e-08 0 1.65645e-08 0.0007 1.65675e-08 0 1.67415e-08 0 1.67445e-08 0.0007 1.67475e-08 0 1.69215e-08 0 1.69245e-08 0.0007 1.69275e-08 0 1.71015e-08 0 1.71045e-08 0.0007 1.71075e-08 0 1.72815e-08 0 1.72845e-08 0.0007 1.72875e-08 0 1.74615e-08 0 1.74645e-08 0.0007 1.74675e-08 0 1.76415e-08 0 1.76445e-08 0.0007 1.76475e-08 0 1.78215e-08 0 1.78245e-08 0.0007 1.78275e-08 0 1.80015e-08 0 1.80045e-08 0.0007 1.80075e-08 0 1.81815e-08 0 1.81845e-08 0.0007 1.81875e-08 0 1.83615e-08 0 1.83645e-08 0.0007 1.83675e-08 0 1.85415e-08 0 1.85445e-08 0.0007 1.85475e-08 0 1.87215e-08 0 1.87245e-08 0.0007 1.87275e-08 0 1.89015e-08 0 1.89045e-08 0.0007 1.89075e-08 0 1.90815e-08 0 1.90845e-08 0.0007 1.90875e-08 0 1.92615e-08 0 1.92645e-08 0.0007 1.92675e-08 0 1.94415e-08 0 1.94445e-08 0.0007 1.94475e-08 0 1.96215e-08 0 1.96245e-08 0.0007 1.96275e-08 0 1.98015e-08 0 1.98045e-08 0.0007 1.98075e-08 0 1.99815e-08 0 1.99845e-08 0.0007 1.99875e-08 0 2.01615e-08 0 2.01645e-08 0.0007 2.01675e-08 0 2.03415e-08 0 2.03445e-08 0.0007 2.03475e-08 0 2.05215e-08 0 2.05245e-08 0.0007 2.05275e-08 0 2.07015e-08 0 2.07045e-08 0.0007 2.07075e-08 0 2.08815e-08 0 2.08845e-08 0.0007 2.08875e-08 0 2.10615e-08 0 2.10645e-08 0.0007 2.10675e-08 0 2.12415e-08 0 2.12445e-08 0.0007 2.12475e-08 0 2.14215e-08 0 2.14245e-08 0.0007 2.14275e-08 0 2.16015e-08 0 2.16045e-08 0.0007 2.16075e-08 0 2.17815e-08 0 2.17845e-08 0.0007 2.17875e-08 0 2.19615e-08 0 2.19645e-08 0.0007 2.19675e-08 0 2.21415e-08 0 2.21445e-08 0.0007 2.21475e-08 0 2.23215e-08 0 2.23245e-08 0.0007 2.23275e-08 0 2.25015e-08 0 2.25045e-08 0.0007 2.25075e-08 0 2.26815e-08 0 2.26845e-08 0.0007 2.26875e-08 0 2.28615e-08 0 2.28645e-08 0.0007 2.28675e-08 0 2.30415e-08 0 2.30445e-08 0.0007 2.30475e-08 0 2.32215e-08 0 2.32245e-08 0.0007 2.32275e-08 0 2.34015e-08 0 2.34045e-08 0.0007 2.34075e-08 0 2.35815e-08 0 2.35845e-08 0.0007 2.35875e-08 0 2.37615e-08 0 2.37645e-08 0.0007 2.37675e-08 0 2.39415e-08 0 2.39445e-08 0.0007 2.39475e-08 0 2.41215e-08 0 2.41245e-08 0.0007 2.41275e-08 0 2.43015e-08 0 2.43045e-08 0.0007 2.43075e-08 0 2.44815e-08 0 2.44845e-08 0.0007 2.44875e-08 0 2.46615e-08 0 2.46645e-08 0.0007 2.46675e-08 0 2.48415e-08 0 2.48445e-08 0.0007 2.48475e-08 0 2.50215e-08 0 2.50245e-08 0.0007 2.50275e-08 0 2.52015e-08 0 2.52045e-08 0.0007 2.52075e-08 0 2.53815e-08 0 2.53845e-08 0.0007 2.53875e-08 0 2.55615e-08 0 2.55645e-08 0.0007 2.55675e-08 0 2.57415e-08 0 2.57445e-08 0.0007 2.57475e-08 0 2.59215e-08 0 2.59245e-08 0.0007 2.59275e-08 0 2.61015e-08 0 2.61045e-08 0.0007 2.61075e-08 0 2.62815e-08 0 2.62845e-08 0.0007 2.62875e-08 0 2.64615e-08 0 2.64645e-08 0.0007 2.64675e-08 0 2.66415e-08 0 2.66445e-08 0.0007 2.66475e-08 0 2.68215e-08 0 2.68245e-08 0.0007 2.68275e-08 0 2.70015e-08 0 2.70045e-08 0.0007 2.70075e-08 0 2.71815e-08 0 2.71845e-08 0.0007 2.71875e-08 0 2.73615e-08 0 2.73645e-08 0.0007 2.73675e-08 0 2.75415e-08 0 2.75445e-08 0.0007 2.75475e-08 0 2.77215e-08 0 2.77245e-08 0.0007 2.77275e-08 0 2.79015e-08 0 2.79045e-08 0.0007 2.79075e-08 0 2.80815e-08 0 2.80845e-08 0.0007 2.80875e-08 0 2.82615e-08 0 2.82645e-08 0.0007 2.82675e-08 0 2.84415e-08 0 2.84445e-08 0.0007 2.84475e-08 0 2.86215e-08 0 2.86245e-08 0.0007 2.86275e-08 0 2.88015e-08 0 2.88045e-08 0.0007 2.88075e-08 0 2.89815e-08 0 2.89845e-08 0.0007 2.89875e-08 0 2.91615e-08 0 2.91645e-08 0.0007 2.91675e-08 0 2.93415e-08 0 2.93445e-08 0.0007 2.93475e-08 0 2.95215e-08 0 2.95245e-08 0.0007 2.95275e-08 0 2.97015e-08 0 2.97045e-08 0.0007 2.97075e-08 0 2.98815e-08 0 2.98845e-08 0.0007 2.98875e-08 0 3.00615e-08 0 3.00645e-08 0.0007 3.00675e-08 0 3.02415e-08 0 3.02445e-08 0.0007 3.02475e-08 0 3.04215e-08 0 3.04245e-08 0.0007 3.04275e-08 0 3.06015e-08 0 3.06045e-08 0.0007 3.06075e-08 0 3.07815e-08 0 3.07845e-08 0.0007 3.07875e-08 0 3.09615e-08 0 3.09645e-08 0.0007 3.09675e-08 0 3.11415e-08 0 3.11445e-08 0.0007 3.11475e-08 0 3.13215e-08 0 3.13245e-08 0.0007 3.13275e-08 0 3.15015e-08 0 3.15045e-08 0.0007 3.15075e-08 0 3.16815e-08 0 3.16845e-08 0.0007 3.16875e-08 0 3.18615e-08 0 3.18645e-08 0.0007 3.18675e-08 0 3.20415e-08 0 3.20445e-08 0.0007 3.20475e-08 0 3.22215e-08 0 3.22245e-08 0.0007 3.22275e-08 0 3.24015e-08 0 3.24045e-08 0.0007 3.24075e-08 0 3.25815e-08 0 3.25845e-08 0.0007 3.25875e-08 0 3.27615e-08 0 3.27645e-08 0.0007 3.27675e-08 0 3.29415e-08 0 3.29445e-08 0.0007 3.29475e-08 0 3.31215e-08 0 3.31245e-08 0.0007 3.31275e-08 0 3.33015e-08 0 3.33045e-08 0.0007 3.33075e-08 0 3.34815e-08 0 3.34845e-08 0.0007 3.34875e-08 0 3.36615e-08 0 3.36645e-08 0.0007 3.36675e-08 0 3.38415e-08 0 3.38445e-08 0.0007 3.38475e-08 0 3.40215e-08 0 3.40245e-08 0.0007 3.40275e-08 0 3.42015e-08 0 3.42045e-08 0.0007 3.42075e-08 0 3.43815e-08 0 3.43845e-08 0.0007 3.43875e-08 0 3.45615e-08 0 3.45645e-08 0.0007 3.45675e-08 0 3.47415e-08 0 3.47445e-08 0.0007 3.47475e-08 0 3.49215e-08 0 3.49245e-08 0.0007 3.49275e-08 0 3.51015e-08 0 3.51045e-08 0.0007 3.51075e-08 0 3.52815e-08 0 3.52845e-08 0.0007 3.52875e-08 0 3.54615e-08 0 3.54645e-08 0.0007 3.54675e-08 0 3.56415e-08 0 3.56445e-08 0.0007 3.56475e-08 0 3.58215e-08 0 3.58245e-08 0.0007 3.58275e-08 0 3.60015e-08 0 3.60045e-08 0.0007 3.60075e-08 0 3.61815e-08 0 3.61845e-08 0.0007 3.61875e-08 0 3.63615e-08 0 3.63645e-08 0.0007 3.63675e-08 0 3.65415e-08 0 3.65445e-08 0.0007 3.65475e-08 0 3.67215e-08 0 3.67245e-08 0.0007 3.67275e-08 0 3.69015e-08 0 3.69045e-08 0.0007 3.69075e-08 0 3.70815e-08 0 3.70845e-08 0.0007 3.70875e-08 0 3.72615e-08 0 3.72645e-08 0.0007 3.72675e-08 0 3.74415e-08 0 3.74445e-08 0.0007 3.74475e-08 0 3.76215e-08 0 3.76245e-08 0.0007 3.76275e-08 0 3.78015e-08 0 3.78045e-08 0.0007 3.78075e-08 0 3.79815e-08 0 3.79845e-08 0.0007 3.79875e-08 0 3.81615e-08 0 3.81645e-08 0.0007 3.81675e-08 0 3.83415e-08 0 3.83445e-08 0.0007 3.83475e-08 0 3.85215e-08 0 3.85245e-08 0.0007 3.85275e-08 0 3.87015e-08 0 3.87045e-08 0.0007 3.87075e-08 0 3.88815e-08 0 3.88845e-08 0.0007 3.88875e-08 0 3.90615e-08 0 3.90645e-08 0.0007 3.90675e-08 0 3.92415e-08 0 3.92445e-08 0.0007 3.92475e-08 0 3.94215e-08 0 3.94245e-08 0.0007 3.94275e-08 0 3.96015e-08 0 3.96045e-08 0.0007 3.96075e-08 0 3.97815e-08 0 3.97845e-08 0.0007 3.97875e-08 0 3.99615e-08 0 3.99645e-08 0.0007 3.99675e-08 0 4.01415e-08 0 4.01445e-08 0.0007 4.01475e-08 0 4.03215e-08 0 4.03245e-08 0.0007 4.03275e-08 0 4.05015e-08 0 4.05045e-08 0.0007 4.05075e-08 0 4.06815e-08 0 4.06845e-08 0.0007 4.06875e-08 0 4.08615e-08 0 4.08645e-08 0.0007 4.08675e-08 0 4.10415e-08 0 4.10445e-08 0.0007 4.10475e-08 0 4.12215e-08 0 4.12245e-08 0.0007 4.12275e-08 0 4.14015e-08 0 4.14045e-08 0.0007 4.14075e-08 0 4.15815e-08 0 4.15845e-08 0.0007 4.15875e-08 0 4.17615e-08 0 4.17645e-08 0.0007 4.17675e-08 0 4.19415e-08 0 4.19445e-08 0.0007 4.19475e-08 0 4.21215e-08 0 4.21245e-08 0.0007 4.21275e-08 0 4.23015e-08 0 4.23045e-08 0.0007 4.23075e-08 0 4.24815e-08 0 4.24845e-08 0.0007 4.24875e-08 0 4.26615e-08 0 4.26645e-08 0.0007 4.26675e-08 0 4.28415e-08 0 4.28445e-08 0.0007 4.28475e-08 0 4.30215e-08 0 4.30245e-08 0.0007 4.30275e-08 0 4.32015e-08 0 4.32045e-08 0.0007 4.32075e-08 0 4.33815e-08 0 4.33845e-08 0.0007 4.33875e-08 0 4.35615e-08 0 4.35645e-08 0.0007 4.35675e-08 0 4.37415e-08 0 4.37445e-08 0.0007 4.37475e-08 0 4.39215e-08 0 4.39245e-08 0.0007 4.39275e-08 0 4.41015e-08 0 4.41045e-08 0.0007 4.41075e-08 0 4.42815e-08 0 4.42845e-08 0.0007 4.42875e-08 0 4.44615e-08 0 4.44645e-08 0.0007 4.44675e-08 0 4.46415e-08 0 4.46445e-08 0.0007 4.46475e-08 0 4.48215e-08 0 4.48245e-08 0.0007 4.48275e-08 0 4.50015e-08 0 4.50045e-08 0.0007 4.50075e-08 0 4.51815e-08 0 4.51845e-08 0.0007 4.51875e-08 0 4.53615e-08 0 4.53645e-08 0.0007 4.53675e-08 0 4.55415e-08 0 4.55445e-08 0.0007 4.55475e-08 0 4.57215e-08 0 4.57245e-08 0.0007 4.57275e-08 0 4.59015e-08 0 4.59045e-08 0.0007 4.59075e-08 0)
B_S2|1 _S2|1 _S2|2 JJMIT AREA=2.5
B_S2|2 _S2|4 _S2|5 JJMIT AREA=2.09
B_S2|3 _S2|25 _S2|6 JJMIT AREA=1.71
B_S2|4 _S2|9 _S2|10 JJMIT AREA=2.5
B_S2|5 _S2|12 _S2|13 JJMIT AREA=2.09
B_S2|6 _S2|26 _S2|14 JJMIT AREA=1.71
B_S2|7 _S2|27 _S2|16 JJMIT AREA=1.62
B_S2|8 _S2|17 _S2|18 JJMIT AREA=2.5
B_S2|9 _S2|20 _S2|16 JJMIT AREA=1.45
B_S2|10 _S2|16 _S2|21 JJMIT AREA=0.89
B_S2|11 _S2|22 _S2|23 JJMIT AREA=2.5
I_S2|B1 0 _S2|3  PWL(0 0 5e-12 0.000175)
I_S2|B2 0 _S2|7  PWL(0 0 5e-12 0.000112)
I_S2|B3 0 _S2|11  PWL(0 0 5e-12 0.000175)
I_S2|B4 0 _S2|15  PWL(0 0 5e-12 0.000112)
I_S2|B5 0 _S2|19  PWL(0 0 5e-12 0.000175)
I_S2|B6 0 _S2|24  PWL(0 0 5e-12 0.000175)
L_S2|B1 _S2|3 _S2|1  2e-12
L_S2|B2 _S2|7 _S2|6  2e-12
L_S2|B3 _S2|11 _S2|9  2e-12
L_S2|B4 _S2|15 _S2|14  2e-12
L_S2|B5 _S2|19 _S2|17  2e-12
L_S2|B6 _S2|24 _S2|22  2e-12
L_S2|1 G1_2_RX _S2|1  2.06e-12
L_S2|2 _S2|1 _S2|4  3.233e-12
L_S2|3 _S2|4 _S2|25  1.419e-12
L_S2|4 _S2|6 _S2|8  6.051e-12
L_S2|5 IP2_2_OUT_RX _S2|9  2.092e-12
L_S2|6 _S2|9 _S2|12  3.221e-12
L_S2|7 _S2|12 _S2|26  1.384e-12
L_S2|8 _S2|14 _S2|8  6.059e-12
L_S2|9 _S2|8 _S2|27  1.301e-12
L_S2|10 T14 _S2|17  2.082e-12
L_S2|11 _S2|17 _S2|20  1.43e-12
L_S2|12 _S2|16 _S2|22  3.892e-12
L_S2|13 _S2|22 S2  2.077e-12
L_S2|P1 _S2|2 0  5.508e-13
L_S2|P2 _S2|5 0  4.769e-13
L_S2|P4 _S2|10 0  4.767e-13
L_S2|P5 _S2|13 0  4.812e-13
L_S2|P8 _S2|18 0  4.526e-13
L_S2|P10 _S2|21 0  5.69e-13
L_S2|P11 _S2|23 0  4.746e-13
R_S2|B1 _S2|1 _S2|101  2.7439617672
L_S2|RB1 _S2|101 0  2.050338398468e-12
R_S2|B2 _S2|4 _S2|104  3.2822509177033496
L_S2|RB2 _S2|104 0  2.3544717685023925e-12
R_S2|B3 _S2|4 _S2|106  4.011640010526316
L_S2|RB3 _S2|106 _S2|6  2.766576605947368e-12
R_S2|B4 _S2|9 _S2|109  2.7439617672
L_S2|RB4 _S2|109 0  2.050338398468e-12
R_S2|B5 _S2|12 _S2|112  3.2822509177033496
L_S2|RB5 _S2|112 0  2.3544717685023925e-12
R_S2|B6 _S2|12 _S2|114  4.011640010526316
L_S2|RB6 _S2|114 _S2|14  2.766576605947368e-12
R_S2|B7 _S2|8 _S2|108  4.2345089
L_S2|RB7 _S2|108 _S2|16  2.8924975284999997e-12
R_S2|B8 _S2|17 _S2|117  2.7439617672
L_S2|RB8 _S2|117 0  2.050338398468e-12
R_S2|B9 _S2|20 _S2|120  4.730968564137931
L_S2|RB9 _S2|120 _S2|16  3.172997238737931e-12
R_S2|B10 _S2|16 _S2|116  7.707757773033708
L_S2|RB10 _S2|116 0  4.854883141764045e-12
R_S2|B11 _S2|22 _S2|122  2.7439617672
L_S2|RB11 _S2|122 0  2.050338398468e-12
IT15|T 0 T15  PWL(0 0 1.5e-12 0 4.5e-12 0.0007 7.5e-12 0 1.815e-10 0 1.845e-10 0.0007 1.875e-10 0 3.615e-10 0 3.645e-10 0.0007 3.675e-10 0 5.415e-10 0 5.445e-10 0.0007 5.475e-10 0 7.215e-10 0 7.245e-10 0.0007 7.275e-10 0 9.015e-10 0 9.045e-10 0.0007 9.075e-10 0 1.0815e-09 0 1.0845e-09 0.0007 1.0875e-09 0 1.2615e-09 0 1.2645e-09 0.0007 1.2675e-09 0 1.4415e-09 0 1.4445e-09 0.0007 1.4475e-09 0 1.6215e-09 0 1.6245e-09 0.0007 1.6275e-09 0 1.8015e-09 0 1.8045e-09 0.0007 1.8075e-09 0 1.9815e-09 0 1.9845e-09 0.0007 1.9875e-09 0 2.1615e-09 0 2.1645e-09 0.0007 2.1675e-09 0 2.3415e-09 0 2.3445e-09 0.0007 2.3475e-09 0 2.5215e-09 0 2.5245e-09 0.0007 2.5275e-09 0 2.7015e-09 0 2.7045e-09 0.0007 2.7075e-09 0 2.8815e-09 0 2.8845e-09 0.0007 2.8875e-09 0 3.0615e-09 0 3.0645e-09 0.0007 3.0675e-09 0 3.2415e-09 0 3.2445e-09 0.0007 3.2475e-09 0 3.4215e-09 0 3.4245e-09 0.0007 3.4275e-09 0 3.6015e-09 0 3.6045e-09 0.0007 3.6075e-09 0 3.7815e-09 0 3.7845e-09 0.0007 3.7875e-09 0 3.9615e-09 0 3.9645e-09 0.0007 3.9675e-09 0 4.1415e-09 0 4.1445e-09 0.0007 4.1475e-09 0 4.3215e-09 0 4.3245e-09 0.0007 4.3275e-09 0 4.5015e-09 0 4.5045e-09 0.0007 4.5075e-09 0 4.6815e-09 0 4.6845e-09 0.0007 4.6875e-09 0 4.8615e-09 0 4.8645e-09 0.0007 4.8675e-09 0 5.0415e-09 0 5.0445e-09 0.0007 5.0475e-09 0 5.2215e-09 0 5.2245e-09 0.0007 5.2275e-09 0 5.4015e-09 0 5.4045e-09 0.0007 5.4075e-09 0 5.5815e-09 0 5.5845e-09 0.0007 5.5875e-09 0 5.7615e-09 0 5.7645e-09 0.0007 5.7675e-09 0 5.9415e-09 0 5.9445e-09 0.0007 5.9475e-09 0 6.1215e-09 0 6.1245e-09 0.0007 6.1275e-09 0 6.3015e-09 0 6.3045e-09 0.0007 6.3075e-09 0 6.4815e-09 0 6.4845e-09 0.0007 6.4875e-09 0 6.6615e-09 0 6.6645e-09 0.0007 6.6675e-09 0 6.8415e-09 0 6.8445e-09 0.0007 6.8475e-09 0 7.0215e-09 0 7.0245e-09 0.0007 7.0275e-09 0 7.2015e-09 0 7.2045e-09 0.0007 7.2075e-09 0 7.3815e-09 0 7.3845e-09 0.0007 7.3875e-09 0 7.5615e-09 0 7.5645e-09 0.0007 7.5675e-09 0 7.7415e-09 0 7.7445e-09 0.0007 7.7475e-09 0 7.9215e-09 0 7.9245e-09 0.0007 7.9275e-09 0 8.1015e-09 0 8.1045e-09 0.0007 8.1075e-09 0 8.2815e-09 0 8.2845e-09 0.0007 8.2875e-09 0 8.4615e-09 0 8.4645e-09 0.0007 8.4675e-09 0 8.6415e-09 0 8.6445e-09 0.0007 8.6475e-09 0 8.8215e-09 0 8.8245e-09 0.0007 8.8275e-09 0 9.0015e-09 0 9.0045e-09 0.0007 9.0075e-09 0 9.1815e-09 0 9.1845e-09 0.0007 9.1875e-09 0 9.3615e-09 0 9.3645e-09 0.0007 9.3675e-09 0 9.5415e-09 0 9.5445e-09 0.0007 9.5475e-09 0 9.7215e-09 0 9.7245e-09 0.0007 9.7275e-09 0 9.9015e-09 0 9.9045e-09 0.0007 9.9075e-09 0 1.00815e-08 0 1.00845e-08 0.0007 1.00875e-08 0 1.02615e-08 0 1.02645e-08 0.0007 1.02675e-08 0 1.04415e-08 0 1.04445e-08 0.0007 1.04475e-08 0 1.06215e-08 0 1.06245e-08 0.0007 1.06275e-08 0 1.08015e-08 0 1.08045e-08 0.0007 1.08075e-08 0 1.09815e-08 0 1.09845e-08 0.0007 1.09875e-08 0 1.11615e-08 0 1.11645e-08 0.0007 1.11675e-08 0 1.13415e-08 0 1.13445e-08 0.0007 1.13475e-08 0 1.15215e-08 0 1.15245e-08 0.0007 1.15275e-08 0 1.17015e-08 0 1.17045e-08 0.0007 1.17075e-08 0 1.18815e-08 0 1.18845e-08 0.0007 1.18875e-08 0 1.20615e-08 0 1.20645e-08 0.0007 1.20675e-08 0 1.22415e-08 0 1.22445e-08 0.0007 1.22475e-08 0 1.24215e-08 0 1.24245e-08 0.0007 1.24275e-08 0 1.26015e-08 0 1.26045e-08 0.0007 1.26075e-08 0 1.27815e-08 0 1.27845e-08 0.0007 1.27875e-08 0 1.29615e-08 0 1.29645e-08 0.0007 1.29675e-08 0 1.31415e-08 0 1.31445e-08 0.0007 1.31475e-08 0 1.33215e-08 0 1.33245e-08 0.0007 1.33275e-08 0 1.35015e-08 0 1.35045e-08 0.0007 1.35075e-08 0 1.36815e-08 0 1.36845e-08 0.0007 1.36875e-08 0 1.38615e-08 0 1.38645e-08 0.0007 1.38675e-08 0 1.40415e-08 0 1.40445e-08 0.0007 1.40475e-08 0 1.42215e-08 0 1.42245e-08 0.0007 1.42275e-08 0 1.44015e-08 0 1.44045e-08 0.0007 1.44075e-08 0 1.45815e-08 0 1.45845e-08 0.0007 1.45875e-08 0 1.47615e-08 0 1.47645e-08 0.0007 1.47675e-08 0 1.49415e-08 0 1.49445e-08 0.0007 1.49475e-08 0 1.51215e-08 0 1.51245e-08 0.0007 1.51275e-08 0 1.53015e-08 0 1.53045e-08 0.0007 1.53075e-08 0 1.54815e-08 0 1.54845e-08 0.0007 1.54875e-08 0 1.56615e-08 0 1.56645e-08 0.0007 1.56675e-08 0 1.58415e-08 0 1.58445e-08 0.0007 1.58475e-08 0 1.60215e-08 0 1.60245e-08 0.0007 1.60275e-08 0 1.62015e-08 0 1.62045e-08 0.0007 1.62075e-08 0 1.63815e-08 0 1.63845e-08 0.0007 1.63875e-08 0 1.65615e-08 0 1.65645e-08 0.0007 1.65675e-08 0 1.67415e-08 0 1.67445e-08 0.0007 1.67475e-08 0 1.69215e-08 0 1.69245e-08 0.0007 1.69275e-08 0 1.71015e-08 0 1.71045e-08 0.0007 1.71075e-08 0 1.72815e-08 0 1.72845e-08 0.0007 1.72875e-08 0 1.74615e-08 0 1.74645e-08 0.0007 1.74675e-08 0 1.76415e-08 0 1.76445e-08 0.0007 1.76475e-08 0 1.78215e-08 0 1.78245e-08 0.0007 1.78275e-08 0 1.80015e-08 0 1.80045e-08 0.0007 1.80075e-08 0 1.81815e-08 0 1.81845e-08 0.0007 1.81875e-08 0 1.83615e-08 0 1.83645e-08 0.0007 1.83675e-08 0 1.85415e-08 0 1.85445e-08 0.0007 1.85475e-08 0 1.87215e-08 0 1.87245e-08 0.0007 1.87275e-08 0 1.89015e-08 0 1.89045e-08 0.0007 1.89075e-08 0 1.90815e-08 0 1.90845e-08 0.0007 1.90875e-08 0 1.92615e-08 0 1.92645e-08 0.0007 1.92675e-08 0 1.94415e-08 0 1.94445e-08 0.0007 1.94475e-08 0 1.96215e-08 0 1.96245e-08 0.0007 1.96275e-08 0 1.98015e-08 0 1.98045e-08 0.0007 1.98075e-08 0 1.99815e-08 0 1.99845e-08 0.0007 1.99875e-08 0 2.01615e-08 0 2.01645e-08 0.0007 2.01675e-08 0 2.03415e-08 0 2.03445e-08 0.0007 2.03475e-08 0 2.05215e-08 0 2.05245e-08 0.0007 2.05275e-08 0 2.07015e-08 0 2.07045e-08 0.0007 2.07075e-08 0 2.08815e-08 0 2.08845e-08 0.0007 2.08875e-08 0 2.10615e-08 0 2.10645e-08 0.0007 2.10675e-08 0 2.12415e-08 0 2.12445e-08 0.0007 2.12475e-08 0 2.14215e-08 0 2.14245e-08 0.0007 2.14275e-08 0 2.16015e-08 0 2.16045e-08 0.0007 2.16075e-08 0 2.17815e-08 0 2.17845e-08 0.0007 2.17875e-08 0 2.19615e-08 0 2.19645e-08 0.0007 2.19675e-08 0 2.21415e-08 0 2.21445e-08 0.0007 2.21475e-08 0 2.23215e-08 0 2.23245e-08 0.0007 2.23275e-08 0 2.25015e-08 0 2.25045e-08 0.0007 2.25075e-08 0 2.26815e-08 0 2.26845e-08 0.0007 2.26875e-08 0 2.28615e-08 0 2.28645e-08 0.0007 2.28675e-08 0 2.30415e-08 0 2.30445e-08 0.0007 2.30475e-08 0 2.32215e-08 0 2.32245e-08 0.0007 2.32275e-08 0 2.34015e-08 0 2.34045e-08 0.0007 2.34075e-08 0 2.35815e-08 0 2.35845e-08 0.0007 2.35875e-08 0 2.37615e-08 0 2.37645e-08 0.0007 2.37675e-08 0 2.39415e-08 0 2.39445e-08 0.0007 2.39475e-08 0 2.41215e-08 0 2.41245e-08 0.0007 2.41275e-08 0 2.43015e-08 0 2.43045e-08 0.0007 2.43075e-08 0 2.44815e-08 0 2.44845e-08 0.0007 2.44875e-08 0 2.46615e-08 0 2.46645e-08 0.0007 2.46675e-08 0 2.48415e-08 0 2.48445e-08 0.0007 2.48475e-08 0 2.50215e-08 0 2.50245e-08 0.0007 2.50275e-08 0 2.52015e-08 0 2.52045e-08 0.0007 2.52075e-08 0 2.53815e-08 0 2.53845e-08 0.0007 2.53875e-08 0 2.55615e-08 0 2.55645e-08 0.0007 2.55675e-08 0 2.57415e-08 0 2.57445e-08 0.0007 2.57475e-08 0 2.59215e-08 0 2.59245e-08 0.0007 2.59275e-08 0 2.61015e-08 0 2.61045e-08 0.0007 2.61075e-08 0 2.62815e-08 0 2.62845e-08 0.0007 2.62875e-08 0 2.64615e-08 0 2.64645e-08 0.0007 2.64675e-08 0 2.66415e-08 0 2.66445e-08 0.0007 2.66475e-08 0 2.68215e-08 0 2.68245e-08 0.0007 2.68275e-08 0 2.70015e-08 0 2.70045e-08 0.0007 2.70075e-08 0 2.71815e-08 0 2.71845e-08 0.0007 2.71875e-08 0 2.73615e-08 0 2.73645e-08 0.0007 2.73675e-08 0 2.75415e-08 0 2.75445e-08 0.0007 2.75475e-08 0 2.77215e-08 0 2.77245e-08 0.0007 2.77275e-08 0 2.79015e-08 0 2.79045e-08 0.0007 2.79075e-08 0 2.80815e-08 0 2.80845e-08 0.0007 2.80875e-08 0 2.82615e-08 0 2.82645e-08 0.0007 2.82675e-08 0 2.84415e-08 0 2.84445e-08 0.0007 2.84475e-08 0 2.86215e-08 0 2.86245e-08 0.0007 2.86275e-08 0 2.88015e-08 0 2.88045e-08 0.0007 2.88075e-08 0 2.89815e-08 0 2.89845e-08 0.0007 2.89875e-08 0 2.91615e-08 0 2.91645e-08 0.0007 2.91675e-08 0 2.93415e-08 0 2.93445e-08 0.0007 2.93475e-08 0 2.95215e-08 0 2.95245e-08 0.0007 2.95275e-08 0 2.97015e-08 0 2.97045e-08 0.0007 2.97075e-08 0 2.98815e-08 0 2.98845e-08 0.0007 2.98875e-08 0 3.00615e-08 0 3.00645e-08 0.0007 3.00675e-08 0 3.02415e-08 0 3.02445e-08 0.0007 3.02475e-08 0 3.04215e-08 0 3.04245e-08 0.0007 3.04275e-08 0 3.06015e-08 0 3.06045e-08 0.0007 3.06075e-08 0 3.07815e-08 0 3.07845e-08 0.0007 3.07875e-08 0 3.09615e-08 0 3.09645e-08 0.0007 3.09675e-08 0 3.11415e-08 0 3.11445e-08 0.0007 3.11475e-08 0 3.13215e-08 0 3.13245e-08 0.0007 3.13275e-08 0 3.15015e-08 0 3.15045e-08 0.0007 3.15075e-08 0 3.16815e-08 0 3.16845e-08 0.0007 3.16875e-08 0 3.18615e-08 0 3.18645e-08 0.0007 3.18675e-08 0 3.20415e-08 0 3.20445e-08 0.0007 3.20475e-08 0 3.22215e-08 0 3.22245e-08 0.0007 3.22275e-08 0 3.24015e-08 0 3.24045e-08 0.0007 3.24075e-08 0 3.25815e-08 0 3.25845e-08 0.0007 3.25875e-08 0 3.27615e-08 0 3.27645e-08 0.0007 3.27675e-08 0 3.29415e-08 0 3.29445e-08 0.0007 3.29475e-08 0 3.31215e-08 0 3.31245e-08 0.0007 3.31275e-08 0 3.33015e-08 0 3.33045e-08 0.0007 3.33075e-08 0 3.34815e-08 0 3.34845e-08 0.0007 3.34875e-08 0 3.36615e-08 0 3.36645e-08 0.0007 3.36675e-08 0 3.38415e-08 0 3.38445e-08 0.0007 3.38475e-08 0 3.40215e-08 0 3.40245e-08 0.0007 3.40275e-08 0 3.42015e-08 0 3.42045e-08 0.0007 3.42075e-08 0 3.43815e-08 0 3.43845e-08 0.0007 3.43875e-08 0 3.45615e-08 0 3.45645e-08 0.0007 3.45675e-08 0 3.47415e-08 0 3.47445e-08 0.0007 3.47475e-08 0 3.49215e-08 0 3.49245e-08 0.0007 3.49275e-08 0 3.51015e-08 0 3.51045e-08 0.0007 3.51075e-08 0 3.52815e-08 0 3.52845e-08 0.0007 3.52875e-08 0 3.54615e-08 0 3.54645e-08 0.0007 3.54675e-08 0 3.56415e-08 0 3.56445e-08 0.0007 3.56475e-08 0 3.58215e-08 0 3.58245e-08 0.0007 3.58275e-08 0 3.60015e-08 0 3.60045e-08 0.0007 3.60075e-08 0 3.61815e-08 0 3.61845e-08 0.0007 3.61875e-08 0 3.63615e-08 0 3.63645e-08 0.0007 3.63675e-08 0 3.65415e-08 0 3.65445e-08 0.0007 3.65475e-08 0 3.67215e-08 0 3.67245e-08 0.0007 3.67275e-08 0 3.69015e-08 0 3.69045e-08 0.0007 3.69075e-08 0 3.70815e-08 0 3.70845e-08 0.0007 3.70875e-08 0 3.72615e-08 0 3.72645e-08 0.0007 3.72675e-08 0 3.74415e-08 0 3.74445e-08 0.0007 3.74475e-08 0 3.76215e-08 0 3.76245e-08 0.0007 3.76275e-08 0 3.78015e-08 0 3.78045e-08 0.0007 3.78075e-08 0 3.79815e-08 0 3.79845e-08 0.0007 3.79875e-08 0 3.81615e-08 0 3.81645e-08 0.0007 3.81675e-08 0 3.83415e-08 0 3.83445e-08 0.0007 3.83475e-08 0 3.85215e-08 0 3.85245e-08 0.0007 3.85275e-08 0 3.87015e-08 0 3.87045e-08 0.0007 3.87075e-08 0 3.88815e-08 0 3.88845e-08 0.0007 3.88875e-08 0 3.90615e-08 0 3.90645e-08 0.0007 3.90675e-08 0 3.92415e-08 0 3.92445e-08 0.0007 3.92475e-08 0 3.94215e-08 0 3.94245e-08 0.0007 3.94275e-08 0 3.96015e-08 0 3.96045e-08 0.0007 3.96075e-08 0 3.97815e-08 0 3.97845e-08 0.0007 3.97875e-08 0 3.99615e-08 0 3.99645e-08 0.0007 3.99675e-08 0 4.01415e-08 0 4.01445e-08 0.0007 4.01475e-08 0 4.03215e-08 0 4.03245e-08 0.0007 4.03275e-08 0 4.05015e-08 0 4.05045e-08 0.0007 4.05075e-08 0 4.06815e-08 0 4.06845e-08 0.0007 4.06875e-08 0 4.08615e-08 0 4.08645e-08 0.0007 4.08675e-08 0 4.10415e-08 0 4.10445e-08 0.0007 4.10475e-08 0 4.12215e-08 0 4.12245e-08 0.0007 4.12275e-08 0 4.14015e-08 0 4.14045e-08 0.0007 4.14075e-08 0 4.15815e-08 0 4.15845e-08 0.0007 4.15875e-08 0 4.17615e-08 0 4.17645e-08 0.0007 4.17675e-08 0 4.19415e-08 0 4.19445e-08 0.0007 4.19475e-08 0 4.21215e-08 0 4.21245e-08 0.0007 4.21275e-08 0 4.23015e-08 0 4.23045e-08 0.0007 4.23075e-08 0 4.24815e-08 0 4.24845e-08 0.0007 4.24875e-08 0 4.26615e-08 0 4.26645e-08 0.0007 4.26675e-08 0 4.28415e-08 0 4.28445e-08 0.0007 4.28475e-08 0 4.30215e-08 0 4.30245e-08 0.0007 4.30275e-08 0 4.32015e-08 0 4.32045e-08 0.0007 4.32075e-08 0 4.33815e-08 0 4.33845e-08 0.0007 4.33875e-08 0 4.35615e-08 0 4.35645e-08 0.0007 4.35675e-08 0 4.37415e-08 0 4.37445e-08 0.0007 4.37475e-08 0 4.39215e-08 0 4.39245e-08 0.0007 4.39275e-08 0 4.41015e-08 0 4.41045e-08 0.0007 4.41075e-08 0 4.42815e-08 0 4.42845e-08 0.0007 4.42875e-08 0 4.44615e-08 0 4.44645e-08 0.0007 4.44675e-08 0 4.46415e-08 0 4.46445e-08 0.0007 4.46475e-08 0 4.48215e-08 0 4.48245e-08 0.0007 4.48275e-08 0 4.50015e-08 0 4.50045e-08 0.0007 4.50075e-08 0 4.51815e-08 0 4.51845e-08 0.0007 4.51875e-08 0 4.53615e-08 0 4.53645e-08 0.0007 4.53675e-08 0 4.55415e-08 0 4.55445e-08 0.0007 4.55475e-08 0 4.57215e-08 0 4.57245e-08 0.0007 4.57275e-08 0 4.59015e-08 0 4.59045e-08 0.0007 4.59075e-08 0)
B_S3|1 _S3|1 _S3|2 JJMIT AREA=2.5
B_S3|2 _S3|4 _S3|5 JJMIT AREA=2.09
B_S3|3 _S3|25 _S3|6 JJMIT AREA=1.71
B_S3|4 _S3|9 _S3|10 JJMIT AREA=2.5
B_S3|5 _S3|12 _S3|13 JJMIT AREA=2.09
B_S3|6 _S3|26 _S3|14 JJMIT AREA=1.71
B_S3|7 _S3|27 _S3|16 JJMIT AREA=1.62
B_S3|8 _S3|17 _S3|18 JJMIT AREA=2.5
B_S3|9 _S3|20 _S3|16 JJMIT AREA=1.45
B_S3|10 _S3|16 _S3|21 JJMIT AREA=0.89
B_S3|11 _S3|22 _S3|23 JJMIT AREA=2.5
I_S3|B1 0 _S3|3  PWL(0 0 5e-12 0.000175)
I_S3|B2 0 _S3|7  PWL(0 0 5e-12 0.000112)
I_S3|B3 0 _S3|11  PWL(0 0 5e-12 0.000175)
I_S3|B4 0 _S3|15  PWL(0 0 5e-12 0.000112)
I_S3|B5 0 _S3|19  PWL(0 0 5e-12 0.000175)
I_S3|B6 0 _S3|24  PWL(0 0 5e-12 0.000175)
L_S3|B1 _S3|3 _S3|1  2e-12
L_S3|B2 _S3|7 _S3|6  2e-12
L_S3|B3 _S3|11 _S3|9  2e-12
L_S3|B4 _S3|15 _S3|14  2e-12
L_S3|B5 _S3|19 _S3|17  2e-12
L_S3|B6 _S3|24 _S3|22  2e-12
L_S3|1 G2_2_RX _S3|1  2.06e-12
L_S3|2 _S3|1 _S3|4  3.233e-12
L_S3|3 _S3|4 _S3|25  1.419e-12
L_S3|4 _S3|6 _S3|8  6.051e-12
L_S3|5 IP3_2_OUT_RX _S3|9  2.092e-12
L_S3|6 _S3|9 _S3|12  3.221e-12
L_S3|7 _S3|12 _S3|26  1.384e-12
L_S3|8 _S3|14 _S3|8  6.059e-12
L_S3|9 _S3|8 _S3|27  1.301e-12
L_S3|10 T15 _S3|17  2.082e-12
L_S3|11 _S3|17 _S3|20  1.43e-12
L_S3|12 _S3|16 _S3|22  3.892e-12
L_S3|13 _S3|22 S3  2.077e-12
L_S3|P1 _S3|2 0  5.508e-13
L_S3|P2 _S3|5 0  4.769e-13
L_S3|P4 _S3|10 0  4.767e-13
L_S3|P5 _S3|13 0  4.812e-13
L_S3|P8 _S3|18 0  4.526e-13
L_S3|P10 _S3|21 0  5.69e-13
L_S3|P11 _S3|23 0  4.746e-13
R_S3|B1 _S3|1 _S3|101  2.7439617672
L_S3|RB1 _S3|101 0  2.050338398468e-12
R_S3|B2 _S3|4 _S3|104  3.2822509177033496
L_S3|RB2 _S3|104 0  2.3544717685023925e-12
R_S3|B3 _S3|4 _S3|106  4.011640010526316
L_S3|RB3 _S3|106 _S3|6  2.766576605947368e-12
R_S3|B4 _S3|9 _S3|109  2.7439617672
L_S3|RB4 _S3|109 0  2.050338398468e-12
R_S3|B5 _S3|12 _S3|112  3.2822509177033496
L_S3|RB5 _S3|112 0  2.3544717685023925e-12
R_S3|B6 _S3|12 _S3|114  4.011640010526316
L_S3|RB6 _S3|114 _S3|14  2.766576605947368e-12
R_S3|B7 _S3|8 _S3|108  4.2345089
L_S3|RB7 _S3|108 _S3|16  2.8924975284999997e-12
R_S3|B8 _S3|17 _S3|117  2.7439617672
L_S3|RB8 _S3|117 0  2.050338398468e-12
R_S3|B9 _S3|20 _S3|120  4.730968564137931
L_S3|RB9 _S3|120 _S3|16  3.172997238737931e-12
R_S3|B10 _S3|16 _S3|116  7.707757773033708
L_S3|RB10 _S3|116 0  4.854883141764045e-12
R_S3|B11 _S3|22 _S3|122  2.7439617672
L_S3|RB11 _S3|122 0  2.050338398468e-12
IT16|T 0 T16  PWL(0 0 1.5e-12 0 4.5e-12 0.0007 7.5e-12 0 1.815e-10 0 1.845e-10 0.0007 1.875e-10 0 3.615e-10 0 3.645e-10 0.0007 3.675e-10 0 5.415e-10 0 5.445e-10 0.0007 5.475e-10 0 7.215e-10 0 7.245e-10 0.0007 7.275e-10 0 9.015e-10 0 9.045e-10 0.0007 9.075e-10 0 1.0815e-09 0 1.0845e-09 0.0007 1.0875e-09 0 1.2615e-09 0 1.2645e-09 0.0007 1.2675e-09 0 1.4415e-09 0 1.4445e-09 0.0007 1.4475e-09 0 1.6215e-09 0 1.6245e-09 0.0007 1.6275e-09 0 1.8015e-09 0 1.8045e-09 0.0007 1.8075e-09 0 1.9815e-09 0 1.9845e-09 0.0007 1.9875e-09 0 2.1615e-09 0 2.1645e-09 0.0007 2.1675e-09 0 2.3415e-09 0 2.3445e-09 0.0007 2.3475e-09 0 2.5215e-09 0 2.5245e-09 0.0007 2.5275e-09 0 2.7015e-09 0 2.7045e-09 0.0007 2.7075e-09 0 2.8815e-09 0 2.8845e-09 0.0007 2.8875e-09 0 3.0615e-09 0 3.0645e-09 0.0007 3.0675e-09 0 3.2415e-09 0 3.2445e-09 0.0007 3.2475e-09 0 3.4215e-09 0 3.4245e-09 0.0007 3.4275e-09 0 3.6015e-09 0 3.6045e-09 0.0007 3.6075e-09 0 3.7815e-09 0 3.7845e-09 0.0007 3.7875e-09 0 3.9615e-09 0 3.9645e-09 0.0007 3.9675e-09 0 4.1415e-09 0 4.1445e-09 0.0007 4.1475e-09 0 4.3215e-09 0 4.3245e-09 0.0007 4.3275e-09 0 4.5015e-09 0 4.5045e-09 0.0007 4.5075e-09 0 4.6815e-09 0 4.6845e-09 0.0007 4.6875e-09 0 4.8615e-09 0 4.8645e-09 0.0007 4.8675e-09 0 5.0415e-09 0 5.0445e-09 0.0007 5.0475e-09 0 5.2215e-09 0 5.2245e-09 0.0007 5.2275e-09 0 5.4015e-09 0 5.4045e-09 0.0007 5.4075e-09 0 5.5815e-09 0 5.5845e-09 0.0007 5.5875e-09 0 5.7615e-09 0 5.7645e-09 0.0007 5.7675e-09 0 5.9415e-09 0 5.9445e-09 0.0007 5.9475e-09 0 6.1215e-09 0 6.1245e-09 0.0007 6.1275e-09 0 6.3015e-09 0 6.3045e-09 0.0007 6.3075e-09 0 6.4815e-09 0 6.4845e-09 0.0007 6.4875e-09 0 6.6615e-09 0 6.6645e-09 0.0007 6.6675e-09 0 6.8415e-09 0 6.8445e-09 0.0007 6.8475e-09 0 7.0215e-09 0 7.0245e-09 0.0007 7.0275e-09 0 7.2015e-09 0 7.2045e-09 0.0007 7.2075e-09 0 7.3815e-09 0 7.3845e-09 0.0007 7.3875e-09 0 7.5615e-09 0 7.5645e-09 0.0007 7.5675e-09 0 7.7415e-09 0 7.7445e-09 0.0007 7.7475e-09 0 7.9215e-09 0 7.9245e-09 0.0007 7.9275e-09 0 8.1015e-09 0 8.1045e-09 0.0007 8.1075e-09 0 8.2815e-09 0 8.2845e-09 0.0007 8.2875e-09 0 8.4615e-09 0 8.4645e-09 0.0007 8.4675e-09 0 8.6415e-09 0 8.6445e-09 0.0007 8.6475e-09 0 8.8215e-09 0 8.8245e-09 0.0007 8.8275e-09 0 9.0015e-09 0 9.0045e-09 0.0007 9.0075e-09 0 9.1815e-09 0 9.1845e-09 0.0007 9.1875e-09 0 9.3615e-09 0 9.3645e-09 0.0007 9.3675e-09 0 9.5415e-09 0 9.5445e-09 0.0007 9.5475e-09 0 9.7215e-09 0 9.7245e-09 0.0007 9.7275e-09 0 9.9015e-09 0 9.9045e-09 0.0007 9.9075e-09 0 1.00815e-08 0 1.00845e-08 0.0007 1.00875e-08 0 1.02615e-08 0 1.02645e-08 0.0007 1.02675e-08 0 1.04415e-08 0 1.04445e-08 0.0007 1.04475e-08 0 1.06215e-08 0 1.06245e-08 0.0007 1.06275e-08 0 1.08015e-08 0 1.08045e-08 0.0007 1.08075e-08 0 1.09815e-08 0 1.09845e-08 0.0007 1.09875e-08 0 1.11615e-08 0 1.11645e-08 0.0007 1.11675e-08 0 1.13415e-08 0 1.13445e-08 0.0007 1.13475e-08 0 1.15215e-08 0 1.15245e-08 0.0007 1.15275e-08 0 1.17015e-08 0 1.17045e-08 0.0007 1.17075e-08 0 1.18815e-08 0 1.18845e-08 0.0007 1.18875e-08 0 1.20615e-08 0 1.20645e-08 0.0007 1.20675e-08 0 1.22415e-08 0 1.22445e-08 0.0007 1.22475e-08 0 1.24215e-08 0 1.24245e-08 0.0007 1.24275e-08 0 1.26015e-08 0 1.26045e-08 0.0007 1.26075e-08 0 1.27815e-08 0 1.27845e-08 0.0007 1.27875e-08 0 1.29615e-08 0 1.29645e-08 0.0007 1.29675e-08 0 1.31415e-08 0 1.31445e-08 0.0007 1.31475e-08 0 1.33215e-08 0 1.33245e-08 0.0007 1.33275e-08 0 1.35015e-08 0 1.35045e-08 0.0007 1.35075e-08 0 1.36815e-08 0 1.36845e-08 0.0007 1.36875e-08 0 1.38615e-08 0 1.38645e-08 0.0007 1.38675e-08 0 1.40415e-08 0 1.40445e-08 0.0007 1.40475e-08 0 1.42215e-08 0 1.42245e-08 0.0007 1.42275e-08 0 1.44015e-08 0 1.44045e-08 0.0007 1.44075e-08 0 1.45815e-08 0 1.45845e-08 0.0007 1.45875e-08 0 1.47615e-08 0 1.47645e-08 0.0007 1.47675e-08 0 1.49415e-08 0 1.49445e-08 0.0007 1.49475e-08 0 1.51215e-08 0 1.51245e-08 0.0007 1.51275e-08 0 1.53015e-08 0 1.53045e-08 0.0007 1.53075e-08 0 1.54815e-08 0 1.54845e-08 0.0007 1.54875e-08 0 1.56615e-08 0 1.56645e-08 0.0007 1.56675e-08 0 1.58415e-08 0 1.58445e-08 0.0007 1.58475e-08 0 1.60215e-08 0 1.60245e-08 0.0007 1.60275e-08 0 1.62015e-08 0 1.62045e-08 0.0007 1.62075e-08 0 1.63815e-08 0 1.63845e-08 0.0007 1.63875e-08 0 1.65615e-08 0 1.65645e-08 0.0007 1.65675e-08 0 1.67415e-08 0 1.67445e-08 0.0007 1.67475e-08 0 1.69215e-08 0 1.69245e-08 0.0007 1.69275e-08 0 1.71015e-08 0 1.71045e-08 0.0007 1.71075e-08 0 1.72815e-08 0 1.72845e-08 0.0007 1.72875e-08 0 1.74615e-08 0 1.74645e-08 0.0007 1.74675e-08 0 1.76415e-08 0 1.76445e-08 0.0007 1.76475e-08 0 1.78215e-08 0 1.78245e-08 0.0007 1.78275e-08 0 1.80015e-08 0 1.80045e-08 0.0007 1.80075e-08 0 1.81815e-08 0 1.81845e-08 0.0007 1.81875e-08 0 1.83615e-08 0 1.83645e-08 0.0007 1.83675e-08 0 1.85415e-08 0 1.85445e-08 0.0007 1.85475e-08 0 1.87215e-08 0 1.87245e-08 0.0007 1.87275e-08 0 1.89015e-08 0 1.89045e-08 0.0007 1.89075e-08 0 1.90815e-08 0 1.90845e-08 0.0007 1.90875e-08 0 1.92615e-08 0 1.92645e-08 0.0007 1.92675e-08 0 1.94415e-08 0 1.94445e-08 0.0007 1.94475e-08 0 1.96215e-08 0 1.96245e-08 0.0007 1.96275e-08 0 1.98015e-08 0 1.98045e-08 0.0007 1.98075e-08 0 1.99815e-08 0 1.99845e-08 0.0007 1.99875e-08 0 2.01615e-08 0 2.01645e-08 0.0007 2.01675e-08 0 2.03415e-08 0 2.03445e-08 0.0007 2.03475e-08 0 2.05215e-08 0 2.05245e-08 0.0007 2.05275e-08 0 2.07015e-08 0 2.07045e-08 0.0007 2.07075e-08 0 2.08815e-08 0 2.08845e-08 0.0007 2.08875e-08 0 2.10615e-08 0 2.10645e-08 0.0007 2.10675e-08 0 2.12415e-08 0 2.12445e-08 0.0007 2.12475e-08 0 2.14215e-08 0 2.14245e-08 0.0007 2.14275e-08 0 2.16015e-08 0 2.16045e-08 0.0007 2.16075e-08 0 2.17815e-08 0 2.17845e-08 0.0007 2.17875e-08 0 2.19615e-08 0 2.19645e-08 0.0007 2.19675e-08 0 2.21415e-08 0 2.21445e-08 0.0007 2.21475e-08 0 2.23215e-08 0 2.23245e-08 0.0007 2.23275e-08 0 2.25015e-08 0 2.25045e-08 0.0007 2.25075e-08 0 2.26815e-08 0 2.26845e-08 0.0007 2.26875e-08 0 2.28615e-08 0 2.28645e-08 0.0007 2.28675e-08 0 2.30415e-08 0 2.30445e-08 0.0007 2.30475e-08 0 2.32215e-08 0 2.32245e-08 0.0007 2.32275e-08 0 2.34015e-08 0 2.34045e-08 0.0007 2.34075e-08 0 2.35815e-08 0 2.35845e-08 0.0007 2.35875e-08 0 2.37615e-08 0 2.37645e-08 0.0007 2.37675e-08 0 2.39415e-08 0 2.39445e-08 0.0007 2.39475e-08 0 2.41215e-08 0 2.41245e-08 0.0007 2.41275e-08 0 2.43015e-08 0 2.43045e-08 0.0007 2.43075e-08 0 2.44815e-08 0 2.44845e-08 0.0007 2.44875e-08 0 2.46615e-08 0 2.46645e-08 0.0007 2.46675e-08 0 2.48415e-08 0 2.48445e-08 0.0007 2.48475e-08 0 2.50215e-08 0 2.50245e-08 0.0007 2.50275e-08 0 2.52015e-08 0 2.52045e-08 0.0007 2.52075e-08 0 2.53815e-08 0 2.53845e-08 0.0007 2.53875e-08 0 2.55615e-08 0 2.55645e-08 0.0007 2.55675e-08 0 2.57415e-08 0 2.57445e-08 0.0007 2.57475e-08 0 2.59215e-08 0 2.59245e-08 0.0007 2.59275e-08 0 2.61015e-08 0 2.61045e-08 0.0007 2.61075e-08 0 2.62815e-08 0 2.62845e-08 0.0007 2.62875e-08 0 2.64615e-08 0 2.64645e-08 0.0007 2.64675e-08 0 2.66415e-08 0 2.66445e-08 0.0007 2.66475e-08 0 2.68215e-08 0 2.68245e-08 0.0007 2.68275e-08 0 2.70015e-08 0 2.70045e-08 0.0007 2.70075e-08 0 2.71815e-08 0 2.71845e-08 0.0007 2.71875e-08 0 2.73615e-08 0 2.73645e-08 0.0007 2.73675e-08 0 2.75415e-08 0 2.75445e-08 0.0007 2.75475e-08 0 2.77215e-08 0 2.77245e-08 0.0007 2.77275e-08 0 2.79015e-08 0 2.79045e-08 0.0007 2.79075e-08 0 2.80815e-08 0 2.80845e-08 0.0007 2.80875e-08 0 2.82615e-08 0 2.82645e-08 0.0007 2.82675e-08 0 2.84415e-08 0 2.84445e-08 0.0007 2.84475e-08 0 2.86215e-08 0 2.86245e-08 0.0007 2.86275e-08 0 2.88015e-08 0 2.88045e-08 0.0007 2.88075e-08 0 2.89815e-08 0 2.89845e-08 0.0007 2.89875e-08 0 2.91615e-08 0 2.91645e-08 0.0007 2.91675e-08 0 2.93415e-08 0 2.93445e-08 0.0007 2.93475e-08 0 2.95215e-08 0 2.95245e-08 0.0007 2.95275e-08 0 2.97015e-08 0 2.97045e-08 0.0007 2.97075e-08 0 2.98815e-08 0 2.98845e-08 0.0007 2.98875e-08 0 3.00615e-08 0 3.00645e-08 0.0007 3.00675e-08 0 3.02415e-08 0 3.02445e-08 0.0007 3.02475e-08 0 3.04215e-08 0 3.04245e-08 0.0007 3.04275e-08 0 3.06015e-08 0 3.06045e-08 0.0007 3.06075e-08 0 3.07815e-08 0 3.07845e-08 0.0007 3.07875e-08 0 3.09615e-08 0 3.09645e-08 0.0007 3.09675e-08 0 3.11415e-08 0 3.11445e-08 0.0007 3.11475e-08 0 3.13215e-08 0 3.13245e-08 0.0007 3.13275e-08 0 3.15015e-08 0 3.15045e-08 0.0007 3.15075e-08 0 3.16815e-08 0 3.16845e-08 0.0007 3.16875e-08 0 3.18615e-08 0 3.18645e-08 0.0007 3.18675e-08 0 3.20415e-08 0 3.20445e-08 0.0007 3.20475e-08 0 3.22215e-08 0 3.22245e-08 0.0007 3.22275e-08 0 3.24015e-08 0 3.24045e-08 0.0007 3.24075e-08 0 3.25815e-08 0 3.25845e-08 0.0007 3.25875e-08 0 3.27615e-08 0 3.27645e-08 0.0007 3.27675e-08 0 3.29415e-08 0 3.29445e-08 0.0007 3.29475e-08 0 3.31215e-08 0 3.31245e-08 0.0007 3.31275e-08 0 3.33015e-08 0 3.33045e-08 0.0007 3.33075e-08 0 3.34815e-08 0 3.34845e-08 0.0007 3.34875e-08 0 3.36615e-08 0 3.36645e-08 0.0007 3.36675e-08 0 3.38415e-08 0 3.38445e-08 0.0007 3.38475e-08 0 3.40215e-08 0 3.40245e-08 0.0007 3.40275e-08 0 3.42015e-08 0 3.42045e-08 0.0007 3.42075e-08 0 3.43815e-08 0 3.43845e-08 0.0007 3.43875e-08 0 3.45615e-08 0 3.45645e-08 0.0007 3.45675e-08 0 3.47415e-08 0 3.47445e-08 0.0007 3.47475e-08 0 3.49215e-08 0 3.49245e-08 0.0007 3.49275e-08 0 3.51015e-08 0 3.51045e-08 0.0007 3.51075e-08 0 3.52815e-08 0 3.52845e-08 0.0007 3.52875e-08 0 3.54615e-08 0 3.54645e-08 0.0007 3.54675e-08 0 3.56415e-08 0 3.56445e-08 0.0007 3.56475e-08 0 3.58215e-08 0 3.58245e-08 0.0007 3.58275e-08 0 3.60015e-08 0 3.60045e-08 0.0007 3.60075e-08 0 3.61815e-08 0 3.61845e-08 0.0007 3.61875e-08 0 3.63615e-08 0 3.63645e-08 0.0007 3.63675e-08 0 3.65415e-08 0 3.65445e-08 0.0007 3.65475e-08 0 3.67215e-08 0 3.67245e-08 0.0007 3.67275e-08 0 3.69015e-08 0 3.69045e-08 0.0007 3.69075e-08 0 3.70815e-08 0 3.70845e-08 0.0007 3.70875e-08 0 3.72615e-08 0 3.72645e-08 0.0007 3.72675e-08 0 3.74415e-08 0 3.74445e-08 0.0007 3.74475e-08 0 3.76215e-08 0 3.76245e-08 0.0007 3.76275e-08 0 3.78015e-08 0 3.78045e-08 0.0007 3.78075e-08 0 3.79815e-08 0 3.79845e-08 0.0007 3.79875e-08 0 3.81615e-08 0 3.81645e-08 0.0007 3.81675e-08 0 3.83415e-08 0 3.83445e-08 0.0007 3.83475e-08 0 3.85215e-08 0 3.85245e-08 0.0007 3.85275e-08 0 3.87015e-08 0 3.87045e-08 0.0007 3.87075e-08 0 3.88815e-08 0 3.88845e-08 0.0007 3.88875e-08 0 3.90615e-08 0 3.90645e-08 0.0007 3.90675e-08 0 3.92415e-08 0 3.92445e-08 0.0007 3.92475e-08 0 3.94215e-08 0 3.94245e-08 0.0007 3.94275e-08 0 3.96015e-08 0 3.96045e-08 0.0007 3.96075e-08 0 3.97815e-08 0 3.97845e-08 0.0007 3.97875e-08 0 3.99615e-08 0 3.99645e-08 0.0007 3.99675e-08 0 4.01415e-08 0 4.01445e-08 0.0007 4.01475e-08 0 4.03215e-08 0 4.03245e-08 0.0007 4.03275e-08 0 4.05015e-08 0 4.05045e-08 0.0007 4.05075e-08 0 4.06815e-08 0 4.06845e-08 0.0007 4.06875e-08 0 4.08615e-08 0 4.08645e-08 0.0007 4.08675e-08 0 4.10415e-08 0 4.10445e-08 0.0007 4.10475e-08 0 4.12215e-08 0 4.12245e-08 0.0007 4.12275e-08 0 4.14015e-08 0 4.14045e-08 0.0007 4.14075e-08 0 4.15815e-08 0 4.15845e-08 0.0007 4.15875e-08 0 4.17615e-08 0 4.17645e-08 0.0007 4.17675e-08 0 4.19415e-08 0 4.19445e-08 0.0007 4.19475e-08 0 4.21215e-08 0 4.21245e-08 0.0007 4.21275e-08 0 4.23015e-08 0 4.23045e-08 0.0007 4.23075e-08 0 4.24815e-08 0 4.24845e-08 0.0007 4.24875e-08 0 4.26615e-08 0 4.26645e-08 0.0007 4.26675e-08 0 4.28415e-08 0 4.28445e-08 0.0007 4.28475e-08 0 4.30215e-08 0 4.30245e-08 0.0007 4.30275e-08 0 4.32015e-08 0 4.32045e-08 0.0007 4.32075e-08 0 4.33815e-08 0 4.33845e-08 0.0007 4.33875e-08 0 4.35615e-08 0 4.35645e-08 0.0007 4.35675e-08 0 4.37415e-08 0 4.37445e-08 0.0007 4.37475e-08 0 4.39215e-08 0 4.39245e-08 0.0007 4.39275e-08 0 4.41015e-08 0 4.41045e-08 0.0007 4.41075e-08 0 4.42815e-08 0 4.42845e-08 0.0007 4.42875e-08 0 4.44615e-08 0 4.44645e-08 0.0007 4.44675e-08 0 4.46415e-08 0 4.46445e-08 0.0007 4.46475e-08 0 4.48215e-08 0 4.48245e-08 0.0007 4.48275e-08 0 4.50015e-08 0 4.50045e-08 0.0007 4.50075e-08 0 4.51815e-08 0 4.51845e-08 0.0007 4.51875e-08 0 4.53615e-08 0 4.53645e-08 0.0007 4.53675e-08 0 4.55415e-08 0 4.55445e-08 0.0007 4.55475e-08 0 4.57215e-08 0 4.57245e-08 0.0007 4.57275e-08 0 4.59015e-08 0 4.59045e-08 0.0007 4.59075e-08 0)
B_S4|1 _S4|1 _S4|2 JJMIT AREA=2.5
B_S4|2 _S4|4 _S4|5 JJMIT AREA=1.61
B_S4|3 _S4|5 _S4|6 JJMIT AREA=1.54
B_S4|4 _S4|8 _S4|9 JJMIT AREA=1.69
B_S4|5 _S4|10 _S4|8 JJMIT AREA=1.38
B_S4|6 _S4|11 _S4|12 JJMIT AREA=2.5
B_S4|7 _S4|14 _S4|15 JJMIT AREA=2.5
I_S4|B1 0 _S4|3  PWL(0 0 5e-12 0.000175)
I_S4|B2 0 _S4|7  PWL(0 0 5e-12 0.000173)
I_S4|B3 0 _S4|13  PWL(0 0 5e-12 0.000175)
I_S4|B4 0 _S4|16  PWL(0 0 5e-12 0.000175)
L_S4|B1 _S4|3 _S4|1  2e-12
L_S4|B2 _S4|7 _S4|5  2e-12
L_S4|B3 _S4|11 _S4|13  2e-12
L_S4|B4 _S4|16 _S4|14  2e-12
L_S4|1 G3_2_RX _S4|1  2.059e-12
L_S4|2 _S4|1 _S4|4  4.123e-12
L_S4|3 _S4|5 _S4|8  6.873e-12
L_S4|4 _S4|10 _S4|11  5.195e-12
L_S4|5 T16 _S4|11  2.071e-12
L_S4|6 _S4|8 _S4|14  3.287e-12
L_S4|7 _S4|14 S4  2.066e-12
L_S4|P1 _S4|2 0  5.042e-13
L_S4|P3 _S4|6 0  5.799e-13
L_S4|P4 _S4|9 0  5.733e-13
L_S4|P6 _S4|12 0  4.605e-13
L_S4|P7 _S4|15 0  4.961e-13
R_S4|B1 _S4|1 _S4|101  2.7439617672
L_S4|RB1 _S4|101 0  1.550338398468e-12
R_S4|B2 _S4|4 _S4|104  4.260810197515528
L_S4|RB2 _S4|104 _S4|5  2.407357761596273e-12
R_S4|B3 _S4|5 _S4|105  4.454483388311688
L_S4|RB3 _S4|105 0  2.516783114396104e-12
R_S4|B4 _S4|8 _S4|108  4.059115040236686
L_S4|RB4 _S4|108 0  2.2933999977337278e-12
R_S4|B5 _S4|10 _S4|110  4.970945230434783
L_S4|RB5 _S4|110 _S4|8  2.8085840551956523e-12
R_S4|B6 _S4|11 _S4|111  2.7439617672
L_S4|RB6 _S4|111 0  1.550338398468e-12
R_S4|B7 _S4|14 _S4|114  2.7439617672
L_S4|RB7 _S4|114 0  1.550338398468e-12
II0|_SPL_A|B1 0 I0|_SPL_A|3  PWL(0 0 5e-12 0.000175)
II0|_SPL_A|B2 0 I0|_SPL_A|6  PWL(0 0 5e-12 0.00028)
II0|_SPL_A|B3 0 I0|_SPL_A|10  PWL(0 0 5e-12 0.000175)
II0|_SPL_A|B4 0 I0|_SPL_A|13  PWL(0 0 5e-12 0.000175)
LI0|_SPL_A|B1 I0|_SPL_A|3 I0|_SPL_A|1  9.175e-13
LI0|_SPL_A|B2 I0|_SPL_A|6 I0|_SPL_A|4  7.666e-13
LI0|_SPL_A|B3 I0|_SPL_A|10 I0|_SPL_A|8  1.928e-12
LI0|_SPL_A|B4 I0|_SPL_A|13 I0|_SPL_A|11  8.786e-13
BI0|_SPL_A|1 I0|_SPL_A|1 I0|_SPL_A|2 JJMIT AREA=2.5
BI0|_SPL_A|2 I0|_SPL_A|4 I0|_SPL_A|5 JJMIT AREA=3.0
BI0|_SPL_A|3 I0|_SPL_A|8 I0|_SPL_A|9 JJMIT AREA=2.5
BI0|_SPL_A|4 I0|_SPL_A|11 I0|_SPL_A|12 JJMIT AREA=2.5
LI0|_SPL_A|1 A0 I0|_SPL_A|1  2.063e-12
LI0|_SPL_A|2 I0|_SPL_A|1 I0|_SPL_A|4  3.637e-12
LI0|_SPL_A|3 I0|_SPL_A|4 I0|_SPL_A|7  1.278e-12
LI0|_SPL_A|4 I0|_SPL_A|7 I0|_SPL_A|8  1.305e-12
LI0|_SPL_A|5 I0|_SPL_A|8 I0|A1  2.05e-12
LI0|_SPL_A|6 I0|_SPL_A|7 I0|_SPL_A|11  1.315e-12
LI0|_SPL_A|7 I0|_SPL_A|11 I0|A2  2.06e-12
LI0|_SPL_A|P1 I0|_SPL_A|2 0  4.676e-13
LI0|_SPL_A|P2 I0|_SPL_A|5 0  4.498e-13
LI0|_SPL_A|P3 I0|_SPL_A|9 0  5.183e-13
LI0|_SPL_A|P4 I0|_SPL_A|12 0  4.639e-13
RI0|_SPL_A|B1 I0|_SPL_A|1 I0|_SPL_A|101  2.7439617672
LI0|_SPL_A|RB1 I0|_SPL_A|101 0  1.550338398468e-12
RI0|_SPL_A|B2 I0|_SPL_A|4 I0|_SPL_A|104  2.286634806
LI0|_SPL_A|RB2 I0|_SPL_A|104 0  1.29194866539e-12
RI0|_SPL_A|B3 I0|_SPL_A|8 I0|_SPL_A|108  2.7439617672
LI0|_SPL_A|RB3 I0|_SPL_A|108 0  1.550338398468e-12
RI0|_SPL_A|B4 I0|_SPL_A|11 I0|_SPL_A|111  2.7439617672
LI0|_SPL_A|RB4 I0|_SPL_A|111 0  1.550338398468e-12
II0|_SPL_B|B1 0 I0|_SPL_B|3  PWL(0 0 5e-12 0.000175)
II0|_SPL_B|B2 0 I0|_SPL_B|6  PWL(0 0 5e-12 0.00028)
II0|_SPL_B|B3 0 I0|_SPL_B|10  PWL(0 0 5e-12 0.000175)
II0|_SPL_B|B4 0 I0|_SPL_B|13  PWL(0 0 5e-12 0.000175)
LI0|_SPL_B|B1 I0|_SPL_B|3 I0|_SPL_B|1  9.175e-13
LI0|_SPL_B|B2 I0|_SPL_B|6 I0|_SPL_B|4  7.666e-13
LI0|_SPL_B|B3 I0|_SPL_B|10 I0|_SPL_B|8  1.928e-12
LI0|_SPL_B|B4 I0|_SPL_B|13 I0|_SPL_B|11  8.786e-13
BI0|_SPL_B|1 I0|_SPL_B|1 I0|_SPL_B|2 JJMIT AREA=2.5
BI0|_SPL_B|2 I0|_SPL_B|4 I0|_SPL_B|5 JJMIT AREA=3.0
BI0|_SPL_B|3 I0|_SPL_B|8 I0|_SPL_B|9 JJMIT AREA=2.5
BI0|_SPL_B|4 I0|_SPL_B|11 I0|_SPL_B|12 JJMIT AREA=2.5
LI0|_SPL_B|1 B0 I0|_SPL_B|1  2.063e-12
LI0|_SPL_B|2 I0|_SPL_B|1 I0|_SPL_B|4  3.637e-12
LI0|_SPL_B|3 I0|_SPL_B|4 I0|_SPL_B|7  1.278e-12
LI0|_SPL_B|4 I0|_SPL_B|7 I0|_SPL_B|8  1.305e-12
LI0|_SPL_B|5 I0|_SPL_B|8 I0|B1  2.05e-12
LI0|_SPL_B|6 I0|_SPL_B|7 I0|_SPL_B|11  1.315e-12
LI0|_SPL_B|7 I0|_SPL_B|11 I0|B2  2.06e-12
LI0|_SPL_B|P1 I0|_SPL_B|2 0  4.676e-13
LI0|_SPL_B|P2 I0|_SPL_B|5 0  4.498e-13
LI0|_SPL_B|P3 I0|_SPL_B|9 0  5.183e-13
LI0|_SPL_B|P4 I0|_SPL_B|12 0  4.639e-13
RI0|_SPL_B|B1 I0|_SPL_B|1 I0|_SPL_B|101  2.7439617672
LI0|_SPL_B|RB1 I0|_SPL_B|101 0  1.550338398468e-12
RI0|_SPL_B|B2 I0|_SPL_B|4 I0|_SPL_B|104  2.286634806
LI0|_SPL_B|RB2 I0|_SPL_B|104 0  1.29194866539e-12
RI0|_SPL_B|B3 I0|_SPL_B|8 I0|_SPL_B|108  2.7439617672
LI0|_SPL_B|RB3 I0|_SPL_B|108 0  1.550338398468e-12
RI0|_SPL_B|B4 I0|_SPL_B|11 I0|_SPL_B|111  2.7439617672
LI0|_SPL_B|RB4 I0|_SPL_B|111 0  1.550338398468e-12
BI0|_DFF_A|1 I0|_DFF_A|1 I0|_DFF_A|2 JJMIT AREA=2.5
BI0|_DFF_A|2 I0|_DFF_A|4 I0|_DFF_A|5 JJMIT AREA=1.61
BI0|_DFF_A|3 I0|_DFF_A|5 I0|_DFF_A|6 JJMIT AREA=1.54
BI0|_DFF_A|4 I0|_DFF_A|8 I0|_DFF_A|9 JJMIT AREA=1.69
BI0|_DFF_A|5 I0|_DFF_A|10 I0|_DFF_A|8 JJMIT AREA=1.38
BI0|_DFF_A|6 I0|_DFF_A|11 I0|_DFF_A|12 JJMIT AREA=2.5
BI0|_DFF_A|7 I0|_DFF_A|14 I0|_DFF_A|15 JJMIT AREA=2.5
II0|_DFF_A|B1 0 I0|_DFF_A|3  PWL(0 0 5e-12 0.000175)
II0|_DFF_A|B2 0 I0|_DFF_A|7  PWL(0 0 5e-12 0.000173)
II0|_DFF_A|B3 0 I0|_DFF_A|13  PWL(0 0 5e-12 0.000175)
II0|_DFF_A|B4 0 I0|_DFF_A|16  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|B1 I0|_DFF_A|3 I0|_DFF_A|1  2e-12
LI0|_DFF_A|B2 I0|_DFF_A|7 I0|_DFF_A|5  2e-12
LI0|_DFF_A|B3 I0|_DFF_A|11 I0|_DFF_A|13  2e-12
LI0|_DFF_A|B4 I0|_DFF_A|16 I0|_DFF_A|14  2e-12
LI0|_DFF_A|1 I0|A1 I0|_DFF_A|1  2.059e-12
LI0|_DFF_A|2 I0|_DFF_A|1 I0|_DFF_A|4  4.123e-12
LI0|_DFF_A|3 I0|_DFF_A|5 I0|_DFF_A|8  6.873e-12
LI0|_DFF_A|4 I0|_DFF_A|10 I0|_DFF_A|11  5.195e-12
LI0|_DFF_A|5 T00 I0|_DFF_A|11  2.071e-12
LI0|_DFF_A|6 I0|_DFF_A|8 I0|_DFF_A|14  3.287e-12
LI0|_DFF_A|7 I0|_DFF_A|14 I0|A1_SYNC  2.066e-12
LI0|_DFF_A|P1 I0|_DFF_A|2 0  5.042e-13
LI0|_DFF_A|P3 I0|_DFF_A|6 0  5.799e-13
LI0|_DFF_A|P4 I0|_DFF_A|9 0  5.733e-13
LI0|_DFF_A|P6 I0|_DFF_A|12 0  4.605e-13
LI0|_DFF_A|P7 I0|_DFF_A|15 0  4.961e-13
RI0|_DFF_A|B1 I0|_DFF_A|1 I0|_DFF_A|101  2.7439617672
LI0|_DFF_A|RB1 I0|_DFF_A|101 0  1.550338398468e-12
RI0|_DFF_A|B2 I0|_DFF_A|4 I0|_DFF_A|104  4.260810197515528
LI0|_DFF_A|RB2 I0|_DFF_A|104 I0|_DFF_A|5  2.407357761596273e-12
RI0|_DFF_A|B3 I0|_DFF_A|5 I0|_DFF_A|105  4.454483388311688
LI0|_DFF_A|RB3 I0|_DFF_A|105 0  2.516783114396104e-12
RI0|_DFF_A|B4 I0|_DFF_A|8 I0|_DFF_A|108  4.059115040236686
LI0|_DFF_A|RB4 I0|_DFF_A|108 0  2.2933999977337278e-12
RI0|_DFF_A|B5 I0|_DFF_A|10 I0|_DFF_A|110  4.970945230434783
LI0|_DFF_A|RB5 I0|_DFF_A|110 I0|_DFF_A|8  2.8085840551956523e-12
RI0|_DFF_A|B6 I0|_DFF_A|11 I0|_DFF_A|111  2.7439617672
LI0|_DFF_A|RB6 I0|_DFF_A|111 0  1.550338398468e-12
RI0|_DFF_A|B7 I0|_DFF_A|14 I0|_DFF_A|114  2.7439617672
LI0|_DFF_A|RB7 I0|_DFF_A|114 0  1.550338398468e-12
BI0|_DFF_B|1 I0|_DFF_B|1 I0|_DFF_B|2 JJMIT AREA=2.5
BI0|_DFF_B|2 I0|_DFF_B|4 I0|_DFF_B|5 JJMIT AREA=1.61
BI0|_DFF_B|3 I0|_DFF_B|5 I0|_DFF_B|6 JJMIT AREA=1.54
BI0|_DFF_B|4 I0|_DFF_B|8 I0|_DFF_B|9 JJMIT AREA=1.69
BI0|_DFF_B|5 I0|_DFF_B|10 I0|_DFF_B|8 JJMIT AREA=1.38
BI0|_DFF_B|6 I0|_DFF_B|11 I0|_DFF_B|12 JJMIT AREA=2.5
BI0|_DFF_B|7 I0|_DFF_B|14 I0|_DFF_B|15 JJMIT AREA=2.5
II0|_DFF_B|B1 0 I0|_DFF_B|3  PWL(0 0 5e-12 0.000175)
II0|_DFF_B|B2 0 I0|_DFF_B|7  PWL(0 0 5e-12 0.000173)
II0|_DFF_B|B3 0 I0|_DFF_B|13  PWL(0 0 5e-12 0.000175)
II0|_DFF_B|B4 0 I0|_DFF_B|16  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|B1 I0|_DFF_B|3 I0|_DFF_B|1  2e-12
LI0|_DFF_B|B2 I0|_DFF_B|7 I0|_DFF_B|5  2e-12
LI0|_DFF_B|B3 I0|_DFF_B|11 I0|_DFF_B|13  2e-12
LI0|_DFF_B|B4 I0|_DFF_B|16 I0|_DFF_B|14  2e-12
LI0|_DFF_B|1 I0|B1 I0|_DFF_B|1  2.059e-12
LI0|_DFF_B|2 I0|_DFF_B|1 I0|_DFF_B|4  4.123e-12
LI0|_DFF_B|3 I0|_DFF_B|5 I0|_DFF_B|8  6.873e-12
LI0|_DFF_B|4 I0|_DFF_B|10 I0|_DFF_B|11  5.195e-12
LI0|_DFF_B|5 T00 I0|_DFF_B|11  2.071e-12
LI0|_DFF_B|6 I0|_DFF_B|8 I0|_DFF_B|14  3.287e-12
LI0|_DFF_B|7 I0|_DFF_B|14 I0|B1_SYNC  2.066e-12
LI0|_DFF_B|P1 I0|_DFF_B|2 0  5.042e-13
LI0|_DFF_B|P3 I0|_DFF_B|6 0  5.799e-13
LI0|_DFF_B|P4 I0|_DFF_B|9 0  5.733e-13
LI0|_DFF_B|P6 I0|_DFF_B|12 0  4.605e-13
LI0|_DFF_B|P7 I0|_DFF_B|15 0  4.961e-13
RI0|_DFF_B|B1 I0|_DFF_B|1 I0|_DFF_B|101  2.7439617672
LI0|_DFF_B|RB1 I0|_DFF_B|101 0  1.550338398468e-12
RI0|_DFF_B|B2 I0|_DFF_B|4 I0|_DFF_B|104  4.260810197515528
LI0|_DFF_B|RB2 I0|_DFF_B|104 I0|_DFF_B|5  2.407357761596273e-12
RI0|_DFF_B|B3 I0|_DFF_B|5 I0|_DFF_B|105  4.454483388311688
LI0|_DFF_B|RB3 I0|_DFF_B|105 0  2.516783114396104e-12
RI0|_DFF_B|B4 I0|_DFF_B|8 I0|_DFF_B|108  4.059115040236686
LI0|_DFF_B|RB4 I0|_DFF_B|108 0  2.2933999977337278e-12
RI0|_DFF_B|B5 I0|_DFF_B|10 I0|_DFF_B|110  4.970945230434783
LI0|_DFF_B|RB5 I0|_DFF_B|110 I0|_DFF_B|8  2.8085840551956523e-12
RI0|_DFF_B|B6 I0|_DFF_B|11 I0|_DFF_B|111  2.7439617672
LI0|_DFF_B|RB6 I0|_DFF_B|111 0  1.550338398468e-12
RI0|_DFF_B|B7 I0|_DFF_B|14 I0|_DFF_B|114  2.7439617672
LI0|_DFF_B|RB7 I0|_DFF_B|114 0  1.550338398468e-12
BI0|_XOR|1 I0|_XOR|1 I0|_XOR|2 JJMIT AREA=2.5
BI0|_XOR|2 I0|_XOR|4 I0|_XOR|5 JJMIT AREA=2.09
BI0|_XOR|3 I0|_XOR|25 I0|_XOR|6 JJMIT AREA=1.71
BI0|_XOR|4 I0|_XOR|9 I0|_XOR|10 JJMIT AREA=2.5
BI0|_XOR|5 I0|_XOR|12 I0|_XOR|13 JJMIT AREA=2.09
BI0|_XOR|6 I0|_XOR|26 I0|_XOR|14 JJMIT AREA=1.71
BI0|_XOR|7 I0|_XOR|27 I0|_XOR|16 JJMIT AREA=1.62
BI0|_XOR|8 I0|_XOR|17 I0|_XOR|18 JJMIT AREA=2.5
BI0|_XOR|9 I0|_XOR|20 I0|_XOR|16 JJMIT AREA=1.45
BI0|_XOR|10 I0|_XOR|16 I0|_XOR|21 JJMIT AREA=0.89
BI0|_XOR|11 I0|_XOR|22 I0|_XOR|23 JJMIT AREA=2.5
II0|_XOR|B1 0 I0|_XOR|3  PWL(0 0 5e-12 0.000175)
II0|_XOR|B2 0 I0|_XOR|7  PWL(0 0 5e-12 0.000112)
II0|_XOR|B3 0 I0|_XOR|11  PWL(0 0 5e-12 0.000175)
II0|_XOR|B4 0 I0|_XOR|15  PWL(0 0 5e-12 0.000112)
II0|_XOR|B5 0 I0|_XOR|19  PWL(0 0 5e-12 0.000175)
II0|_XOR|B6 0 I0|_XOR|24  PWL(0 0 5e-12 0.000175)
LI0|_XOR|B1 I0|_XOR|3 I0|_XOR|1  2e-12
LI0|_XOR|B2 I0|_XOR|7 I0|_XOR|6  2e-12
LI0|_XOR|B3 I0|_XOR|11 I0|_XOR|9  2e-12
LI0|_XOR|B4 I0|_XOR|15 I0|_XOR|14  2e-12
LI0|_XOR|B5 I0|_XOR|19 I0|_XOR|17  2e-12
LI0|_XOR|B6 I0|_XOR|24 I0|_XOR|22  2e-12
LI0|_XOR|1 I0|A2 I0|_XOR|1  2.06e-12
LI0|_XOR|2 I0|_XOR|1 I0|_XOR|4  3.233e-12
LI0|_XOR|3 I0|_XOR|4 I0|_XOR|25  1.419e-12
LI0|_XOR|4 I0|_XOR|6 I0|_XOR|8  6.051e-12
LI0|_XOR|5 I0|B2 I0|_XOR|9  2.092e-12
LI0|_XOR|6 I0|_XOR|9 I0|_XOR|12  3.221e-12
LI0|_XOR|7 I0|_XOR|12 I0|_XOR|26  1.384e-12
LI0|_XOR|8 I0|_XOR|14 I0|_XOR|8  6.059e-12
LI0|_XOR|9 I0|_XOR|8 I0|_XOR|27  1.301e-12
LI0|_XOR|10 T00 I0|_XOR|17  2.082e-12
LI0|_XOR|11 I0|_XOR|17 I0|_XOR|20  1.43e-12
LI0|_XOR|12 I0|_XOR|16 I0|_XOR|22  3.892e-12
LI0|_XOR|13 I0|_XOR|22 IP0_0  2.077e-12
LI0|_XOR|P1 I0|_XOR|2 0  5.508e-13
LI0|_XOR|P2 I0|_XOR|5 0  4.769e-13
LI0|_XOR|P4 I0|_XOR|10 0  4.767e-13
LI0|_XOR|P5 I0|_XOR|13 0  4.812e-13
LI0|_XOR|P8 I0|_XOR|18 0  4.526e-13
LI0|_XOR|P10 I0|_XOR|21 0  5.69e-13
LI0|_XOR|P11 I0|_XOR|23 0  4.746e-13
RI0|_XOR|B1 I0|_XOR|1 I0|_XOR|101  2.7439617672
LI0|_XOR|RB1 I0|_XOR|101 0  2.050338398468e-12
RI0|_XOR|B2 I0|_XOR|4 I0|_XOR|104  3.2822509177033496
LI0|_XOR|RB2 I0|_XOR|104 0  2.3544717685023925e-12
RI0|_XOR|B3 I0|_XOR|4 I0|_XOR|106  4.011640010526316
LI0|_XOR|RB3 I0|_XOR|106 I0|_XOR|6  2.766576605947368e-12
RI0|_XOR|B4 I0|_XOR|9 I0|_XOR|109  2.7439617672
LI0|_XOR|RB4 I0|_XOR|109 0  2.050338398468e-12
RI0|_XOR|B5 I0|_XOR|12 I0|_XOR|112  3.2822509177033496
LI0|_XOR|RB5 I0|_XOR|112 0  2.3544717685023925e-12
RI0|_XOR|B6 I0|_XOR|12 I0|_XOR|114  4.011640010526316
LI0|_XOR|RB6 I0|_XOR|114 I0|_XOR|14  2.766576605947368e-12
RI0|_XOR|B7 I0|_XOR|8 I0|_XOR|108  4.2345089
LI0|_XOR|RB7 I0|_XOR|108 I0|_XOR|16  2.8924975284999997e-12
RI0|_XOR|B8 I0|_XOR|17 I0|_XOR|117  2.7439617672
LI0|_XOR|RB8 I0|_XOR|117 0  2.050338398468e-12
RI0|_XOR|B9 I0|_XOR|20 I0|_XOR|120  4.730968564137931
LI0|_XOR|RB9 I0|_XOR|120 I0|_XOR|16  3.172997238737931e-12
RI0|_XOR|B10 I0|_XOR|16 I0|_XOR|116  7.707757773033708
LI0|_XOR|RB10 I0|_XOR|116 0  4.854883141764045e-12
RI0|_XOR|B11 I0|_XOR|22 I0|_XOR|122  2.7439617672
LI0|_XOR|RB11 I0|_XOR|122 0  2.050338398468e-12
LI0|_AND|A1 I0|A1_SYNC I0|_AND|A1  2.067833848e-12
LI0|_AND|A2 I0|_AND|A1 I0|_AND|A2  4.135667696e-12
LI0|_AND|A3 I0|_AND|A3 I0|_AND|Q3  1.2e-12
LI0|_AND|B1 I0|B1_SYNC I0|_AND|B1  2.067833848e-12
LI0|_AND|B2 I0|_AND|B1 I0|_AND|B2  4.135667696e-12
LI0|_AND|B3 I0|_AND|B3 I0|_AND|Q3  1.2e-12
LI0|_AND|Q3 I0|_AND|Q3 I0|_AND|Q2  4.135667696e-12
LI0|_AND|Q2 I0|_AND|Q2 I0|_AND|Q1  4.135667696e-12
LI0|_AND|Q1 I0|_AND|Q1 IG0_0  2.067833848e-12
II1|_SPL_A|B1 0 I1|_SPL_A|3  PWL(0 0 5e-12 0.000175)
II1|_SPL_A|B2 0 I1|_SPL_A|6  PWL(0 0 5e-12 0.00028)
II1|_SPL_A|B3 0 I1|_SPL_A|10  PWL(0 0 5e-12 0.000175)
II1|_SPL_A|B4 0 I1|_SPL_A|13  PWL(0 0 5e-12 0.000175)
LI1|_SPL_A|B1 I1|_SPL_A|3 I1|_SPL_A|1  9.175e-13
LI1|_SPL_A|B2 I1|_SPL_A|6 I1|_SPL_A|4  7.666e-13
LI1|_SPL_A|B3 I1|_SPL_A|10 I1|_SPL_A|8  1.928e-12
LI1|_SPL_A|B4 I1|_SPL_A|13 I1|_SPL_A|11  8.786e-13
BI1|_SPL_A|1 I1|_SPL_A|1 I1|_SPL_A|2 JJMIT AREA=2.5
BI1|_SPL_A|2 I1|_SPL_A|4 I1|_SPL_A|5 JJMIT AREA=3.0
BI1|_SPL_A|3 I1|_SPL_A|8 I1|_SPL_A|9 JJMIT AREA=2.5
BI1|_SPL_A|4 I1|_SPL_A|11 I1|_SPL_A|12 JJMIT AREA=2.5
LI1|_SPL_A|1 A1 I1|_SPL_A|1  2.063e-12
LI1|_SPL_A|2 I1|_SPL_A|1 I1|_SPL_A|4  3.637e-12
LI1|_SPL_A|3 I1|_SPL_A|4 I1|_SPL_A|7  1.278e-12
LI1|_SPL_A|4 I1|_SPL_A|7 I1|_SPL_A|8  1.305e-12
LI1|_SPL_A|5 I1|_SPL_A|8 I1|A1  2.05e-12
LI1|_SPL_A|6 I1|_SPL_A|7 I1|_SPL_A|11  1.315e-12
LI1|_SPL_A|7 I1|_SPL_A|11 I1|A2  2.06e-12
LI1|_SPL_A|P1 I1|_SPL_A|2 0  4.676e-13
LI1|_SPL_A|P2 I1|_SPL_A|5 0  4.498e-13
LI1|_SPL_A|P3 I1|_SPL_A|9 0  5.183e-13
LI1|_SPL_A|P4 I1|_SPL_A|12 0  4.639e-13
RI1|_SPL_A|B1 I1|_SPL_A|1 I1|_SPL_A|101  2.7439617672
LI1|_SPL_A|RB1 I1|_SPL_A|101 0  1.550338398468e-12
RI1|_SPL_A|B2 I1|_SPL_A|4 I1|_SPL_A|104  2.286634806
LI1|_SPL_A|RB2 I1|_SPL_A|104 0  1.29194866539e-12
RI1|_SPL_A|B3 I1|_SPL_A|8 I1|_SPL_A|108  2.7439617672
LI1|_SPL_A|RB3 I1|_SPL_A|108 0  1.550338398468e-12
RI1|_SPL_A|B4 I1|_SPL_A|11 I1|_SPL_A|111  2.7439617672
LI1|_SPL_A|RB4 I1|_SPL_A|111 0  1.550338398468e-12
II1|_SPL_B|B1 0 I1|_SPL_B|3  PWL(0 0 5e-12 0.000175)
II1|_SPL_B|B2 0 I1|_SPL_B|6  PWL(0 0 5e-12 0.00028)
II1|_SPL_B|B3 0 I1|_SPL_B|10  PWL(0 0 5e-12 0.000175)
II1|_SPL_B|B4 0 I1|_SPL_B|13  PWL(0 0 5e-12 0.000175)
LI1|_SPL_B|B1 I1|_SPL_B|3 I1|_SPL_B|1  9.175e-13
LI1|_SPL_B|B2 I1|_SPL_B|6 I1|_SPL_B|4  7.666e-13
LI1|_SPL_B|B3 I1|_SPL_B|10 I1|_SPL_B|8  1.928e-12
LI1|_SPL_B|B4 I1|_SPL_B|13 I1|_SPL_B|11  8.786e-13
BI1|_SPL_B|1 I1|_SPL_B|1 I1|_SPL_B|2 JJMIT AREA=2.5
BI1|_SPL_B|2 I1|_SPL_B|4 I1|_SPL_B|5 JJMIT AREA=3.0
BI1|_SPL_B|3 I1|_SPL_B|8 I1|_SPL_B|9 JJMIT AREA=2.5
BI1|_SPL_B|4 I1|_SPL_B|11 I1|_SPL_B|12 JJMIT AREA=2.5
LI1|_SPL_B|1 B1 I1|_SPL_B|1  2.063e-12
LI1|_SPL_B|2 I1|_SPL_B|1 I1|_SPL_B|4  3.637e-12
LI1|_SPL_B|3 I1|_SPL_B|4 I1|_SPL_B|7  1.278e-12
LI1|_SPL_B|4 I1|_SPL_B|7 I1|_SPL_B|8  1.305e-12
LI1|_SPL_B|5 I1|_SPL_B|8 I1|B1  2.05e-12
LI1|_SPL_B|6 I1|_SPL_B|7 I1|_SPL_B|11  1.315e-12
LI1|_SPL_B|7 I1|_SPL_B|11 I1|B2  2.06e-12
LI1|_SPL_B|P1 I1|_SPL_B|2 0  4.676e-13
LI1|_SPL_B|P2 I1|_SPL_B|5 0  4.498e-13
LI1|_SPL_B|P3 I1|_SPL_B|9 0  5.183e-13
LI1|_SPL_B|P4 I1|_SPL_B|12 0  4.639e-13
RI1|_SPL_B|B1 I1|_SPL_B|1 I1|_SPL_B|101  2.7439617672
LI1|_SPL_B|RB1 I1|_SPL_B|101 0  1.550338398468e-12
RI1|_SPL_B|B2 I1|_SPL_B|4 I1|_SPL_B|104  2.286634806
LI1|_SPL_B|RB2 I1|_SPL_B|104 0  1.29194866539e-12
RI1|_SPL_B|B3 I1|_SPL_B|8 I1|_SPL_B|108  2.7439617672
LI1|_SPL_B|RB3 I1|_SPL_B|108 0  1.550338398468e-12
RI1|_SPL_B|B4 I1|_SPL_B|11 I1|_SPL_B|111  2.7439617672
LI1|_SPL_B|RB4 I1|_SPL_B|111 0  1.550338398468e-12
BI1|_DFF_A|1 I1|_DFF_A|1 I1|_DFF_A|2 JJMIT AREA=2.5
BI1|_DFF_A|2 I1|_DFF_A|4 I1|_DFF_A|5 JJMIT AREA=1.61
BI1|_DFF_A|3 I1|_DFF_A|5 I1|_DFF_A|6 JJMIT AREA=1.54
BI1|_DFF_A|4 I1|_DFF_A|8 I1|_DFF_A|9 JJMIT AREA=1.69
BI1|_DFF_A|5 I1|_DFF_A|10 I1|_DFF_A|8 JJMIT AREA=1.38
BI1|_DFF_A|6 I1|_DFF_A|11 I1|_DFF_A|12 JJMIT AREA=2.5
BI1|_DFF_A|7 I1|_DFF_A|14 I1|_DFF_A|15 JJMIT AREA=2.5
II1|_DFF_A|B1 0 I1|_DFF_A|3  PWL(0 0 5e-12 0.000175)
II1|_DFF_A|B2 0 I1|_DFF_A|7  PWL(0 0 5e-12 0.000173)
II1|_DFF_A|B3 0 I1|_DFF_A|13  PWL(0 0 5e-12 0.000175)
II1|_DFF_A|B4 0 I1|_DFF_A|16  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|B1 I1|_DFF_A|3 I1|_DFF_A|1  2e-12
LI1|_DFF_A|B2 I1|_DFF_A|7 I1|_DFF_A|5  2e-12
LI1|_DFF_A|B3 I1|_DFF_A|11 I1|_DFF_A|13  2e-12
LI1|_DFF_A|B4 I1|_DFF_A|16 I1|_DFF_A|14  2e-12
LI1|_DFF_A|1 I1|A1 I1|_DFF_A|1  2.059e-12
LI1|_DFF_A|2 I1|_DFF_A|1 I1|_DFF_A|4  4.123e-12
LI1|_DFF_A|3 I1|_DFF_A|5 I1|_DFF_A|8  6.873e-12
LI1|_DFF_A|4 I1|_DFF_A|10 I1|_DFF_A|11  5.195e-12
LI1|_DFF_A|5 T01 I1|_DFF_A|11  2.071e-12
LI1|_DFF_A|6 I1|_DFF_A|8 I1|_DFF_A|14  3.287e-12
LI1|_DFF_A|7 I1|_DFF_A|14 I1|A1_SYNC  2.066e-12
LI1|_DFF_A|P1 I1|_DFF_A|2 0  5.042e-13
LI1|_DFF_A|P3 I1|_DFF_A|6 0  5.799e-13
LI1|_DFF_A|P4 I1|_DFF_A|9 0  5.733e-13
LI1|_DFF_A|P6 I1|_DFF_A|12 0  4.605e-13
LI1|_DFF_A|P7 I1|_DFF_A|15 0  4.961e-13
RI1|_DFF_A|B1 I1|_DFF_A|1 I1|_DFF_A|101  2.7439617672
LI1|_DFF_A|RB1 I1|_DFF_A|101 0  1.550338398468e-12
RI1|_DFF_A|B2 I1|_DFF_A|4 I1|_DFF_A|104  4.260810197515528
LI1|_DFF_A|RB2 I1|_DFF_A|104 I1|_DFF_A|5  2.407357761596273e-12
RI1|_DFF_A|B3 I1|_DFF_A|5 I1|_DFF_A|105  4.454483388311688
LI1|_DFF_A|RB3 I1|_DFF_A|105 0  2.516783114396104e-12
RI1|_DFF_A|B4 I1|_DFF_A|8 I1|_DFF_A|108  4.059115040236686
LI1|_DFF_A|RB4 I1|_DFF_A|108 0  2.2933999977337278e-12
RI1|_DFF_A|B5 I1|_DFF_A|10 I1|_DFF_A|110  4.970945230434783
LI1|_DFF_A|RB5 I1|_DFF_A|110 I1|_DFF_A|8  2.8085840551956523e-12
RI1|_DFF_A|B6 I1|_DFF_A|11 I1|_DFF_A|111  2.7439617672
LI1|_DFF_A|RB6 I1|_DFF_A|111 0  1.550338398468e-12
RI1|_DFF_A|B7 I1|_DFF_A|14 I1|_DFF_A|114  2.7439617672
LI1|_DFF_A|RB7 I1|_DFF_A|114 0  1.550338398468e-12
BI1|_DFF_B|1 I1|_DFF_B|1 I1|_DFF_B|2 JJMIT AREA=2.5
BI1|_DFF_B|2 I1|_DFF_B|4 I1|_DFF_B|5 JJMIT AREA=1.61
BI1|_DFF_B|3 I1|_DFF_B|5 I1|_DFF_B|6 JJMIT AREA=1.54
BI1|_DFF_B|4 I1|_DFF_B|8 I1|_DFF_B|9 JJMIT AREA=1.69
BI1|_DFF_B|5 I1|_DFF_B|10 I1|_DFF_B|8 JJMIT AREA=1.38
BI1|_DFF_B|6 I1|_DFF_B|11 I1|_DFF_B|12 JJMIT AREA=2.5
BI1|_DFF_B|7 I1|_DFF_B|14 I1|_DFF_B|15 JJMIT AREA=2.5
II1|_DFF_B|B1 0 I1|_DFF_B|3  PWL(0 0 5e-12 0.000175)
II1|_DFF_B|B2 0 I1|_DFF_B|7  PWL(0 0 5e-12 0.000173)
II1|_DFF_B|B3 0 I1|_DFF_B|13  PWL(0 0 5e-12 0.000175)
II1|_DFF_B|B4 0 I1|_DFF_B|16  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|B1 I1|_DFF_B|3 I1|_DFF_B|1  2e-12
LI1|_DFF_B|B2 I1|_DFF_B|7 I1|_DFF_B|5  2e-12
LI1|_DFF_B|B3 I1|_DFF_B|11 I1|_DFF_B|13  2e-12
LI1|_DFF_B|B4 I1|_DFF_B|16 I1|_DFF_B|14  2e-12
LI1|_DFF_B|1 I1|B1 I1|_DFF_B|1  2.059e-12
LI1|_DFF_B|2 I1|_DFF_B|1 I1|_DFF_B|4  4.123e-12
LI1|_DFF_B|3 I1|_DFF_B|5 I1|_DFF_B|8  6.873e-12
LI1|_DFF_B|4 I1|_DFF_B|10 I1|_DFF_B|11  5.195e-12
LI1|_DFF_B|5 T01 I1|_DFF_B|11  2.071e-12
LI1|_DFF_B|6 I1|_DFF_B|8 I1|_DFF_B|14  3.287e-12
LI1|_DFF_B|7 I1|_DFF_B|14 I1|B1_SYNC  2.066e-12
LI1|_DFF_B|P1 I1|_DFF_B|2 0  5.042e-13
LI1|_DFF_B|P3 I1|_DFF_B|6 0  5.799e-13
LI1|_DFF_B|P4 I1|_DFF_B|9 0  5.733e-13
LI1|_DFF_B|P6 I1|_DFF_B|12 0  4.605e-13
LI1|_DFF_B|P7 I1|_DFF_B|15 0  4.961e-13
RI1|_DFF_B|B1 I1|_DFF_B|1 I1|_DFF_B|101  2.7439617672
LI1|_DFF_B|RB1 I1|_DFF_B|101 0  1.550338398468e-12
RI1|_DFF_B|B2 I1|_DFF_B|4 I1|_DFF_B|104  4.260810197515528
LI1|_DFF_B|RB2 I1|_DFF_B|104 I1|_DFF_B|5  2.407357761596273e-12
RI1|_DFF_B|B3 I1|_DFF_B|5 I1|_DFF_B|105  4.454483388311688
LI1|_DFF_B|RB3 I1|_DFF_B|105 0  2.516783114396104e-12
RI1|_DFF_B|B4 I1|_DFF_B|8 I1|_DFF_B|108  4.059115040236686
LI1|_DFF_B|RB4 I1|_DFF_B|108 0  2.2933999977337278e-12
RI1|_DFF_B|B5 I1|_DFF_B|10 I1|_DFF_B|110  4.970945230434783
LI1|_DFF_B|RB5 I1|_DFF_B|110 I1|_DFF_B|8  2.8085840551956523e-12
RI1|_DFF_B|B6 I1|_DFF_B|11 I1|_DFF_B|111  2.7439617672
LI1|_DFF_B|RB6 I1|_DFF_B|111 0  1.550338398468e-12
RI1|_DFF_B|B7 I1|_DFF_B|14 I1|_DFF_B|114  2.7439617672
LI1|_DFF_B|RB7 I1|_DFF_B|114 0  1.550338398468e-12
BI1|_XOR|1 I1|_XOR|1 I1|_XOR|2 JJMIT AREA=2.5
BI1|_XOR|2 I1|_XOR|4 I1|_XOR|5 JJMIT AREA=2.09
BI1|_XOR|3 I1|_XOR|25 I1|_XOR|6 JJMIT AREA=1.71
BI1|_XOR|4 I1|_XOR|9 I1|_XOR|10 JJMIT AREA=2.5
BI1|_XOR|5 I1|_XOR|12 I1|_XOR|13 JJMIT AREA=2.09
BI1|_XOR|6 I1|_XOR|26 I1|_XOR|14 JJMIT AREA=1.71
BI1|_XOR|7 I1|_XOR|27 I1|_XOR|16 JJMIT AREA=1.62
BI1|_XOR|8 I1|_XOR|17 I1|_XOR|18 JJMIT AREA=2.5
BI1|_XOR|9 I1|_XOR|20 I1|_XOR|16 JJMIT AREA=1.45
BI1|_XOR|10 I1|_XOR|16 I1|_XOR|21 JJMIT AREA=0.89
BI1|_XOR|11 I1|_XOR|22 I1|_XOR|23 JJMIT AREA=2.5
II1|_XOR|B1 0 I1|_XOR|3  PWL(0 0 5e-12 0.000175)
II1|_XOR|B2 0 I1|_XOR|7  PWL(0 0 5e-12 0.000112)
II1|_XOR|B3 0 I1|_XOR|11  PWL(0 0 5e-12 0.000175)
II1|_XOR|B4 0 I1|_XOR|15  PWL(0 0 5e-12 0.000112)
II1|_XOR|B5 0 I1|_XOR|19  PWL(0 0 5e-12 0.000175)
II1|_XOR|B6 0 I1|_XOR|24  PWL(0 0 5e-12 0.000175)
LI1|_XOR|B1 I1|_XOR|3 I1|_XOR|1  2e-12
LI1|_XOR|B2 I1|_XOR|7 I1|_XOR|6  2e-12
LI1|_XOR|B3 I1|_XOR|11 I1|_XOR|9  2e-12
LI1|_XOR|B4 I1|_XOR|15 I1|_XOR|14  2e-12
LI1|_XOR|B5 I1|_XOR|19 I1|_XOR|17  2e-12
LI1|_XOR|B6 I1|_XOR|24 I1|_XOR|22  2e-12
LI1|_XOR|1 I1|A2 I1|_XOR|1  2.06e-12
LI1|_XOR|2 I1|_XOR|1 I1|_XOR|4  3.233e-12
LI1|_XOR|3 I1|_XOR|4 I1|_XOR|25  1.419e-12
LI1|_XOR|4 I1|_XOR|6 I1|_XOR|8  6.051e-12
LI1|_XOR|5 I1|B2 I1|_XOR|9  2.092e-12
LI1|_XOR|6 I1|_XOR|9 I1|_XOR|12  3.221e-12
LI1|_XOR|7 I1|_XOR|12 I1|_XOR|26  1.384e-12
LI1|_XOR|8 I1|_XOR|14 I1|_XOR|8  6.059e-12
LI1|_XOR|9 I1|_XOR|8 I1|_XOR|27  1.301e-12
LI1|_XOR|10 T01 I1|_XOR|17  2.082e-12
LI1|_XOR|11 I1|_XOR|17 I1|_XOR|20  1.43e-12
LI1|_XOR|12 I1|_XOR|16 I1|_XOR|22  3.892e-12
LI1|_XOR|13 I1|_XOR|22 IP1_0  2.077e-12
LI1|_XOR|P1 I1|_XOR|2 0  5.508e-13
LI1|_XOR|P2 I1|_XOR|5 0  4.769e-13
LI1|_XOR|P4 I1|_XOR|10 0  4.767e-13
LI1|_XOR|P5 I1|_XOR|13 0  4.812e-13
LI1|_XOR|P8 I1|_XOR|18 0  4.526e-13
LI1|_XOR|P10 I1|_XOR|21 0  5.69e-13
LI1|_XOR|P11 I1|_XOR|23 0  4.746e-13
RI1|_XOR|B1 I1|_XOR|1 I1|_XOR|101  2.7439617672
LI1|_XOR|RB1 I1|_XOR|101 0  2.050338398468e-12
RI1|_XOR|B2 I1|_XOR|4 I1|_XOR|104  3.2822509177033496
LI1|_XOR|RB2 I1|_XOR|104 0  2.3544717685023925e-12
RI1|_XOR|B3 I1|_XOR|4 I1|_XOR|106  4.011640010526316
LI1|_XOR|RB3 I1|_XOR|106 I1|_XOR|6  2.766576605947368e-12
RI1|_XOR|B4 I1|_XOR|9 I1|_XOR|109  2.7439617672
LI1|_XOR|RB4 I1|_XOR|109 0  2.050338398468e-12
RI1|_XOR|B5 I1|_XOR|12 I1|_XOR|112  3.2822509177033496
LI1|_XOR|RB5 I1|_XOR|112 0  2.3544717685023925e-12
RI1|_XOR|B6 I1|_XOR|12 I1|_XOR|114  4.011640010526316
LI1|_XOR|RB6 I1|_XOR|114 I1|_XOR|14  2.766576605947368e-12
RI1|_XOR|B7 I1|_XOR|8 I1|_XOR|108  4.2345089
LI1|_XOR|RB7 I1|_XOR|108 I1|_XOR|16  2.8924975284999997e-12
RI1|_XOR|B8 I1|_XOR|17 I1|_XOR|117  2.7439617672
LI1|_XOR|RB8 I1|_XOR|117 0  2.050338398468e-12
RI1|_XOR|B9 I1|_XOR|20 I1|_XOR|120  4.730968564137931
LI1|_XOR|RB9 I1|_XOR|120 I1|_XOR|16  3.172997238737931e-12
RI1|_XOR|B10 I1|_XOR|16 I1|_XOR|116  7.707757773033708
LI1|_XOR|RB10 I1|_XOR|116 0  4.854883141764045e-12
RI1|_XOR|B11 I1|_XOR|22 I1|_XOR|122  2.7439617672
LI1|_XOR|RB11 I1|_XOR|122 0  2.050338398468e-12
LI1|_AND|A1 I1|A1_SYNC I1|_AND|A1  2.067833848e-12
LI1|_AND|A2 I1|_AND|A1 I1|_AND|A2  4.135667696e-12
LI1|_AND|A3 I1|_AND|A3 I1|_AND|Q3  1.2e-12
LI1|_AND|B1 I1|B1_SYNC I1|_AND|B1  2.067833848e-12
LI1|_AND|B2 I1|_AND|B1 I1|_AND|B2  4.135667696e-12
LI1|_AND|B3 I1|_AND|B3 I1|_AND|Q3  1.2e-12
LI1|_AND|Q3 I1|_AND|Q3 I1|_AND|Q2  4.135667696e-12
LI1|_AND|Q2 I1|_AND|Q2 I1|_AND|Q1  4.135667696e-12
LI1|_AND|Q1 I1|_AND|Q1 IG1_0  2.067833848e-12
II2|_SPL_A|B1 0 I2|_SPL_A|3  PWL(0 0 5e-12 0.000175)
II2|_SPL_A|B2 0 I2|_SPL_A|6  PWL(0 0 5e-12 0.00028)
II2|_SPL_A|B3 0 I2|_SPL_A|10  PWL(0 0 5e-12 0.000175)
II2|_SPL_A|B4 0 I2|_SPL_A|13  PWL(0 0 5e-12 0.000175)
LI2|_SPL_A|B1 I2|_SPL_A|3 I2|_SPL_A|1  9.175e-13
LI2|_SPL_A|B2 I2|_SPL_A|6 I2|_SPL_A|4  7.666e-13
LI2|_SPL_A|B3 I2|_SPL_A|10 I2|_SPL_A|8  1.928e-12
LI2|_SPL_A|B4 I2|_SPL_A|13 I2|_SPL_A|11  8.786e-13
BI2|_SPL_A|1 I2|_SPL_A|1 I2|_SPL_A|2 JJMIT AREA=2.5
BI2|_SPL_A|2 I2|_SPL_A|4 I2|_SPL_A|5 JJMIT AREA=3.0
BI2|_SPL_A|3 I2|_SPL_A|8 I2|_SPL_A|9 JJMIT AREA=2.5
BI2|_SPL_A|4 I2|_SPL_A|11 I2|_SPL_A|12 JJMIT AREA=2.5
LI2|_SPL_A|1 A2 I2|_SPL_A|1  2.063e-12
LI2|_SPL_A|2 I2|_SPL_A|1 I2|_SPL_A|4  3.637e-12
LI2|_SPL_A|3 I2|_SPL_A|4 I2|_SPL_A|7  1.278e-12
LI2|_SPL_A|4 I2|_SPL_A|7 I2|_SPL_A|8  1.305e-12
LI2|_SPL_A|5 I2|_SPL_A|8 I2|A1  2.05e-12
LI2|_SPL_A|6 I2|_SPL_A|7 I2|_SPL_A|11  1.315e-12
LI2|_SPL_A|7 I2|_SPL_A|11 I2|A2  2.06e-12
LI2|_SPL_A|P1 I2|_SPL_A|2 0  4.676e-13
LI2|_SPL_A|P2 I2|_SPL_A|5 0  4.498e-13
LI2|_SPL_A|P3 I2|_SPL_A|9 0  5.183e-13
LI2|_SPL_A|P4 I2|_SPL_A|12 0  4.639e-13
RI2|_SPL_A|B1 I2|_SPL_A|1 I2|_SPL_A|101  2.7439617672
LI2|_SPL_A|RB1 I2|_SPL_A|101 0  1.550338398468e-12
RI2|_SPL_A|B2 I2|_SPL_A|4 I2|_SPL_A|104  2.286634806
LI2|_SPL_A|RB2 I2|_SPL_A|104 0  1.29194866539e-12
RI2|_SPL_A|B3 I2|_SPL_A|8 I2|_SPL_A|108  2.7439617672
LI2|_SPL_A|RB3 I2|_SPL_A|108 0  1.550338398468e-12
RI2|_SPL_A|B4 I2|_SPL_A|11 I2|_SPL_A|111  2.7439617672
LI2|_SPL_A|RB4 I2|_SPL_A|111 0  1.550338398468e-12
II2|_SPL_B|B1 0 I2|_SPL_B|3  PWL(0 0 5e-12 0.000175)
II2|_SPL_B|B2 0 I2|_SPL_B|6  PWL(0 0 5e-12 0.00028)
II2|_SPL_B|B3 0 I2|_SPL_B|10  PWL(0 0 5e-12 0.000175)
II2|_SPL_B|B4 0 I2|_SPL_B|13  PWL(0 0 5e-12 0.000175)
LI2|_SPL_B|B1 I2|_SPL_B|3 I2|_SPL_B|1  9.175e-13
LI2|_SPL_B|B2 I2|_SPL_B|6 I2|_SPL_B|4  7.666e-13
LI2|_SPL_B|B3 I2|_SPL_B|10 I2|_SPL_B|8  1.928e-12
LI2|_SPL_B|B4 I2|_SPL_B|13 I2|_SPL_B|11  8.786e-13
BI2|_SPL_B|1 I2|_SPL_B|1 I2|_SPL_B|2 JJMIT AREA=2.5
BI2|_SPL_B|2 I2|_SPL_B|4 I2|_SPL_B|5 JJMIT AREA=3.0
BI2|_SPL_B|3 I2|_SPL_B|8 I2|_SPL_B|9 JJMIT AREA=2.5
BI2|_SPL_B|4 I2|_SPL_B|11 I2|_SPL_B|12 JJMIT AREA=2.5
LI2|_SPL_B|1 B2 I2|_SPL_B|1  2.063e-12
LI2|_SPL_B|2 I2|_SPL_B|1 I2|_SPL_B|4  3.637e-12
LI2|_SPL_B|3 I2|_SPL_B|4 I2|_SPL_B|7  1.278e-12
LI2|_SPL_B|4 I2|_SPL_B|7 I2|_SPL_B|8  1.305e-12
LI2|_SPL_B|5 I2|_SPL_B|8 I2|B1  2.05e-12
LI2|_SPL_B|6 I2|_SPL_B|7 I2|_SPL_B|11  1.315e-12
LI2|_SPL_B|7 I2|_SPL_B|11 I2|B2  2.06e-12
LI2|_SPL_B|P1 I2|_SPL_B|2 0  4.676e-13
LI2|_SPL_B|P2 I2|_SPL_B|5 0  4.498e-13
LI2|_SPL_B|P3 I2|_SPL_B|9 0  5.183e-13
LI2|_SPL_B|P4 I2|_SPL_B|12 0  4.639e-13
RI2|_SPL_B|B1 I2|_SPL_B|1 I2|_SPL_B|101  2.7439617672
LI2|_SPL_B|RB1 I2|_SPL_B|101 0  1.550338398468e-12
RI2|_SPL_B|B2 I2|_SPL_B|4 I2|_SPL_B|104  2.286634806
LI2|_SPL_B|RB2 I2|_SPL_B|104 0  1.29194866539e-12
RI2|_SPL_B|B3 I2|_SPL_B|8 I2|_SPL_B|108  2.7439617672
LI2|_SPL_B|RB3 I2|_SPL_B|108 0  1.550338398468e-12
RI2|_SPL_B|B4 I2|_SPL_B|11 I2|_SPL_B|111  2.7439617672
LI2|_SPL_B|RB4 I2|_SPL_B|111 0  1.550338398468e-12
BI2|_DFF_A|1 I2|_DFF_A|1 I2|_DFF_A|2 JJMIT AREA=2.5
BI2|_DFF_A|2 I2|_DFF_A|4 I2|_DFF_A|5 JJMIT AREA=1.61
BI2|_DFF_A|3 I2|_DFF_A|5 I2|_DFF_A|6 JJMIT AREA=1.54
BI2|_DFF_A|4 I2|_DFF_A|8 I2|_DFF_A|9 JJMIT AREA=1.69
BI2|_DFF_A|5 I2|_DFF_A|10 I2|_DFF_A|8 JJMIT AREA=1.38
BI2|_DFF_A|6 I2|_DFF_A|11 I2|_DFF_A|12 JJMIT AREA=2.5
BI2|_DFF_A|7 I2|_DFF_A|14 I2|_DFF_A|15 JJMIT AREA=2.5
II2|_DFF_A|B1 0 I2|_DFF_A|3  PWL(0 0 5e-12 0.000175)
II2|_DFF_A|B2 0 I2|_DFF_A|7  PWL(0 0 5e-12 0.000173)
II2|_DFF_A|B3 0 I2|_DFF_A|13  PWL(0 0 5e-12 0.000175)
II2|_DFF_A|B4 0 I2|_DFF_A|16  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|B1 I2|_DFF_A|3 I2|_DFF_A|1  2e-12
LI2|_DFF_A|B2 I2|_DFF_A|7 I2|_DFF_A|5  2e-12
LI2|_DFF_A|B3 I2|_DFF_A|11 I2|_DFF_A|13  2e-12
LI2|_DFF_A|B4 I2|_DFF_A|16 I2|_DFF_A|14  2e-12
LI2|_DFF_A|1 I2|A1 I2|_DFF_A|1  2.059e-12
LI2|_DFF_A|2 I2|_DFF_A|1 I2|_DFF_A|4  4.123e-12
LI2|_DFF_A|3 I2|_DFF_A|5 I2|_DFF_A|8  6.873e-12
LI2|_DFF_A|4 I2|_DFF_A|10 I2|_DFF_A|11  5.195e-12
LI2|_DFF_A|5 T02 I2|_DFF_A|11  2.071e-12
LI2|_DFF_A|6 I2|_DFF_A|8 I2|_DFF_A|14  3.287e-12
LI2|_DFF_A|7 I2|_DFF_A|14 I2|A1_SYNC  2.066e-12
LI2|_DFF_A|P1 I2|_DFF_A|2 0  5.042e-13
LI2|_DFF_A|P3 I2|_DFF_A|6 0  5.799e-13
LI2|_DFF_A|P4 I2|_DFF_A|9 0  5.733e-13
LI2|_DFF_A|P6 I2|_DFF_A|12 0  4.605e-13
LI2|_DFF_A|P7 I2|_DFF_A|15 0  4.961e-13
RI2|_DFF_A|B1 I2|_DFF_A|1 I2|_DFF_A|101  2.7439617672
LI2|_DFF_A|RB1 I2|_DFF_A|101 0  1.550338398468e-12
RI2|_DFF_A|B2 I2|_DFF_A|4 I2|_DFF_A|104  4.260810197515528
LI2|_DFF_A|RB2 I2|_DFF_A|104 I2|_DFF_A|5  2.407357761596273e-12
RI2|_DFF_A|B3 I2|_DFF_A|5 I2|_DFF_A|105  4.454483388311688
LI2|_DFF_A|RB3 I2|_DFF_A|105 0  2.516783114396104e-12
RI2|_DFF_A|B4 I2|_DFF_A|8 I2|_DFF_A|108  4.059115040236686
LI2|_DFF_A|RB4 I2|_DFF_A|108 0  2.2933999977337278e-12
RI2|_DFF_A|B5 I2|_DFF_A|10 I2|_DFF_A|110  4.970945230434783
LI2|_DFF_A|RB5 I2|_DFF_A|110 I2|_DFF_A|8  2.8085840551956523e-12
RI2|_DFF_A|B6 I2|_DFF_A|11 I2|_DFF_A|111  2.7439617672
LI2|_DFF_A|RB6 I2|_DFF_A|111 0  1.550338398468e-12
RI2|_DFF_A|B7 I2|_DFF_A|14 I2|_DFF_A|114  2.7439617672
LI2|_DFF_A|RB7 I2|_DFF_A|114 0  1.550338398468e-12
BI2|_DFF_B|1 I2|_DFF_B|1 I2|_DFF_B|2 JJMIT AREA=2.5
BI2|_DFF_B|2 I2|_DFF_B|4 I2|_DFF_B|5 JJMIT AREA=1.61
BI2|_DFF_B|3 I2|_DFF_B|5 I2|_DFF_B|6 JJMIT AREA=1.54
BI2|_DFF_B|4 I2|_DFF_B|8 I2|_DFF_B|9 JJMIT AREA=1.69
BI2|_DFF_B|5 I2|_DFF_B|10 I2|_DFF_B|8 JJMIT AREA=1.38
BI2|_DFF_B|6 I2|_DFF_B|11 I2|_DFF_B|12 JJMIT AREA=2.5
BI2|_DFF_B|7 I2|_DFF_B|14 I2|_DFF_B|15 JJMIT AREA=2.5
II2|_DFF_B|B1 0 I2|_DFF_B|3  PWL(0 0 5e-12 0.000175)
II2|_DFF_B|B2 0 I2|_DFF_B|7  PWL(0 0 5e-12 0.000173)
II2|_DFF_B|B3 0 I2|_DFF_B|13  PWL(0 0 5e-12 0.000175)
II2|_DFF_B|B4 0 I2|_DFF_B|16  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|B1 I2|_DFF_B|3 I2|_DFF_B|1  2e-12
LI2|_DFF_B|B2 I2|_DFF_B|7 I2|_DFF_B|5  2e-12
LI2|_DFF_B|B3 I2|_DFF_B|11 I2|_DFF_B|13  2e-12
LI2|_DFF_B|B4 I2|_DFF_B|16 I2|_DFF_B|14  2e-12
LI2|_DFF_B|1 I2|B1 I2|_DFF_B|1  2.059e-12
LI2|_DFF_B|2 I2|_DFF_B|1 I2|_DFF_B|4  4.123e-12
LI2|_DFF_B|3 I2|_DFF_B|5 I2|_DFF_B|8  6.873e-12
LI2|_DFF_B|4 I2|_DFF_B|10 I2|_DFF_B|11  5.195e-12
LI2|_DFF_B|5 T02 I2|_DFF_B|11  2.071e-12
LI2|_DFF_B|6 I2|_DFF_B|8 I2|_DFF_B|14  3.287e-12
LI2|_DFF_B|7 I2|_DFF_B|14 I2|B1_SYNC  2.066e-12
LI2|_DFF_B|P1 I2|_DFF_B|2 0  5.042e-13
LI2|_DFF_B|P3 I2|_DFF_B|6 0  5.799e-13
LI2|_DFF_B|P4 I2|_DFF_B|9 0  5.733e-13
LI2|_DFF_B|P6 I2|_DFF_B|12 0  4.605e-13
LI2|_DFF_B|P7 I2|_DFF_B|15 0  4.961e-13
RI2|_DFF_B|B1 I2|_DFF_B|1 I2|_DFF_B|101  2.7439617672
LI2|_DFF_B|RB1 I2|_DFF_B|101 0  1.550338398468e-12
RI2|_DFF_B|B2 I2|_DFF_B|4 I2|_DFF_B|104  4.260810197515528
LI2|_DFF_B|RB2 I2|_DFF_B|104 I2|_DFF_B|5  2.407357761596273e-12
RI2|_DFF_B|B3 I2|_DFF_B|5 I2|_DFF_B|105  4.454483388311688
LI2|_DFF_B|RB3 I2|_DFF_B|105 0  2.516783114396104e-12
RI2|_DFF_B|B4 I2|_DFF_B|8 I2|_DFF_B|108  4.059115040236686
LI2|_DFF_B|RB4 I2|_DFF_B|108 0  2.2933999977337278e-12
RI2|_DFF_B|B5 I2|_DFF_B|10 I2|_DFF_B|110  4.970945230434783
LI2|_DFF_B|RB5 I2|_DFF_B|110 I2|_DFF_B|8  2.8085840551956523e-12
RI2|_DFF_B|B6 I2|_DFF_B|11 I2|_DFF_B|111  2.7439617672
LI2|_DFF_B|RB6 I2|_DFF_B|111 0  1.550338398468e-12
RI2|_DFF_B|B7 I2|_DFF_B|14 I2|_DFF_B|114  2.7439617672
LI2|_DFF_B|RB7 I2|_DFF_B|114 0  1.550338398468e-12
BI2|_XOR|1 I2|_XOR|1 I2|_XOR|2 JJMIT AREA=2.5
BI2|_XOR|2 I2|_XOR|4 I2|_XOR|5 JJMIT AREA=2.09
BI2|_XOR|3 I2|_XOR|25 I2|_XOR|6 JJMIT AREA=1.71
BI2|_XOR|4 I2|_XOR|9 I2|_XOR|10 JJMIT AREA=2.5
BI2|_XOR|5 I2|_XOR|12 I2|_XOR|13 JJMIT AREA=2.09
BI2|_XOR|6 I2|_XOR|26 I2|_XOR|14 JJMIT AREA=1.71
BI2|_XOR|7 I2|_XOR|27 I2|_XOR|16 JJMIT AREA=1.62
BI2|_XOR|8 I2|_XOR|17 I2|_XOR|18 JJMIT AREA=2.5
BI2|_XOR|9 I2|_XOR|20 I2|_XOR|16 JJMIT AREA=1.45
BI2|_XOR|10 I2|_XOR|16 I2|_XOR|21 JJMIT AREA=0.89
BI2|_XOR|11 I2|_XOR|22 I2|_XOR|23 JJMIT AREA=2.5
II2|_XOR|B1 0 I2|_XOR|3  PWL(0 0 5e-12 0.000175)
II2|_XOR|B2 0 I2|_XOR|7  PWL(0 0 5e-12 0.000112)
II2|_XOR|B3 0 I2|_XOR|11  PWL(0 0 5e-12 0.000175)
II2|_XOR|B4 0 I2|_XOR|15  PWL(0 0 5e-12 0.000112)
II2|_XOR|B5 0 I2|_XOR|19  PWL(0 0 5e-12 0.000175)
II2|_XOR|B6 0 I2|_XOR|24  PWL(0 0 5e-12 0.000175)
LI2|_XOR|B1 I2|_XOR|3 I2|_XOR|1  2e-12
LI2|_XOR|B2 I2|_XOR|7 I2|_XOR|6  2e-12
LI2|_XOR|B3 I2|_XOR|11 I2|_XOR|9  2e-12
LI2|_XOR|B4 I2|_XOR|15 I2|_XOR|14  2e-12
LI2|_XOR|B5 I2|_XOR|19 I2|_XOR|17  2e-12
LI2|_XOR|B6 I2|_XOR|24 I2|_XOR|22  2e-12
LI2|_XOR|1 I2|A2 I2|_XOR|1  2.06e-12
LI2|_XOR|2 I2|_XOR|1 I2|_XOR|4  3.233e-12
LI2|_XOR|3 I2|_XOR|4 I2|_XOR|25  1.419e-12
LI2|_XOR|4 I2|_XOR|6 I2|_XOR|8  6.051e-12
LI2|_XOR|5 I2|B2 I2|_XOR|9  2.092e-12
LI2|_XOR|6 I2|_XOR|9 I2|_XOR|12  3.221e-12
LI2|_XOR|7 I2|_XOR|12 I2|_XOR|26  1.384e-12
LI2|_XOR|8 I2|_XOR|14 I2|_XOR|8  6.059e-12
LI2|_XOR|9 I2|_XOR|8 I2|_XOR|27  1.301e-12
LI2|_XOR|10 T02 I2|_XOR|17  2.082e-12
LI2|_XOR|11 I2|_XOR|17 I2|_XOR|20  1.43e-12
LI2|_XOR|12 I2|_XOR|16 I2|_XOR|22  3.892e-12
LI2|_XOR|13 I2|_XOR|22 IP2_0  2.077e-12
LI2|_XOR|P1 I2|_XOR|2 0  5.508e-13
LI2|_XOR|P2 I2|_XOR|5 0  4.769e-13
LI2|_XOR|P4 I2|_XOR|10 0  4.767e-13
LI2|_XOR|P5 I2|_XOR|13 0  4.812e-13
LI2|_XOR|P8 I2|_XOR|18 0  4.526e-13
LI2|_XOR|P10 I2|_XOR|21 0  5.69e-13
LI2|_XOR|P11 I2|_XOR|23 0  4.746e-13
RI2|_XOR|B1 I2|_XOR|1 I2|_XOR|101  2.7439617672
LI2|_XOR|RB1 I2|_XOR|101 0  2.050338398468e-12
RI2|_XOR|B2 I2|_XOR|4 I2|_XOR|104  3.2822509177033496
LI2|_XOR|RB2 I2|_XOR|104 0  2.3544717685023925e-12
RI2|_XOR|B3 I2|_XOR|4 I2|_XOR|106  4.011640010526316
LI2|_XOR|RB3 I2|_XOR|106 I2|_XOR|6  2.766576605947368e-12
RI2|_XOR|B4 I2|_XOR|9 I2|_XOR|109  2.7439617672
LI2|_XOR|RB4 I2|_XOR|109 0  2.050338398468e-12
RI2|_XOR|B5 I2|_XOR|12 I2|_XOR|112  3.2822509177033496
LI2|_XOR|RB5 I2|_XOR|112 0  2.3544717685023925e-12
RI2|_XOR|B6 I2|_XOR|12 I2|_XOR|114  4.011640010526316
LI2|_XOR|RB6 I2|_XOR|114 I2|_XOR|14  2.766576605947368e-12
RI2|_XOR|B7 I2|_XOR|8 I2|_XOR|108  4.2345089
LI2|_XOR|RB7 I2|_XOR|108 I2|_XOR|16  2.8924975284999997e-12
RI2|_XOR|B8 I2|_XOR|17 I2|_XOR|117  2.7439617672
LI2|_XOR|RB8 I2|_XOR|117 0  2.050338398468e-12
RI2|_XOR|B9 I2|_XOR|20 I2|_XOR|120  4.730968564137931
LI2|_XOR|RB9 I2|_XOR|120 I2|_XOR|16  3.172997238737931e-12
RI2|_XOR|B10 I2|_XOR|16 I2|_XOR|116  7.707757773033708
LI2|_XOR|RB10 I2|_XOR|116 0  4.854883141764045e-12
RI2|_XOR|B11 I2|_XOR|22 I2|_XOR|122  2.7439617672
LI2|_XOR|RB11 I2|_XOR|122 0  2.050338398468e-12
LI2|_AND|A1 I2|A1_SYNC I2|_AND|A1  2.067833848e-12
LI2|_AND|A2 I2|_AND|A1 I2|_AND|A2  4.135667696e-12
LI2|_AND|A3 I2|_AND|A3 I2|_AND|Q3  1.2e-12
LI2|_AND|B1 I2|B1_SYNC I2|_AND|B1  2.067833848e-12
LI2|_AND|B2 I2|_AND|B1 I2|_AND|B2  4.135667696e-12
LI2|_AND|B3 I2|_AND|B3 I2|_AND|Q3  1.2e-12
LI2|_AND|Q3 I2|_AND|Q3 I2|_AND|Q2  4.135667696e-12
LI2|_AND|Q2 I2|_AND|Q2 I2|_AND|Q1  4.135667696e-12
LI2|_AND|Q1 I2|_AND|Q1 IG2_0  2.067833848e-12
II3|_SPL_A|B1 0 I3|_SPL_A|3  PWL(0 0 5e-12 0.000175)
II3|_SPL_A|B2 0 I3|_SPL_A|6  PWL(0 0 5e-12 0.00028)
II3|_SPL_A|B3 0 I3|_SPL_A|10  PWL(0 0 5e-12 0.000175)
II3|_SPL_A|B4 0 I3|_SPL_A|13  PWL(0 0 5e-12 0.000175)
LI3|_SPL_A|B1 I3|_SPL_A|3 I3|_SPL_A|1  9.175e-13
LI3|_SPL_A|B2 I3|_SPL_A|6 I3|_SPL_A|4  7.666e-13
LI3|_SPL_A|B3 I3|_SPL_A|10 I3|_SPL_A|8  1.928e-12
LI3|_SPL_A|B4 I3|_SPL_A|13 I3|_SPL_A|11  8.786e-13
BI3|_SPL_A|1 I3|_SPL_A|1 I3|_SPL_A|2 JJMIT AREA=2.5
BI3|_SPL_A|2 I3|_SPL_A|4 I3|_SPL_A|5 JJMIT AREA=3.0
BI3|_SPL_A|3 I3|_SPL_A|8 I3|_SPL_A|9 JJMIT AREA=2.5
BI3|_SPL_A|4 I3|_SPL_A|11 I3|_SPL_A|12 JJMIT AREA=2.5
LI3|_SPL_A|1 A3 I3|_SPL_A|1  2.063e-12
LI3|_SPL_A|2 I3|_SPL_A|1 I3|_SPL_A|4  3.637e-12
LI3|_SPL_A|3 I3|_SPL_A|4 I3|_SPL_A|7  1.278e-12
LI3|_SPL_A|4 I3|_SPL_A|7 I3|_SPL_A|8  1.305e-12
LI3|_SPL_A|5 I3|_SPL_A|8 I3|A1  2.05e-12
LI3|_SPL_A|6 I3|_SPL_A|7 I3|_SPL_A|11  1.315e-12
LI3|_SPL_A|7 I3|_SPL_A|11 I3|A2  2.06e-12
LI3|_SPL_A|P1 I3|_SPL_A|2 0  4.676e-13
LI3|_SPL_A|P2 I3|_SPL_A|5 0  4.498e-13
LI3|_SPL_A|P3 I3|_SPL_A|9 0  5.183e-13
LI3|_SPL_A|P4 I3|_SPL_A|12 0  4.639e-13
RI3|_SPL_A|B1 I3|_SPL_A|1 I3|_SPL_A|101  2.7439617672
LI3|_SPL_A|RB1 I3|_SPL_A|101 0  1.550338398468e-12
RI3|_SPL_A|B2 I3|_SPL_A|4 I3|_SPL_A|104  2.286634806
LI3|_SPL_A|RB2 I3|_SPL_A|104 0  1.29194866539e-12
RI3|_SPL_A|B3 I3|_SPL_A|8 I3|_SPL_A|108  2.7439617672
LI3|_SPL_A|RB3 I3|_SPL_A|108 0  1.550338398468e-12
RI3|_SPL_A|B4 I3|_SPL_A|11 I3|_SPL_A|111  2.7439617672
LI3|_SPL_A|RB4 I3|_SPL_A|111 0  1.550338398468e-12
II3|_SPL_B|B1 0 I3|_SPL_B|3  PWL(0 0 5e-12 0.000175)
II3|_SPL_B|B2 0 I3|_SPL_B|6  PWL(0 0 5e-12 0.00028)
II3|_SPL_B|B3 0 I3|_SPL_B|10  PWL(0 0 5e-12 0.000175)
II3|_SPL_B|B4 0 I3|_SPL_B|13  PWL(0 0 5e-12 0.000175)
LI3|_SPL_B|B1 I3|_SPL_B|3 I3|_SPL_B|1  9.175e-13
LI3|_SPL_B|B2 I3|_SPL_B|6 I3|_SPL_B|4  7.666e-13
LI3|_SPL_B|B3 I3|_SPL_B|10 I3|_SPL_B|8  1.928e-12
LI3|_SPL_B|B4 I3|_SPL_B|13 I3|_SPL_B|11  8.786e-13
BI3|_SPL_B|1 I3|_SPL_B|1 I3|_SPL_B|2 JJMIT AREA=2.5
BI3|_SPL_B|2 I3|_SPL_B|4 I3|_SPL_B|5 JJMIT AREA=3.0
BI3|_SPL_B|3 I3|_SPL_B|8 I3|_SPL_B|9 JJMIT AREA=2.5
BI3|_SPL_B|4 I3|_SPL_B|11 I3|_SPL_B|12 JJMIT AREA=2.5
LI3|_SPL_B|1 B3 I3|_SPL_B|1  2.063e-12
LI3|_SPL_B|2 I3|_SPL_B|1 I3|_SPL_B|4  3.637e-12
LI3|_SPL_B|3 I3|_SPL_B|4 I3|_SPL_B|7  1.278e-12
LI3|_SPL_B|4 I3|_SPL_B|7 I3|_SPL_B|8  1.305e-12
LI3|_SPL_B|5 I3|_SPL_B|8 I3|B1  2.05e-12
LI3|_SPL_B|6 I3|_SPL_B|7 I3|_SPL_B|11  1.315e-12
LI3|_SPL_B|7 I3|_SPL_B|11 I3|B2  2.06e-12
LI3|_SPL_B|P1 I3|_SPL_B|2 0  4.676e-13
LI3|_SPL_B|P2 I3|_SPL_B|5 0  4.498e-13
LI3|_SPL_B|P3 I3|_SPL_B|9 0  5.183e-13
LI3|_SPL_B|P4 I3|_SPL_B|12 0  4.639e-13
RI3|_SPL_B|B1 I3|_SPL_B|1 I3|_SPL_B|101  2.7439617672
LI3|_SPL_B|RB1 I3|_SPL_B|101 0  1.550338398468e-12
RI3|_SPL_B|B2 I3|_SPL_B|4 I3|_SPL_B|104  2.286634806
LI3|_SPL_B|RB2 I3|_SPL_B|104 0  1.29194866539e-12
RI3|_SPL_B|B3 I3|_SPL_B|8 I3|_SPL_B|108  2.7439617672
LI3|_SPL_B|RB3 I3|_SPL_B|108 0  1.550338398468e-12
RI3|_SPL_B|B4 I3|_SPL_B|11 I3|_SPL_B|111  2.7439617672
LI3|_SPL_B|RB4 I3|_SPL_B|111 0  1.550338398468e-12
BI3|_DFF_A|1 I3|_DFF_A|1 I3|_DFF_A|2 JJMIT AREA=2.5
BI3|_DFF_A|2 I3|_DFF_A|4 I3|_DFF_A|5 JJMIT AREA=1.61
BI3|_DFF_A|3 I3|_DFF_A|5 I3|_DFF_A|6 JJMIT AREA=1.54
BI3|_DFF_A|4 I3|_DFF_A|8 I3|_DFF_A|9 JJMIT AREA=1.69
BI3|_DFF_A|5 I3|_DFF_A|10 I3|_DFF_A|8 JJMIT AREA=1.38
BI3|_DFF_A|6 I3|_DFF_A|11 I3|_DFF_A|12 JJMIT AREA=2.5
BI3|_DFF_A|7 I3|_DFF_A|14 I3|_DFF_A|15 JJMIT AREA=2.5
II3|_DFF_A|B1 0 I3|_DFF_A|3  PWL(0 0 5e-12 0.000175)
II3|_DFF_A|B2 0 I3|_DFF_A|7  PWL(0 0 5e-12 0.000173)
II3|_DFF_A|B3 0 I3|_DFF_A|13  PWL(0 0 5e-12 0.000175)
II3|_DFF_A|B4 0 I3|_DFF_A|16  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|B1 I3|_DFF_A|3 I3|_DFF_A|1  2e-12
LI3|_DFF_A|B2 I3|_DFF_A|7 I3|_DFF_A|5  2e-12
LI3|_DFF_A|B3 I3|_DFF_A|11 I3|_DFF_A|13  2e-12
LI3|_DFF_A|B4 I3|_DFF_A|16 I3|_DFF_A|14  2e-12
LI3|_DFF_A|1 I3|A1 I3|_DFF_A|1  2.059e-12
LI3|_DFF_A|2 I3|_DFF_A|1 I3|_DFF_A|4  4.123e-12
LI3|_DFF_A|3 I3|_DFF_A|5 I3|_DFF_A|8  6.873e-12
LI3|_DFF_A|4 I3|_DFF_A|10 I3|_DFF_A|11  5.195e-12
LI3|_DFF_A|5 T03 I3|_DFF_A|11  2.071e-12
LI3|_DFF_A|6 I3|_DFF_A|8 I3|_DFF_A|14  3.287e-12
LI3|_DFF_A|7 I3|_DFF_A|14 I3|A1_SYNC  2.066e-12
LI3|_DFF_A|P1 I3|_DFF_A|2 0  5.042e-13
LI3|_DFF_A|P3 I3|_DFF_A|6 0  5.799e-13
LI3|_DFF_A|P4 I3|_DFF_A|9 0  5.733e-13
LI3|_DFF_A|P6 I3|_DFF_A|12 0  4.605e-13
LI3|_DFF_A|P7 I3|_DFF_A|15 0  4.961e-13
RI3|_DFF_A|B1 I3|_DFF_A|1 I3|_DFF_A|101  2.7439617672
LI3|_DFF_A|RB1 I3|_DFF_A|101 0  1.550338398468e-12
RI3|_DFF_A|B2 I3|_DFF_A|4 I3|_DFF_A|104  4.260810197515528
LI3|_DFF_A|RB2 I3|_DFF_A|104 I3|_DFF_A|5  2.407357761596273e-12
RI3|_DFF_A|B3 I3|_DFF_A|5 I3|_DFF_A|105  4.454483388311688
LI3|_DFF_A|RB3 I3|_DFF_A|105 0  2.516783114396104e-12
RI3|_DFF_A|B4 I3|_DFF_A|8 I3|_DFF_A|108  4.059115040236686
LI3|_DFF_A|RB4 I3|_DFF_A|108 0  2.2933999977337278e-12
RI3|_DFF_A|B5 I3|_DFF_A|10 I3|_DFF_A|110  4.970945230434783
LI3|_DFF_A|RB5 I3|_DFF_A|110 I3|_DFF_A|8  2.8085840551956523e-12
RI3|_DFF_A|B6 I3|_DFF_A|11 I3|_DFF_A|111  2.7439617672
LI3|_DFF_A|RB6 I3|_DFF_A|111 0  1.550338398468e-12
RI3|_DFF_A|B7 I3|_DFF_A|14 I3|_DFF_A|114  2.7439617672
LI3|_DFF_A|RB7 I3|_DFF_A|114 0  1.550338398468e-12
BI3|_DFF_B|1 I3|_DFF_B|1 I3|_DFF_B|2 JJMIT AREA=2.5
BI3|_DFF_B|2 I3|_DFF_B|4 I3|_DFF_B|5 JJMIT AREA=1.61
BI3|_DFF_B|3 I3|_DFF_B|5 I3|_DFF_B|6 JJMIT AREA=1.54
BI3|_DFF_B|4 I3|_DFF_B|8 I3|_DFF_B|9 JJMIT AREA=1.69
BI3|_DFF_B|5 I3|_DFF_B|10 I3|_DFF_B|8 JJMIT AREA=1.38
BI3|_DFF_B|6 I3|_DFF_B|11 I3|_DFF_B|12 JJMIT AREA=2.5
BI3|_DFF_B|7 I3|_DFF_B|14 I3|_DFF_B|15 JJMIT AREA=2.5
II3|_DFF_B|B1 0 I3|_DFF_B|3  PWL(0 0 5e-12 0.000175)
II3|_DFF_B|B2 0 I3|_DFF_B|7  PWL(0 0 5e-12 0.000173)
II3|_DFF_B|B3 0 I3|_DFF_B|13  PWL(0 0 5e-12 0.000175)
II3|_DFF_B|B4 0 I3|_DFF_B|16  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|B1 I3|_DFF_B|3 I3|_DFF_B|1  2e-12
LI3|_DFF_B|B2 I3|_DFF_B|7 I3|_DFF_B|5  2e-12
LI3|_DFF_B|B3 I3|_DFF_B|11 I3|_DFF_B|13  2e-12
LI3|_DFF_B|B4 I3|_DFF_B|16 I3|_DFF_B|14  2e-12
LI3|_DFF_B|1 I3|B1 I3|_DFF_B|1  2.059e-12
LI3|_DFF_B|2 I3|_DFF_B|1 I3|_DFF_B|4  4.123e-12
LI3|_DFF_B|3 I3|_DFF_B|5 I3|_DFF_B|8  6.873e-12
LI3|_DFF_B|4 I3|_DFF_B|10 I3|_DFF_B|11  5.195e-12
LI3|_DFF_B|5 T03 I3|_DFF_B|11  2.071e-12
LI3|_DFF_B|6 I3|_DFF_B|8 I3|_DFF_B|14  3.287e-12
LI3|_DFF_B|7 I3|_DFF_B|14 I3|B1_SYNC  2.066e-12
LI3|_DFF_B|P1 I3|_DFF_B|2 0  5.042e-13
LI3|_DFF_B|P3 I3|_DFF_B|6 0  5.799e-13
LI3|_DFF_B|P4 I3|_DFF_B|9 0  5.733e-13
LI3|_DFF_B|P6 I3|_DFF_B|12 0  4.605e-13
LI3|_DFF_B|P7 I3|_DFF_B|15 0  4.961e-13
RI3|_DFF_B|B1 I3|_DFF_B|1 I3|_DFF_B|101  2.7439617672
LI3|_DFF_B|RB1 I3|_DFF_B|101 0  1.550338398468e-12
RI3|_DFF_B|B2 I3|_DFF_B|4 I3|_DFF_B|104  4.260810197515528
LI3|_DFF_B|RB2 I3|_DFF_B|104 I3|_DFF_B|5  2.407357761596273e-12
RI3|_DFF_B|B3 I3|_DFF_B|5 I3|_DFF_B|105  4.454483388311688
LI3|_DFF_B|RB3 I3|_DFF_B|105 0  2.516783114396104e-12
RI3|_DFF_B|B4 I3|_DFF_B|8 I3|_DFF_B|108  4.059115040236686
LI3|_DFF_B|RB4 I3|_DFF_B|108 0  2.2933999977337278e-12
RI3|_DFF_B|B5 I3|_DFF_B|10 I3|_DFF_B|110  4.970945230434783
LI3|_DFF_B|RB5 I3|_DFF_B|110 I3|_DFF_B|8  2.8085840551956523e-12
RI3|_DFF_B|B6 I3|_DFF_B|11 I3|_DFF_B|111  2.7439617672
LI3|_DFF_B|RB6 I3|_DFF_B|111 0  1.550338398468e-12
RI3|_DFF_B|B7 I3|_DFF_B|14 I3|_DFF_B|114  2.7439617672
LI3|_DFF_B|RB7 I3|_DFF_B|114 0  1.550338398468e-12
BI3|_XOR|1 I3|_XOR|1 I3|_XOR|2 JJMIT AREA=2.5
BI3|_XOR|2 I3|_XOR|4 I3|_XOR|5 JJMIT AREA=2.09
BI3|_XOR|3 I3|_XOR|25 I3|_XOR|6 JJMIT AREA=1.71
BI3|_XOR|4 I3|_XOR|9 I3|_XOR|10 JJMIT AREA=2.5
BI3|_XOR|5 I3|_XOR|12 I3|_XOR|13 JJMIT AREA=2.09
BI3|_XOR|6 I3|_XOR|26 I3|_XOR|14 JJMIT AREA=1.71
BI3|_XOR|7 I3|_XOR|27 I3|_XOR|16 JJMIT AREA=1.62
BI3|_XOR|8 I3|_XOR|17 I3|_XOR|18 JJMIT AREA=2.5
BI3|_XOR|9 I3|_XOR|20 I3|_XOR|16 JJMIT AREA=1.45
BI3|_XOR|10 I3|_XOR|16 I3|_XOR|21 JJMIT AREA=0.89
BI3|_XOR|11 I3|_XOR|22 I3|_XOR|23 JJMIT AREA=2.5
II3|_XOR|B1 0 I3|_XOR|3  PWL(0 0 5e-12 0.000175)
II3|_XOR|B2 0 I3|_XOR|7  PWL(0 0 5e-12 0.000112)
II3|_XOR|B3 0 I3|_XOR|11  PWL(0 0 5e-12 0.000175)
II3|_XOR|B4 0 I3|_XOR|15  PWL(0 0 5e-12 0.000112)
II3|_XOR|B5 0 I3|_XOR|19  PWL(0 0 5e-12 0.000175)
II3|_XOR|B6 0 I3|_XOR|24  PWL(0 0 5e-12 0.000175)
LI3|_XOR|B1 I3|_XOR|3 I3|_XOR|1  2e-12
LI3|_XOR|B2 I3|_XOR|7 I3|_XOR|6  2e-12
LI3|_XOR|B3 I3|_XOR|11 I3|_XOR|9  2e-12
LI3|_XOR|B4 I3|_XOR|15 I3|_XOR|14  2e-12
LI3|_XOR|B5 I3|_XOR|19 I3|_XOR|17  2e-12
LI3|_XOR|B6 I3|_XOR|24 I3|_XOR|22  2e-12
LI3|_XOR|1 I3|A2 I3|_XOR|1  2.06e-12
LI3|_XOR|2 I3|_XOR|1 I3|_XOR|4  3.233e-12
LI3|_XOR|3 I3|_XOR|4 I3|_XOR|25  1.419e-12
LI3|_XOR|4 I3|_XOR|6 I3|_XOR|8  6.051e-12
LI3|_XOR|5 I3|B2 I3|_XOR|9  2.092e-12
LI3|_XOR|6 I3|_XOR|9 I3|_XOR|12  3.221e-12
LI3|_XOR|7 I3|_XOR|12 I3|_XOR|26  1.384e-12
LI3|_XOR|8 I3|_XOR|14 I3|_XOR|8  6.059e-12
LI3|_XOR|9 I3|_XOR|8 I3|_XOR|27  1.301e-12
LI3|_XOR|10 T03 I3|_XOR|17  2.082e-12
LI3|_XOR|11 I3|_XOR|17 I3|_XOR|20  1.43e-12
LI3|_XOR|12 I3|_XOR|16 I3|_XOR|22  3.892e-12
LI3|_XOR|13 I3|_XOR|22 IP3_0  2.077e-12
LI3|_XOR|P1 I3|_XOR|2 0  5.508e-13
LI3|_XOR|P2 I3|_XOR|5 0  4.769e-13
LI3|_XOR|P4 I3|_XOR|10 0  4.767e-13
LI3|_XOR|P5 I3|_XOR|13 0  4.812e-13
LI3|_XOR|P8 I3|_XOR|18 0  4.526e-13
LI3|_XOR|P10 I3|_XOR|21 0  5.69e-13
LI3|_XOR|P11 I3|_XOR|23 0  4.746e-13
RI3|_XOR|B1 I3|_XOR|1 I3|_XOR|101  2.7439617672
LI3|_XOR|RB1 I3|_XOR|101 0  2.050338398468e-12
RI3|_XOR|B2 I3|_XOR|4 I3|_XOR|104  3.2822509177033496
LI3|_XOR|RB2 I3|_XOR|104 0  2.3544717685023925e-12
RI3|_XOR|B3 I3|_XOR|4 I3|_XOR|106  4.011640010526316
LI3|_XOR|RB3 I3|_XOR|106 I3|_XOR|6  2.766576605947368e-12
RI3|_XOR|B4 I3|_XOR|9 I3|_XOR|109  2.7439617672
LI3|_XOR|RB4 I3|_XOR|109 0  2.050338398468e-12
RI3|_XOR|B5 I3|_XOR|12 I3|_XOR|112  3.2822509177033496
LI3|_XOR|RB5 I3|_XOR|112 0  2.3544717685023925e-12
RI3|_XOR|B6 I3|_XOR|12 I3|_XOR|114  4.011640010526316
LI3|_XOR|RB6 I3|_XOR|114 I3|_XOR|14  2.766576605947368e-12
RI3|_XOR|B7 I3|_XOR|8 I3|_XOR|108  4.2345089
LI3|_XOR|RB7 I3|_XOR|108 I3|_XOR|16  2.8924975284999997e-12
RI3|_XOR|B8 I3|_XOR|17 I3|_XOR|117  2.7439617672
LI3|_XOR|RB8 I3|_XOR|117 0  2.050338398468e-12
RI3|_XOR|B9 I3|_XOR|20 I3|_XOR|120  4.730968564137931
LI3|_XOR|RB9 I3|_XOR|120 I3|_XOR|16  3.172997238737931e-12
RI3|_XOR|B10 I3|_XOR|16 I3|_XOR|116  7.707757773033708
LI3|_XOR|RB10 I3|_XOR|116 0  4.854883141764045e-12
RI3|_XOR|B11 I3|_XOR|22 I3|_XOR|122  2.7439617672
LI3|_XOR|RB11 I3|_XOR|122 0  2.050338398468e-12
LI3|_AND|A1 I3|A1_SYNC I3|_AND|A1  2.067833848e-12
LI3|_AND|A2 I3|_AND|A1 I3|_AND|A2  4.135667696e-12
LI3|_AND|A3 I3|_AND|A3 I3|_AND|Q3  1.2e-12
LI3|_AND|B1 I3|B1_SYNC I3|_AND|B1  2.067833848e-12
LI3|_AND|B2 I3|_AND|B1 I3|_AND|B2  4.135667696e-12
LI3|_AND|B3 I3|_AND|B3 I3|_AND|Q3  1.2e-12
LI3|_AND|Q3 I3|_AND|Q3 I3|_AND|Q2  4.135667696e-12
LI3|_AND|Q2 I3|_AND|Q2 I3|_AND|Q1  4.135667696e-12
LI3|_AND|Q1 I3|_AND|Q1 IG3_0  2.067833848e-12
B_PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP0_0|_TX|B1 0 _PTL_IP0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP0_0|_TX|B2 0 _PTL_IP0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|3  1.684e-12
L_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|6  3.596e-12
L_PTL_IP0_0|_TX|1 IP0_0 _PTL_IP0_0|_TX|1  2.063e-12
L_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|4  4.123e-12
L_PTL_IP0_0|_TX|3 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|7  2.193e-12
R_PTL_IP0_0|_TX|D _PTL_IP0_0|_TX|7 _PTL_IP0_0|A_PTL  1.36
L_PTL_IP0_0|_TX|P1 _PTL_IP0_0|_TX|2 0  5.254e-13
L_PTL_IP0_0|_TX|P2 _PTL_IP0_0|_TX|5 0  5.141e-13
R_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|101  2.7439617672
R_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|104  2.7439617672
L_PTL_IP0_0|_TX|RB1 _PTL_IP0_0|_TX|101 0  1.550338398468e-12
L_PTL_IP0_0|_TX|RB2 _PTL_IP0_0|_TX|104 0  1.550338398468e-12
B_PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP0_0|_RX|B1 0 _PTL_IP0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|3  2.777e-12
I_PTL_IP0_0|_RX|B2 0 _PTL_IP0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|6  2.685e-12
I_PTL_IP0_0|_RX|B3 0 _PTL_IP0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|9  2.764e-12
L_PTL_IP0_0|_RX|1 _PTL_IP0_0|A_PTL _PTL_IP0_0|_RX|1  1.346e-12
L_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|4  6.348e-12
L_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7  5.197e-12
L_PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7 IP0_0_RX  2.058e-12
L_PTL_IP0_0|_RX|P1 _PTL_IP0_0|_RX|2 0  4.795e-13
L_PTL_IP0_0|_RX|P2 _PTL_IP0_0|_RX|5 0  5.431e-13
L_PTL_IP0_0|_RX|P3 _PTL_IP0_0|_RX|8 0  5.339e-13
R_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|101  4.225701121488
R_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|104  3.429952209
R_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|107  2.7439617672
L_PTL_IP0_0|_RX|RB1 _PTL_IP0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP0_0|_RX|RB2 _PTL_IP0_0|_RX|104 0  1.937922998085e-12
L_PTL_IP0_0|_RX|RB3 _PTL_IP0_0|_RX|107 0  1.550338398468e-12
B_PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG0_0|_TX|B1 0 _PTL_IG0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG0_0|_TX|B2 0 _PTL_IG0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|3  1.684e-12
L_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|6  3.596e-12
L_PTL_IG0_0|_TX|1 IG0_0 _PTL_IG0_0|_TX|1  2.063e-12
L_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|4  4.123e-12
L_PTL_IG0_0|_TX|3 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|7  2.193e-12
R_PTL_IG0_0|_TX|D _PTL_IG0_0|_TX|7 _PTL_IG0_0|A_PTL  1.36
L_PTL_IG0_0|_TX|P1 _PTL_IG0_0|_TX|2 0  5.254e-13
L_PTL_IG0_0|_TX|P2 _PTL_IG0_0|_TX|5 0  5.141e-13
R_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|101  2.7439617672
R_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|104  2.7439617672
L_PTL_IG0_0|_TX|RB1 _PTL_IG0_0|_TX|101 0  1.550338398468e-12
L_PTL_IG0_0|_TX|RB2 _PTL_IG0_0|_TX|104 0  1.550338398468e-12
B_PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG0_0|_RX|B1 0 _PTL_IG0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|3  2.777e-12
I_PTL_IG0_0|_RX|B2 0 _PTL_IG0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|6  2.685e-12
I_PTL_IG0_0|_RX|B3 0 _PTL_IG0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|9  2.764e-12
L_PTL_IG0_0|_RX|1 _PTL_IG0_0|A_PTL _PTL_IG0_0|_RX|1  1.346e-12
L_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|4  6.348e-12
L_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7  5.197e-12
L_PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7 IG0_0_RX  2.058e-12
L_PTL_IG0_0|_RX|P1 _PTL_IG0_0|_RX|2 0  4.795e-13
L_PTL_IG0_0|_RX|P2 _PTL_IG0_0|_RX|5 0  5.431e-13
L_PTL_IG0_0|_RX|P3 _PTL_IG0_0|_RX|8 0  5.339e-13
R_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|101  4.225701121488
R_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|104  3.429952209
R_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|107  2.7439617672
L_PTL_IG0_0|_RX|RB1 _PTL_IG0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG0_0|_RX|RB2 _PTL_IG0_0|_RX|104 0  1.937922998085e-12
L_PTL_IG0_0|_RX|RB3 _PTL_IG0_0|_RX|107 0  1.550338398468e-12
B_PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_0|_TX|B1 0 _PTL_IP1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_0|_TX|B2 0 _PTL_IP1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|3  1.684e-12
L_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|6  3.596e-12
L_PTL_IP1_0|_TX|1 IP1_0 _PTL_IP1_0|_TX|1  2.063e-12
L_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|4  4.123e-12
L_PTL_IP1_0|_TX|3 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|7  2.193e-12
R_PTL_IP1_0|_TX|D _PTL_IP1_0|_TX|7 _PTL_IP1_0|A_PTL  1.36
L_PTL_IP1_0|_TX|P1 _PTL_IP1_0|_TX|2 0  5.254e-13
L_PTL_IP1_0|_TX|P2 _PTL_IP1_0|_TX|5 0  5.141e-13
R_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|101  2.7439617672
R_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|104  2.7439617672
L_PTL_IP1_0|_TX|RB1 _PTL_IP1_0|_TX|101 0  1.550338398468e-12
L_PTL_IP1_0|_TX|RB2 _PTL_IP1_0|_TX|104 0  1.550338398468e-12
B_PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_0|_RX|B1 0 _PTL_IP1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|3  2.777e-12
I_PTL_IP1_0|_RX|B2 0 _PTL_IP1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|6  2.685e-12
I_PTL_IP1_0|_RX|B3 0 _PTL_IP1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|9  2.764e-12
L_PTL_IP1_0|_RX|1 _PTL_IP1_0|A_PTL _PTL_IP1_0|_RX|1  1.346e-12
L_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|4  6.348e-12
L_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7  5.197e-12
L_PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7 IP1_0_RX  2.058e-12
L_PTL_IP1_0|_RX|P1 _PTL_IP1_0|_RX|2 0  4.795e-13
L_PTL_IP1_0|_RX|P2 _PTL_IP1_0|_RX|5 0  5.431e-13
L_PTL_IP1_0|_RX|P3 _PTL_IP1_0|_RX|8 0  5.339e-13
R_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|101  4.225701121488
R_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|104  3.429952209
R_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|107  2.7439617672
L_PTL_IP1_0|_RX|RB1 _PTL_IP1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_0|_RX|RB2 _PTL_IP1_0|_RX|104 0  1.937922998085e-12
L_PTL_IP1_0|_RX|RB3 _PTL_IP1_0|_RX|107 0  1.550338398468e-12
B_PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG1_0|_TX|B1 0 _PTL_IG1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG1_0|_TX|B2 0 _PTL_IG1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|3  1.684e-12
L_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|6  3.596e-12
L_PTL_IG1_0|_TX|1 IG1_0 _PTL_IG1_0|_TX|1  2.063e-12
L_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|4  4.123e-12
L_PTL_IG1_0|_TX|3 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|7  2.193e-12
R_PTL_IG1_0|_TX|D _PTL_IG1_0|_TX|7 _PTL_IG1_0|A_PTL  1.36
L_PTL_IG1_0|_TX|P1 _PTL_IG1_0|_TX|2 0  5.254e-13
L_PTL_IG1_0|_TX|P2 _PTL_IG1_0|_TX|5 0  5.141e-13
R_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|101  2.7439617672
R_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|104  2.7439617672
L_PTL_IG1_0|_TX|RB1 _PTL_IG1_0|_TX|101 0  1.550338398468e-12
L_PTL_IG1_0|_TX|RB2 _PTL_IG1_0|_TX|104 0  1.550338398468e-12
B_PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG1_0|_RX|B1 0 _PTL_IG1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|3  2.777e-12
I_PTL_IG1_0|_RX|B2 0 _PTL_IG1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|6  2.685e-12
I_PTL_IG1_0|_RX|B3 0 _PTL_IG1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|9  2.764e-12
L_PTL_IG1_0|_RX|1 _PTL_IG1_0|A_PTL _PTL_IG1_0|_RX|1  1.346e-12
L_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|4  6.348e-12
L_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7  5.197e-12
L_PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7 IG1_0_RX  2.058e-12
L_PTL_IG1_0|_RX|P1 _PTL_IG1_0|_RX|2 0  4.795e-13
L_PTL_IG1_0|_RX|P2 _PTL_IG1_0|_RX|5 0  5.431e-13
L_PTL_IG1_0|_RX|P3 _PTL_IG1_0|_RX|8 0  5.339e-13
R_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|101  4.225701121488
R_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|104  3.429952209
R_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|107  2.7439617672
L_PTL_IG1_0|_RX|RB1 _PTL_IG1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG1_0|_RX|RB2 _PTL_IG1_0|_RX|104 0  1.937922998085e-12
L_PTL_IG1_0|_RX|RB3 _PTL_IG1_0|_RX|107 0  1.550338398468e-12
B_PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_0|_TX|B1 0 _PTL_IP2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_0|_TX|B2 0 _PTL_IP2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|3  1.684e-12
L_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|6  3.596e-12
L_PTL_IP2_0|_TX|1 IP2_0 _PTL_IP2_0|_TX|1  2.063e-12
L_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|4  4.123e-12
L_PTL_IP2_0|_TX|3 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|7  2.193e-12
R_PTL_IP2_0|_TX|D _PTL_IP2_0|_TX|7 _PTL_IP2_0|A_PTL  1.36
L_PTL_IP2_0|_TX|P1 _PTL_IP2_0|_TX|2 0  5.254e-13
L_PTL_IP2_0|_TX|P2 _PTL_IP2_0|_TX|5 0  5.141e-13
R_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|101  2.7439617672
R_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|104  2.7439617672
L_PTL_IP2_0|_TX|RB1 _PTL_IP2_0|_TX|101 0  1.550338398468e-12
L_PTL_IP2_0|_TX|RB2 _PTL_IP2_0|_TX|104 0  1.550338398468e-12
B_PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_0|_RX|B1 0 _PTL_IP2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|3  2.777e-12
I_PTL_IP2_0|_RX|B2 0 _PTL_IP2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|6  2.685e-12
I_PTL_IP2_0|_RX|B3 0 _PTL_IP2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|9  2.764e-12
L_PTL_IP2_0|_RX|1 _PTL_IP2_0|A_PTL _PTL_IP2_0|_RX|1  1.346e-12
L_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|4  6.348e-12
L_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7  5.197e-12
L_PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7 IP2_0_RX  2.058e-12
L_PTL_IP2_0|_RX|P1 _PTL_IP2_0|_RX|2 0  4.795e-13
L_PTL_IP2_0|_RX|P2 _PTL_IP2_0|_RX|5 0  5.431e-13
L_PTL_IP2_0|_RX|P3 _PTL_IP2_0|_RX|8 0  5.339e-13
R_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|101  4.225701121488
R_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|104  3.429952209
R_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|107  2.7439617672
L_PTL_IP2_0|_RX|RB1 _PTL_IP2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_0|_RX|RB2 _PTL_IP2_0|_RX|104 0  1.937922998085e-12
L_PTL_IP2_0|_RX|RB3 _PTL_IP2_0|_RX|107 0  1.550338398468e-12
B_PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG2_0|_TX|B1 0 _PTL_IG2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG2_0|_TX|B2 0 _PTL_IG2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|3  1.684e-12
L_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|6  3.596e-12
L_PTL_IG2_0|_TX|1 IG2_0 _PTL_IG2_0|_TX|1  2.063e-12
L_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|4  4.123e-12
L_PTL_IG2_0|_TX|3 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|7  2.193e-12
R_PTL_IG2_0|_TX|D _PTL_IG2_0|_TX|7 _PTL_IG2_0|A_PTL  1.36
L_PTL_IG2_0|_TX|P1 _PTL_IG2_0|_TX|2 0  5.254e-13
L_PTL_IG2_0|_TX|P2 _PTL_IG2_0|_TX|5 0  5.141e-13
R_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|101  2.7439617672
R_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|104  2.7439617672
L_PTL_IG2_0|_TX|RB1 _PTL_IG2_0|_TX|101 0  1.550338398468e-12
L_PTL_IG2_0|_TX|RB2 _PTL_IG2_0|_TX|104 0  1.550338398468e-12
B_PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG2_0|_RX|B1 0 _PTL_IG2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|3  2.777e-12
I_PTL_IG2_0|_RX|B2 0 _PTL_IG2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|6  2.685e-12
I_PTL_IG2_0|_RX|B3 0 _PTL_IG2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|9  2.764e-12
L_PTL_IG2_0|_RX|1 _PTL_IG2_0|A_PTL _PTL_IG2_0|_RX|1  1.346e-12
L_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|4  6.348e-12
L_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7  5.197e-12
L_PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7 IG2_0_RX  2.058e-12
L_PTL_IG2_0|_RX|P1 _PTL_IG2_0|_RX|2 0  4.795e-13
L_PTL_IG2_0|_RX|P2 _PTL_IG2_0|_RX|5 0  5.431e-13
L_PTL_IG2_0|_RX|P3 _PTL_IG2_0|_RX|8 0  5.339e-13
R_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|101  4.225701121488
R_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|104  3.429952209
R_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|107  2.7439617672
L_PTL_IG2_0|_RX|RB1 _PTL_IG2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG2_0|_RX|RB2 _PTL_IG2_0|_RX|104 0  1.937922998085e-12
L_PTL_IG2_0|_RX|RB3 _PTL_IG2_0|_RX|107 0  1.550338398468e-12
B_PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_0|_TX|B1 0 _PTL_IP3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_0|_TX|B2 0 _PTL_IP3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|3  1.684e-12
L_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|6  3.596e-12
L_PTL_IP3_0|_TX|1 IP3_0 _PTL_IP3_0|_TX|1  2.063e-12
L_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|4  4.123e-12
L_PTL_IP3_0|_TX|3 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|7  2.193e-12
R_PTL_IP3_0|_TX|D _PTL_IP3_0|_TX|7 _PTL_IP3_0|A_PTL  1.36
L_PTL_IP3_0|_TX|P1 _PTL_IP3_0|_TX|2 0  5.254e-13
L_PTL_IP3_0|_TX|P2 _PTL_IP3_0|_TX|5 0  5.141e-13
R_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|101  2.7439617672
R_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|104  2.7439617672
L_PTL_IP3_0|_TX|RB1 _PTL_IP3_0|_TX|101 0  1.550338398468e-12
L_PTL_IP3_0|_TX|RB2 _PTL_IP3_0|_TX|104 0  1.550338398468e-12
B_PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_0|_RX|B1 0 _PTL_IP3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|3  2.777e-12
I_PTL_IP3_0|_RX|B2 0 _PTL_IP3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|6  2.685e-12
I_PTL_IP3_0|_RX|B3 0 _PTL_IP3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|9  2.764e-12
L_PTL_IP3_0|_RX|1 _PTL_IP3_0|A_PTL _PTL_IP3_0|_RX|1  1.346e-12
L_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|4  6.348e-12
L_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7  5.197e-12
L_PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7 IP3_0_RX  2.058e-12
L_PTL_IP3_0|_RX|P1 _PTL_IP3_0|_RX|2 0  4.795e-13
L_PTL_IP3_0|_RX|P2 _PTL_IP3_0|_RX|5 0  5.431e-13
L_PTL_IP3_0|_RX|P3 _PTL_IP3_0|_RX|8 0  5.339e-13
R_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|101  4.225701121488
R_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|104  3.429952209
R_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|107  2.7439617672
L_PTL_IP3_0|_RX|RB1 _PTL_IP3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_0|_RX|RB2 _PTL_IP3_0|_RX|104 0  1.937922998085e-12
L_PTL_IP3_0|_RX|RB3 _PTL_IP3_0|_RX|107 0  1.550338398468e-12
B_PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG3_0|_TX|B1 0 _PTL_IG3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG3_0|_TX|B2 0 _PTL_IG3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|3  1.684e-12
L_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|6  3.596e-12
L_PTL_IG3_0|_TX|1 IG3_0 _PTL_IG3_0|_TX|1  2.063e-12
L_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|4  4.123e-12
L_PTL_IG3_0|_TX|3 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|7  2.193e-12
R_PTL_IG3_0|_TX|D _PTL_IG3_0|_TX|7 _PTL_IG3_0|A_PTL  1.36
L_PTL_IG3_0|_TX|P1 _PTL_IG3_0|_TX|2 0  5.254e-13
L_PTL_IG3_0|_TX|P2 _PTL_IG3_0|_TX|5 0  5.141e-13
R_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|101  2.7439617672
R_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|104  2.7439617672
L_PTL_IG3_0|_TX|RB1 _PTL_IG3_0|_TX|101 0  1.550338398468e-12
L_PTL_IG3_0|_TX|RB2 _PTL_IG3_0|_TX|104 0  1.550338398468e-12
B_PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG3_0|_RX|B1 0 _PTL_IG3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|3  2.777e-12
I_PTL_IG3_0|_RX|B2 0 _PTL_IG3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|6  2.685e-12
I_PTL_IG3_0|_RX|B3 0 _PTL_IG3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|9  2.764e-12
L_PTL_IG3_0|_RX|1 _PTL_IG3_0|A_PTL _PTL_IG3_0|_RX|1  1.346e-12
L_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|4  6.348e-12
L_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7  5.197e-12
L_PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7 IG3_0_RX  2.058e-12
L_PTL_IG3_0|_RX|P1 _PTL_IG3_0|_RX|2 0  4.795e-13
L_PTL_IG3_0|_RX|P2 _PTL_IG3_0|_RX|5 0  5.431e-13
L_PTL_IG3_0|_RX|P3 _PTL_IG3_0|_RX|8 0  5.339e-13
R_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|101  4.225701121488
R_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|104  3.429952209
R_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|107  2.7439617672
L_PTL_IG3_0|_RX|RB1 _PTL_IG3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG3_0|_RX|RB2 _PTL_IG3_0|_RX|104 0  1.937922998085e-12
L_PTL_IG3_0|_RX|RB3 _PTL_IG3_0|_RX|107 0  1.550338398468e-12
LSPL_IP2_0|SPL1|1 IP2_0_RX SPL_IP2_0|SPL1|D1  2e-12
LSPL_IP2_0|SPL1|2 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|D2  4.135667696e-12
LSPL_IP2_0|SPL1|3 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL1|4 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL1|5 SPL_IP2_0|SPL1|QA1 IP2_0_TO2  2e-12
LSPL_IP2_0|SPL1|6 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL1|7 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|QTMP  2e-12
LSPL_IP2_0|SPL2|1 SPL_IP2_0|QTMP SPL_IP2_0|SPL2|D1  2e-12
LSPL_IP2_0|SPL2|2 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|D2  4.135667696e-12
LSPL_IP2_0|SPL2|3 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL2|4 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL2|5 SPL_IP2_0|SPL2|QA1 IP2_0_TO3  2e-12
LSPL_IP2_0|SPL2|6 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL2|7 SPL_IP2_0|SPL2|QB1 IP2_0_OUT  2e-12
B_PG0_01|P|1 _PG0_01|P|1 _PG0_01|P|2 JJMIT AREA=2.5
B_PG0_01|P|2 _PG0_01|P|4 _PG0_01|P|5 JJMIT AREA=1.61
B_PG0_01|P|3 _PG0_01|P|5 _PG0_01|P|6 JJMIT AREA=1.54
B_PG0_01|P|4 _PG0_01|P|8 _PG0_01|P|9 JJMIT AREA=1.69
B_PG0_01|P|5 _PG0_01|P|10 _PG0_01|P|8 JJMIT AREA=1.38
B_PG0_01|P|6 _PG0_01|P|11 _PG0_01|P|12 JJMIT AREA=2.5
B_PG0_01|P|7 _PG0_01|P|14 _PG0_01|P|15 JJMIT AREA=2.5
I_PG0_01|P|B1 0 _PG0_01|P|3  PWL(0 0 5e-12 0.000175)
I_PG0_01|P|B2 0 _PG0_01|P|7  PWL(0 0 5e-12 0.000173)
I_PG0_01|P|B3 0 _PG0_01|P|13  PWL(0 0 5e-12 0.000175)
I_PG0_01|P|B4 0 _PG0_01|P|16  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|B1 _PG0_01|P|3 _PG0_01|P|1  2e-12
L_PG0_01|P|B2 _PG0_01|P|7 _PG0_01|P|5  2e-12
L_PG0_01|P|B3 _PG0_01|P|11 _PG0_01|P|13  2e-12
L_PG0_01|P|B4 _PG0_01|P|16 _PG0_01|P|14  2e-12
L_PG0_01|P|1 IP0_0_RX _PG0_01|P|1  2.059e-12
L_PG0_01|P|2 _PG0_01|P|1 _PG0_01|P|4  4.123e-12
L_PG0_01|P|3 _PG0_01|P|5 _PG0_01|P|8  6.873e-12
L_PG0_01|P|4 _PG0_01|P|10 _PG0_01|P|11  5.195e-12
L_PG0_01|P|5 T04 _PG0_01|P|11  2.071e-12
L_PG0_01|P|6 _PG0_01|P|8 _PG0_01|P|14  3.287e-12
L_PG0_01|P|7 _PG0_01|P|14 P0_1  2.066e-12
L_PG0_01|P|P1 _PG0_01|P|2 0  5.042e-13
L_PG0_01|P|P3 _PG0_01|P|6 0  5.799e-13
L_PG0_01|P|P4 _PG0_01|P|9 0  5.733e-13
L_PG0_01|P|P6 _PG0_01|P|12 0  4.605e-13
L_PG0_01|P|P7 _PG0_01|P|15 0  4.961e-13
R_PG0_01|P|B1 _PG0_01|P|1 _PG0_01|P|101  2.7439617672
L_PG0_01|P|RB1 _PG0_01|P|101 0  1.550338398468e-12
R_PG0_01|P|B2 _PG0_01|P|4 _PG0_01|P|104  4.260810197515528
L_PG0_01|P|RB2 _PG0_01|P|104 _PG0_01|P|5  2.407357761596273e-12
R_PG0_01|P|B3 _PG0_01|P|5 _PG0_01|P|105  4.454483388311688
L_PG0_01|P|RB3 _PG0_01|P|105 0  2.516783114396104e-12
R_PG0_01|P|B4 _PG0_01|P|8 _PG0_01|P|108  4.059115040236686
L_PG0_01|P|RB4 _PG0_01|P|108 0  2.2933999977337278e-12
R_PG0_01|P|B5 _PG0_01|P|10 _PG0_01|P|110  4.970945230434783
L_PG0_01|P|RB5 _PG0_01|P|110 _PG0_01|P|8  2.8085840551956523e-12
R_PG0_01|P|B6 _PG0_01|P|11 _PG0_01|P|111  2.7439617672
L_PG0_01|P|RB6 _PG0_01|P|111 0  1.550338398468e-12
R_PG0_01|P|B7 _PG0_01|P|14 _PG0_01|P|114  2.7439617672
L_PG0_01|P|RB7 _PG0_01|P|114 0  1.550338398468e-12
B_PG0_01|G|1 _PG0_01|G|1 _PG0_01|G|2 JJMIT AREA=2.5
B_PG0_01|G|2 _PG0_01|G|4 _PG0_01|G|5 JJMIT AREA=1.61
B_PG0_01|G|3 _PG0_01|G|5 _PG0_01|G|6 JJMIT AREA=1.54
B_PG0_01|G|4 _PG0_01|G|8 _PG0_01|G|9 JJMIT AREA=1.69
B_PG0_01|G|5 _PG0_01|G|10 _PG0_01|G|8 JJMIT AREA=1.38
B_PG0_01|G|6 _PG0_01|G|11 _PG0_01|G|12 JJMIT AREA=2.5
B_PG0_01|G|7 _PG0_01|G|14 _PG0_01|G|15 JJMIT AREA=2.5
I_PG0_01|G|B1 0 _PG0_01|G|3  PWL(0 0 5e-12 0.000175)
I_PG0_01|G|B2 0 _PG0_01|G|7  PWL(0 0 5e-12 0.000173)
I_PG0_01|G|B3 0 _PG0_01|G|13  PWL(0 0 5e-12 0.000175)
I_PG0_01|G|B4 0 _PG0_01|G|16  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|B1 _PG0_01|G|3 _PG0_01|G|1  2e-12
L_PG0_01|G|B2 _PG0_01|G|7 _PG0_01|G|5  2e-12
L_PG0_01|G|B3 _PG0_01|G|11 _PG0_01|G|13  2e-12
L_PG0_01|G|B4 _PG0_01|G|16 _PG0_01|G|14  2e-12
L_PG0_01|G|1 IG0_0_TO0 _PG0_01|G|1  2.059e-12
L_PG0_01|G|2 _PG0_01|G|1 _PG0_01|G|4  4.123e-12
L_PG0_01|G|3 _PG0_01|G|5 _PG0_01|G|8  6.873e-12
L_PG0_01|G|4 _PG0_01|G|10 _PG0_01|G|11  5.195e-12
L_PG0_01|G|5 T04 _PG0_01|G|11  2.071e-12
L_PG0_01|G|6 _PG0_01|G|8 _PG0_01|G|14  3.287e-12
L_PG0_01|G|7 _PG0_01|G|14 G0_1  2.066e-12
L_PG0_01|G|P1 _PG0_01|G|2 0  5.042e-13
L_PG0_01|G|P3 _PG0_01|G|6 0  5.799e-13
L_PG0_01|G|P4 _PG0_01|G|9 0  5.733e-13
L_PG0_01|G|P6 _PG0_01|G|12 0  4.605e-13
L_PG0_01|G|P7 _PG0_01|G|15 0  4.961e-13
R_PG0_01|G|B1 _PG0_01|G|1 _PG0_01|G|101  2.7439617672
L_PG0_01|G|RB1 _PG0_01|G|101 0  1.550338398468e-12
R_PG0_01|G|B2 _PG0_01|G|4 _PG0_01|G|104  4.260810197515528
L_PG0_01|G|RB2 _PG0_01|G|104 _PG0_01|G|5  2.407357761596273e-12
R_PG0_01|G|B3 _PG0_01|G|5 _PG0_01|G|105  4.454483388311688
L_PG0_01|G|RB3 _PG0_01|G|105 0  2.516783114396104e-12
R_PG0_01|G|B4 _PG0_01|G|8 _PG0_01|G|108  4.059115040236686
L_PG0_01|G|RB4 _PG0_01|G|108 0  2.2933999977337278e-12
R_PG0_01|G|B5 _PG0_01|G|10 _PG0_01|G|110  4.970945230434783
L_PG0_01|G|RB5 _PG0_01|G|110 _PG0_01|G|8  2.8085840551956523e-12
R_PG0_01|G|B6 _PG0_01|G|11 _PG0_01|G|111  2.7439617672
L_PG0_01|G|RB6 _PG0_01|G|111 0  1.550338398468e-12
R_PG0_01|G|B7 _PG0_01|G|14 _PG0_01|G|114  2.7439617672
L_PG0_01|G|RB7 _PG0_01|G|114 0  1.550338398468e-12
I_PG1_01|_SPL_G1|B1 0 _PG1_01|_SPL_G1|3  PWL(0 0 5e-12 0.000175)
I_PG1_01|_SPL_G1|B2 0 _PG1_01|_SPL_G1|6  PWL(0 0 5e-12 0.00028)
I_PG1_01|_SPL_G1|B3 0 _PG1_01|_SPL_G1|10  PWL(0 0 5e-12 0.000175)
I_PG1_01|_SPL_G1|B4 0 _PG1_01|_SPL_G1|13  PWL(0 0 5e-12 0.000175)
L_PG1_01|_SPL_G1|B1 _PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|1  9.175e-13
L_PG1_01|_SPL_G1|B2 _PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|4  7.666e-13
L_PG1_01|_SPL_G1|B3 _PG1_01|_SPL_G1|10 _PG1_01|_SPL_G1|8  1.928e-12
L_PG1_01|_SPL_G1|B4 _PG1_01|_SPL_G1|13 _PG1_01|_SPL_G1|11  8.786e-13
B_PG1_01|_SPL_G1|1 _PG1_01|_SPL_G1|1 _PG1_01|_SPL_G1|2 JJMIT AREA=2.5
B_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|5 JJMIT AREA=3.0
B_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|8 _PG1_01|_SPL_G1|9 JJMIT AREA=2.5
B_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|11 _PG1_01|_SPL_G1|12 JJMIT AREA=2.5
L_PG1_01|_SPL_G1|1 IG1_0_RX _PG1_01|_SPL_G1|1  2.063e-12
L_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|1 _PG1_01|_SPL_G1|4  3.637e-12
L_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|7  1.278e-12
L_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|8  1.305e-12
L_PG1_01|_SPL_G1|5 _PG1_01|_SPL_G1|8 _PG1_01|G1_COPY_1  2.05e-12
L_PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|11  1.315e-12
L_PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|11 _PG1_01|G1_COPY_2  2.06e-12
L_PG1_01|_SPL_G1|P1 _PG1_01|_SPL_G1|2 0  4.676e-13
L_PG1_01|_SPL_G1|P2 _PG1_01|_SPL_G1|5 0  4.498e-13
L_PG1_01|_SPL_G1|P3 _PG1_01|_SPL_G1|9 0  5.183e-13
L_PG1_01|_SPL_G1|P4 _PG1_01|_SPL_G1|12 0  4.639e-13
R_PG1_01|_SPL_G1|B1 _PG1_01|_SPL_G1|1 _PG1_01|_SPL_G1|101  2.7439617672
L_PG1_01|_SPL_G1|RB1 _PG1_01|_SPL_G1|101 0  1.550338398468e-12
R_PG1_01|_SPL_G1|B2 _PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|104  2.286634806
L_PG1_01|_SPL_G1|RB2 _PG1_01|_SPL_G1|104 0  1.29194866539e-12
R_PG1_01|_SPL_G1|B3 _PG1_01|_SPL_G1|8 _PG1_01|_SPL_G1|108  2.7439617672
L_PG1_01|_SPL_G1|RB3 _PG1_01|_SPL_G1|108 0  1.550338398468e-12
R_PG1_01|_SPL_G1|B4 _PG1_01|_SPL_G1|11 _PG1_01|_SPL_G1|111  2.7439617672
L_PG1_01|_SPL_G1|RB4 _PG1_01|_SPL_G1|111 0  1.550338398468e-12
L_PG1_01|_PG|A1 IP1_0_TO1 _PG1_01|_PG|A1  2.067833848e-12
L_PG1_01|_PG|A2 _PG1_01|_PG|A1 _PG1_01|_PG|A2  4.135667696e-12
L_PG1_01|_PG|A3 _PG1_01|_PG|A3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|B1 _PG1_01|G1_COPY_1 _PG1_01|_PG|B1  2.067833848e-12
L_PG1_01|_PG|B2 _PG1_01|_PG|B1 _PG1_01|_PG|B2  4.135667696e-12
L_PG1_01|_PG|B3 _PG1_01|_PG|B3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|Q3 _PG1_01|_PG|Q3 _PG1_01|_PG|Q2  4.135667696e-12
L_PG1_01|_PG|Q2 _PG1_01|_PG|Q2 _PG1_01|_PG|Q1  4.135667696e-12
L_PG1_01|_PG|Q1 _PG1_01|_PG|Q1 _PG1_01|PG  2.067833848e-12
L_PG1_01|_GG|A1 IG0_0_TO1 _PG1_01|_GG|A1  2.067833848e-12
L_PG1_01|_GG|A2 _PG1_01|_GG|A1 _PG1_01|_GG|A2  4.135667696e-12
L_PG1_01|_GG|A3 _PG1_01|_GG|A3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|B1 _PG1_01|G1_COPY_2 _PG1_01|_GG|B1  2.067833848e-12
L_PG1_01|_GG|B2 _PG1_01|_GG|B1 _PG1_01|_GG|B2  4.135667696e-12
L_PG1_01|_GG|B3 _PG1_01|_GG|B3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|Q3 _PG1_01|_GG|Q3 _PG1_01|_GG|Q2  4.135667696e-12
L_PG1_01|_GG|Q2 _PG1_01|_GG|Q2 _PG1_01|_GG|Q1  4.135667696e-12
L_PG1_01|_GG|Q1 _PG1_01|_GG|Q1 _PG1_01|GG  2.067833848e-12
B_PG1_01|_DFF_PG|1 _PG1_01|_DFF_PG|1 _PG1_01|_DFF_PG|2 JJMIT AREA=2.5
B_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|5 JJMIT AREA=1.61
B_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|6 JJMIT AREA=1.54
B_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|8 _PG1_01|_DFF_PG|9 JJMIT AREA=1.69
B_PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|10 _PG1_01|_DFF_PG|8 JJMIT AREA=1.38
B_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|11 _PG1_01|_DFF_PG|12 JJMIT AREA=2.5
B_PG1_01|_DFF_PG|7 _PG1_01|_DFF_PG|14 _PG1_01|_DFF_PG|15 JJMIT AREA=2.5
I_PG1_01|_DFF_PG|B1 0 _PG1_01|_DFF_PG|3  PWL(0 0 5e-12 0.000175)
I_PG1_01|_DFF_PG|B2 0 _PG1_01|_DFF_PG|7  PWL(0 0 5e-12 0.000173)
I_PG1_01|_DFF_PG|B3 0 _PG1_01|_DFF_PG|13  PWL(0 0 5e-12 0.000175)
I_PG1_01|_DFF_PG|B4 0 _PG1_01|_DFF_PG|16  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|B1 _PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|1  2e-12
L_PG1_01|_DFF_PG|B2 _PG1_01|_DFF_PG|7 _PG1_01|_DFF_PG|5  2e-12
L_PG1_01|_DFF_PG|B3 _PG1_01|_DFF_PG|11 _PG1_01|_DFF_PG|13  2e-12
L_PG1_01|_DFF_PG|B4 _PG1_01|_DFF_PG|16 _PG1_01|_DFF_PG|14  2e-12
L_PG1_01|_DFF_PG|1 _PG1_01|PG _PG1_01|_DFF_PG|1  2.059e-12
L_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|1 _PG1_01|_DFF_PG|4  4.123e-12
L_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|8  6.873e-12
L_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|10 _PG1_01|_DFF_PG|11  5.195e-12
L_PG1_01|_DFF_PG|5 T05 _PG1_01|_DFF_PG|11  2.071e-12
L_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|8 _PG1_01|_DFF_PG|14  3.287e-12
L_PG1_01|_DFF_PG|7 _PG1_01|_DFF_PG|14 _PG1_01|PG_SYNC  2.066e-12
L_PG1_01|_DFF_PG|P1 _PG1_01|_DFF_PG|2 0  5.042e-13
L_PG1_01|_DFF_PG|P3 _PG1_01|_DFF_PG|6 0  5.799e-13
L_PG1_01|_DFF_PG|P4 _PG1_01|_DFF_PG|9 0  5.733e-13
L_PG1_01|_DFF_PG|P6 _PG1_01|_DFF_PG|12 0  4.605e-13
L_PG1_01|_DFF_PG|P7 _PG1_01|_DFF_PG|15 0  4.961e-13
R_PG1_01|_DFF_PG|B1 _PG1_01|_DFF_PG|1 _PG1_01|_DFF_PG|101  2.7439617672
L_PG1_01|_DFF_PG|RB1 _PG1_01|_DFF_PG|101 0  1.550338398468e-12
R_PG1_01|_DFF_PG|B2 _PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|104  4.260810197515528
L_PG1_01|_DFF_PG|RB2 _PG1_01|_DFF_PG|104 _PG1_01|_DFF_PG|5  2.407357761596273e-12
R_PG1_01|_DFF_PG|B3 _PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|105  4.454483388311688
L_PG1_01|_DFF_PG|RB3 _PG1_01|_DFF_PG|105 0  2.516783114396104e-12
R_PG1_01|_DFF_PG|B4 _PG1_01|_DFF_PG|8 _PG1_01|_DFF_PG|108  4.059115040236686
L_PG1_01|_DFF_PG|RB4 _PG1_01|_DFF_PG|108 0  2.2933999977337278e-12
R_PG1_01|_DFF_PG|B5 _PG1_01|_DFF_PG|10 _PG1_01|_DFF_PG|110  4.970945230434783
L_PG1_01|_DFF_PG|RB5 _PG1_01|_DFF_PG|110 _PG1_01|_DFF_PG|8  2.8085840551956523e-12
R_PG1_01|_DFF_PG|B6 _PG1_01|_DFF_PG|11 _PG1_01|_DFF_PG|111  2.7439617672
L_PG1_01|_DFF_PG|RB6 _PG1_01|_DFF_PG|111 0  1.550338398468e-12
R_PG1_01|_DFF_PG|B7 _PG1_01|_DFF_PG|14 _PG1_01|_DFF_PG|114  2.7439617672
L_PG1_01|_DFF_PG|RB7 _PG1_01|_DFF_PG|114 0  1.550338398468e-12
B_PG1_01|_DFF_GG|1 _PG1_01|_DFF_GG|1 _PG1_01|_DFF_GG|2 JJMIT AREA=2.5
B_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|5 JJMIT AREA=1.61
B_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|6 JJMIT AREA=1.54
B_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|8 _PG1_01|_DFF_GG|9 JJMIT AREA=1.69
B_PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|10 _PG1_01|_DFF_GG|8 JJMIT AREA=1.38
B_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|11 _PG1_01|_DFF_GG|12 JJMIT AREA=2.5
B_PG1_01|_DFF_GG|7 _PG1_01|_DFF_GG|14 _PG1_01|_DFF_GG|15 JJMIT AREA=2.5
I_PG1_01|_DFF_GG|B1 0 _PG1_01|_DFF_GG|3  PWL(0 0 5e-12 0.000175)
I_PG1_01|_DFF_GG|B2 0 _PG1_01|_DFF_GG|7  PWL(0 0 5e-12 0.000173)
I_PG1_01|_DFF_GG|B3 0 _PG1_01|_DFF_GG|13  PWL(0 0 5e-12 0.000175)
I_PG1_01|_DFF_GG|B4 0 _PG1_01|_DFF_GG|16  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|B1 _PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|1  2e-12
L_PG1_01|_DFF_GG|B2 _PG1_01|_DFF_GG|7 _PG1_01|_DFF_GG|5  2e-12
L_PG1_01|_DFF_GG|B3 _PG1_01|_DFF_GG|11 _PG1_01|_DFF_GG|13  2e-12
L_PG1_01|_DFF_GG|B4 _PG1_01|_DFF_GG|16 _PG1_01|_DFF_GG|14  2e-12
L_PG1_01|_DFF_GG|1 _PG1_01|GG _PG1_01|_DFF_GG|1  2.059e-12
L_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|1 _PG1_01|_DFF_GG|4  4.123e-12
L_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|8  6.873e-12
L_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|10 _PG1_01|_DFF_GG|11  5.195e-12
L_PG1_01|_DFF_GG|5 T05 _PG1_01|_DFF_GG|11  2.071e-12
L_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|8 _PG1_01|_DFF_GG|14  3.287e-12
L_PG1_01|_DFF_GG|7 _PG1_01|_DFF_GG|14 _PG1_01|GG_SYNC  2.066e-12
L_PG1_01|_DFF_GG|P1 _PG1_01|_DFF_GG|2 0  5.042e-13
L_PG1_01|_DFF_GG|P3 _PG1_01|_DFF_GG|6 0  5.799e-13
L_PG1_01|_DFF_GG|P4 _PG1_01|_DFF_GG|9 0  5.733e-13
L_PG1_01|_DFF_GG|P6 _PG1_01|_DFF_GG|12 0  4.605e-13
L_PG1_01|_DFF_GG|P7 _PG1_01|_DFF_GG|15 0  4.961e-13
R_PG1_01|_DFF_GG|B1 _PG1_01|_DFF_GG|1 _PG1_01|_DFF_GG|101  2.7439617672
L_PG1_01|_DFF_GG|RB1 _PG1_01|_DFF_GG|101 0  1.550338398468e-12
R_PG1_01|_DFF_GG|B2 _PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|104  4.260810197515528
L_PG1_01|_DFF_GG|RB2 _PG1_01|_DFF_GG|104 _PG1_01|_DFF_GG|5  2.407357761596273e-12
R_PG1_01|_DFF_GG|B3 _PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|105  4.454483388311688
L_PG1_01|_DFF_GG|RB3 _PG1_01|_DFF_GG|105 0  2.516783114396104e-12
R_PG1_01|_DFF_GG|B4 _PG1_01|_DFF_GG|8 _PG1_01|_DFF_GG|108  4.059115040236686
L_PG1_01|_DFF_GG|RB4 _PG1_01|_DFF_GG|108 0  2.2933999977337278e-12
R_PG1_01|_DFF_GG|B5 _PG1_01|_DFF_GG|10 _PG1_01|_DFF_GG|110  4.970945230434783
L_PG1_01|_DFF_GG|RB5 _PG1_01|_DFF_GG|110 _PG1_01|_DFF_GG|8  2.8085840551956523e-12
R_PG1_01|_DFF_GG|B6 _PG1_01|_DFF_GG|11 _PG1_01|_DFF_GG|111  2.7439617672
L_PG1_01|_DFF_GG|RB6 _PG1_01|_DFF_GG|111 0  1.550338398468e-12
R_PG1_01|_DFF_GG|B7 _PG1_01|_DFF_GG|14 _PG1_01|_DFF_GG|114  2.7439617672
L_PG1_01|_DFF_GG|RB7 _PG1_01|_DFF_GG|114 0  1.550338398468e-12
L_PG1_01|_AND_G|A1 _PG1_01|PG_SYNC _PG1_01|_AND_G|A1  2.067833848e-12
L_PG1_01|_AND_G|A2 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A2  4.135667696e-12
L_PG1_01|_AND_G|A3 _PG1_01|_AND_G|A3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|B1 _PG1_01|GG_SYNC _PG1_01|_AND_G|B1  2.067833848e-12
L_PG1_01|_AND_G|B2 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B2  4.135667696e-12
L_PG1_01|_AND_G|B3 _PG1_01|_AND_G|B3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q2  4.135667696e-12
L_PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q1  4.135667696e-12
L_PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1 G1_1  2.067833848e-12
B_PG2_01|P|1 _PG2_01|P|1 _PG2_01|P|2 JJMIT AREA=2.5
B_PG2_01|P|2 _PG2_01|P|4 _PG2_01|P|5 JJMIT AREA=1.61
B_PG2_01|P|3 _PG2_01|P|5 _PG2_01|P|6 JJMIT AREA=1.54
B_PG2_01|P|4 _PG2_01|P|8 _PG2_01|P|9 JJMIT AREA=1.69
B_PG2_01|P|5 _PG2_01|P|10 _PG2_01|P|8 JJMIT AREA=1.38
B_PG2_01|P|6 _PG2_01|P|11 _PG2_01|P|12 JJMIT AREA=2.5
B_PG2_01|P|7 _PG2_01|P|14 _PG2_01|P|15 JJMIT AREA=2.5
I_PG2_01|P|B1 0 _PG2_01|P|3  PWL(0 0 5e-12 0.000175)
I_PG2_01|P|B2 0 _PG2_01|P|7  PWL(0 0 5e-12 0.000173)
I_PG2_01|P|B3 0 _PG2_01|P|13  PWL(0 0 5e-12 0.000175)
I_PG2_01|P|B4 0 _PG2_01|P|16  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|B1 _PG2_01|P|3 _PG2_01|P|1  2e-12
L_PG2_01|P|B2 _PG2_01|P|7 _PG2_01|P|5  2e-12
L_PG2_01|P|B3 _PG2_01|P|11 _PG2_01|P|13  2e-12
L_PG2_01|P|B4 _PG2_01|P|16 _PG2_01|P|14  2e-12
L_PG2_01|P|1 IP2_0_TO2 _PG2_01|P|1  2.059e-12
L_PG2_01|P|2 _PG2_01|P|1 _PG2_01|P|4  4.123e-12
L_PG2_01|P|3 _PG2_01|P|5 _PG2_01|P|8  6.873e-12
L_PG2_01|P|4 _PG2_01|P|10 _PG2_01|P|11  5.195e-12
L_PG2_01|P|5 T06 _PG2_01|P|11  2.071e-12
L_PG2_01|P|6 _PG2_01|P|8 _PG2_01|P|14  3.287e-12
L_PG2_01|P|7 _PG2_01|P|14 P2_1  2.066e-12
L_PG2_01|P|P1 _PG2_01|P|2 0  5.042e-13
L_PG2_01|P|P3 _PG2_01|P|6 0  5.799e-13
L_PG2_01|P|P4 _PG2_01|P|9 0  5.733e-13
L_PG2_01|P|P6 _PG2_01|P|12 0  4.605e-13
L_PG2_01|P|P7 _PG2_01|P|15 0  4.961e-13
R_PG2_01|P|B1 _PG2_01|P|1 _PG2_01|P|101  2.7439617672
L_PG2_01|P|RB1 _PG2_01|P|101 0  1.550338398468e-12
R_PG2_01|P|B2 _PG2_01|P|4 _PG2_01|P|104  4.260810197515528
L_PG2_01|P|RB2 _PG2_01|P|104 _PG2_01|P|5  2.407357761596273e-12
R_PG2_01|P|B3 _PG2_01|P|5 _PG2_01|P|105  4.454483388311688
L_PG2_01|P|RB3 _PG2_01|P|105 0  2.516783114396104e-12
R_PG2_01|P|B4 _PG2_01|P|8 _PG2_01|P|108  4.059115040236686
L_PG2_01|P|RB4 _PG2_01|P|108 0  2.2933999977337278e-12
R_PG2_01|P|B5 _PG2_01|P|10 _PG2_01|P|110  4.970945230434783
L_PG2_01|P|RB5 _PG2_01|P|110 _PG2_01|P|8  2.8085840551956523e-12
R_PG2_01|P|B6 _PG2_01|P|11 _PG2_01|P|111  2.7439617672
L_PG2_01|P|RB6 _PG2_01|P|111 0  1.550338398468e-12
R_PG2_01|P|B7 _PG2_01|P|14 _PG2_01|P|114  2.7439617672
L_PG2_01|P|RB7 _PG2_01|P|114 0  1.550338398468e-12
B_PG2_01|G|1 _PG2_01|G|1 _PG2_01|G|2 JJMIT AREA=2.5
B_PG2_01|G|2 _PG2_01|G|4 _PG2_01|G|5 JJMIT AREA=1.61
B_PG2_01|G|3 _PG2_01|G|5 _PG2_01|G|6 JJMIT AREA=1.54
B_PG2_01|G|4 _PG2_01|G|8 _PG2_01|G|9 JJMIT AREA=1.69
B_PG2_01|G|5 _PG2_01|G|10 _PG2_01|G|8 JJMIT AREA=1.38
B_PG2_01|G|6 _PG2_01|G|11 _PG2_01|G|12 JJMIT AREA=2.5
B_PG2_01|G|7 _PG2_01|G|14 _PG2_01|G|15 JJMIT AREA=2.5
I_PG2_01|G|B1 0 _PG2_01|G|3  PWL(0 0 5e-12 0.000175)
I_PG2_01|G|B2 0 _PG2_01|G|7  PWL(0 0 5e-12 0.000173)
I_PG2_01|G|B3 0 _PG2_01|G|13  PWL(0 0 5e-12 0.000175)
I_PG2_01|G|B4 0 _PG2_01|G|16  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|B1 _PG2_01|G|3 _PG2_01|G|1  2e-12
L_PG2_01|G|B2 _PG2_01|G|7 _PG2_01|G|5  2e-12
L_PG2_01|G|B3 _PG2_01|G|11 _PG2_01|G|13  2e-12
L_PG2_01|G|B4 _PG2_01|G|16 _PG2_01|G|14  2e-12
L_PG2_01|G|1 IG2_0_TO2 _PG2_01|G|1  2.059e-12
L_PG2_01|G|2 _PG2_01|G|1 _PG2_01|G|4  4.123e-12
L_PG2_01|G|3 _PG2_01|G|5 _PG2_01|G|8  6.873e-12
L_PG2_01|G|4 _PG2_01|G|10 _PG2_01|G|11  5.195e-12
L_PG2_01|G|5 T06 _PG2_01|G|11  2.071e-12
L_PG2_01|G|6 _PG2_01|G|8 _PG2_01|G|14  3.287e-12
L_PG2_01|G|7 _PG2_01|G|14 G2_1  2.066e-12
L_PG2_01|G|P1 _PG2_01|G|2 0  5.042e-13
L_PG2_01|G|P3 _PG2_01|G|6 0  5.799e-13
L_PG2_01|G|P4 _PG2_01|G|9 0  5.733e-13
L_PG2_01|G|P6 _PG2_01|G|12 0  4.605e-13
L_PG2_01|G|P7 _PG2_01|G|15 0  4.961e-13
R_PG2_01|G|B1 _PG2_01|G|1 _PG2_01|G|101  2.7439617672
L_PG2_01|G|RB1 _PG2_01|G|101 0  1.550338398468e-12
R_PG2_01|G|B2 _PG2_01|G|4 _PG2_01|G|104  4.260810197515528
L_PG2_01|G|RB2 _PG2_01|G|104 _PG2_01|G|5  2.407357761596273e-12
R_PG2_01|G|B3 _PG2_01|G|5 _PG2_01|G|105  4.454483388311688
L_PG2_01|G|RB3 _PG2_01|G|105 0  2.516783114396104e-12
R_PG2_01|G|B4 _PG2_01|G|8 _PG2_01|G|108  4.059115040236686
L_PG2_01|G|RB4 _PG2_01|G|108 0  2.2933999977337278e-12
R_PG2_01|G|B5 _PG2_01|G|10 _PG2_01|G|110  4.970945230434783
L_PG2_01|G|RB5 _PG2_01|G|110 _PG2_01|G|8  2.8085840551956523e-12
R_PG2_01|G|B6 _PG2_01|G|11 _PG2_01|G|111  2.7439617672
L_PG2_01|G|RB6 _PG2_01|G|111 0  1.550338398468e-12
R_PG2_01|G|B7 _PG2_01|G|14 _PG2_01|G|114  2.7439617672
L_PG2_01|G|RB7 _PG2_01|G|114 0  1.550338398468e-12
I_PG3_01|_SPL_G1|B1 0 _PG3_01|_SPL_G1|3  PWL(0 0 5e-12 0.000175)
I_PG3_01|_SPL_G1|B2 0 _PG3_01|_SPL_G1|6  PWL(0 0 5e-12 0.00028)
I_PG3_01|_SPL_G1|B3 0 _PG3_01|_SPL_G1|10  PWL(0 0 5e-12 0.000175)
I_PG3_01|_SPL_G1|B4 0 _PG3_01|_SPL_G1|13  PWL(0 0 5e-12 0.000175)
L_PG3_01|_SPL_G1|B1 _PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|1  9.175e-13
L_PG3_01|_SPL_G1|B2 _PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|4  7.666e-13
L_PG3_01|_SPL_G1|B3 _PG3_01|_SPL_G1|10 _PG3_01|_SPL_G1|8  1.928e-12
L_PG3_01|_SPL_G1|B4 _PG3_01|_SPL_G1|13 _PG3_01|_SPL_G1|11  8.786e-13
B_PG3_01|_SPL_G1|1 _PG3_01|_SPL_G1|1 _PG3_01|_SPL_G1|2 JJMIT AREA=2.5
B_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|5 JJMIT AREA=3.0
B_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|8 _PG3_01|_SPL_G1|9 JJMIT AREA=2.5
B_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|11 _PG3_01|_SPL_G1|12 JJMIT AREA=2.5
L_PG3_01|_SPL_G1|1 IG3_0_RX _PG3_01|_SPL_G1|1  2.063e-12
L_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|1 _PG3_01|_SPL_G1|4  3.637e-12
L_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|7  1.278e-12
L_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|8  1.305e-12
L_PG3_01|_SPL_G1|5 _PG3_01|_SPL_G1|8 _PG3_01|G1_COPY_1  2.05e-12
L_PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|11  1.315e-12
L_PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|11 _PG3_01|G1_COPY_2  2.06e-12
L_PG3_01|_SPL_G1|P1 _PG3_01|_SPL_G1|2 0  4.676e-13
L_PG3_01|_SPL_G1|P2 _PG3_01|_SPL_G1|5 0  4.498e-13
L_PG3_01|_SPL_G1|P3 _PG3_01|_SPL_G1|9 0  5.183e-13
L_PG3_01|_SPL_G1|P4 _PG3_01|_SPL_G1|12 0  4.639e-13
R_PG3_01|_SPL_G1|B1 _PG3_01|_SPL_G1|1 _PG3_01|_SPL_G1|101  2.7439617672
L_PG3_01|_SPL_G1|RB1 _PG3_01|_SPL_G1|101 0  1.550338398468e-12
R_PG3_01|_SPL_G1|B2 _PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|104  2.286634806
L_PG3_01|_SPL_G1|RB2 _PG3_01|_SPL_G1|104 0  1.29194866539e-12
R_PG3_01|_SPL_G1|B3 _PG3_01|_SPL_G1|8 _PG3_01|_SPL_G1|108  2.7439617672
L_PG3_01|_SPL_G1|RB3 _PG3_01|_SPL_G1|108 0  1.550338398468e-12
R_PG3_01|_SPL_G1|B4 _PG3_01|_SPL_G1|11 _PG3_01|_SPL_G1|111  2.7439617672
L_PG3_01|_SPL_G1|RB4 _PG3_01|_SPL_G1|111 0  1.550338398468e-12
I_PG3_01|_SPL_P1|B1 0 _PG3_01|_SPL_P1|3  PWL(0 0 5e-12 0.000175)
I_PG3_01|_SPL_P1|B2 0 _PG3_01|_SPL_P1|6  PWL(0 0 5e-12 0.00028)
I_PG3_01|_SPL_P1|B3 0 _PG3_01|_SPL_P1|10  PWL(0 0 5e-12 0.000175)
I_PG3_01|_SPL_P1|B4 0 _PG3_01|_SPL_P1|13  PWL(0 0 5e-12 0.000175)
L_PG3_01|_SPL_P1|B1 _PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|1  9.175e-13
L_PG3_01|_SPL_P1|B2 _PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|4  7.666e-13
L_PG3_01|_SPL_P1|B3 _PG3_01|_SPL_P1|10 _PG3_01|_SPL_P1|8  1.928e-12
L_PG3_01|_SPL_P1|B4 _PG3_01|_SPL_P1|13 _PG3_01|_SPL_P1|11  8.786e-13
B_PG3_01|_SPL_P1|1 _PG3_01|_SPL_P1|1 _PG3_01|_SPL_P1|2 JJMIT AREA=2.5
B_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|5 JJMIT AREA=3.0
B_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|8 _PG3_01|_SPL_P1|9 JJMIT AREA=2.5
B_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|11 _PG3_01|_SPL_P1|12 JJMIT AREA=2.5
L_PG3_01|_SPL_P1|1 IP3_0_TO1 _PG3_01|_SPL_P1|1  2.063e-12
L_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|1 _PG3_01|_SPL_P1|4  3.637e-12
L_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|7  1.278e-12
L_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|8  1.305e-12
L_PG3_01|_SPL_P1|5 _PG3_01|_SPL_P1|8 _PG3_01|P1_COPY_1  2.05e-12
L_PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|11  1.315e-12
L_PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|11 _PG3_01|P1_COPY_2  2.06e-12
L_PG3_01|_SPL_P1|P1 _PG3_01|_SPL_P1|2 0  4.676e-13
L_PG3_01|_SPL_P1|P2 _PG3_01|_SPL_P1|5 0  4.498e-13
L_PG3_01|_SPL_P1|P3 _PG3_01|_SPL_P1|9 0  5.183e-13
L_PG3_01|_SPL_P1|P4 _PG3_01|_SPL_P1|12 0  4.639e-13
R_PG3_01|_SPL_P1|B1 _PG3_01|_SPL_P1|1 _PG3_01|_SPL_P1|101  2.7439617672
L_PG3_01|_SPL_P1|RB1 _PG3_01|_SPL_P1|101 0  1.550338398468e-12
R_PG3_01|_SPL_P1|B2 _PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|104  2.286634806
L_PG3_01|_SPL_P1|RB2 _PG3_01|_SPL_P1|104 0  1.29194866539e-12
R_PG3_01|_SPL_P1|B3 _PG3_01|_SPL_P1|8 _PG3_01|_SPL_P1|108  2.7439617672
L_PG3_01|_SPL_P1|RB3 _PG3_01|_SPL_P1|108 0  1.550338398468e-12
R_PG3_01|_SPL_P1|B4 _PG3_01|_SPL_P1|11 _PG3_01|_SPL_P1|111  2.7439617672
L_PG3_01|_SPL_P1|RB4 _PG3_01|_SPL_P1|111 0  1.550338398468e-12
L_PG3_01|_PG|A1 _PG3_01|P1_COPY_1 _PG3_01|_PG|A1  2.067833848e-12
L_PG3_01|_PG|A2 _PG3_01|_PG|A1 _PG3_01|_PG|A2  4.135667696e-12
L_PG3_01|_PG|A3 _PG3_01|_PG|A3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|B1 _PG3_01|G1_COPY_1 _PG3_01|_PG|B1  2.067833848e-12
L_PG3_01|_PG|B2 _PG3_01|_PG|B1 _PG3_01|_PG|B2  4.135667696e-12
L_PG3_01|_PG|B3 _PG3_01|_PG|B3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|Q3 _PG3_01|_PG|Q3 _PG3_01|_PG|Q2  4.135667696e-12
L_PG3_01|_PG|Q2 _PG3_01|_PG|Q2 _PG3_01|_PG|Q1  4.135667696e-12
L_PG3_01|_PG|Q1 _PG3_01|_PG|Q1 _PG3_01|PG  2.067833848e-12
L_PG3_01|_GG|A1 IG2_0_TO3 _PG3_01|_GG|A1  2.067833848e-12
L_PG3_01|_GG|A2 _PG3_01|_GG|A1 _PG3_01|_GG|A2  4.135667696e-12
L_PG3_01|_GG|A3 _PG3_01|_GG|A3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|B1 _PG3_01|G1_COPY_2 _PG3_01|_GG|B1  2.067833848e-12
L_PG3_01|_GG|B2 _PG3_01|_GG|B1 _PG3_01|_GG|B2  4.135667696e-12
L_PG3_01|_GG|B3 _PG3_01|_GG|B3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|Q3 _PG3_01|_GG|Q3 _PG3_01|_GG|Q2  4.135667696e-12
L_PG3_01|_GG|Q2 _PG3_01|_GG|Q2 _PG3_01|_GG|Q1  4.135667696e-12
L_PG3_01|_GG|Q1 _PG3_01|_GG|Q1 _PG3_01|GG  2.067833848e-12
B_PG3_01|_DFF_P0|1 _PG3_01|_DFF_P0|1 _PG3_01|_DFF_P0|2 JJMIT AREA=2.5
B_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|5 JJMIT AREA=1.61
B_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|6 JJMIT AREA=1.54
B_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|8 _PG3_01|_DFF_P0|9 JJMIT AREA=1.69
B_PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|10 _PG3_01|_DFF_P0|8 JJMIT AREA=1.38
B_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|11 _PG3_01|_DFF_P0|12 JJMIT AREA=2.5
B_PG3_01|_DFF_P0|7 _PG3_01|_DFF_P0|14 _PG3_01|_DFF_P0|15 JJMIT AREA=2.5
I_PG3_01|_DFF_P0|B1 0 _PG3_01|_DFF_P0|3  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_P0|B2 0 _PG3_01|_DFF_P0|7  PWL(0 0 5e-12 0.000173)
I_PG3_01|_DFF_P0|B3 0 _PG3_01|_DFF_P0|13  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_P0|B4 0 _PG3_01|_DFF_P0|16  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|B1 _PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|1  2e-12
L_PG3_01|_DFF_P0|B2 _PG3_01|_DFF_P0|7 _PG3_01|_DFF_P0|5  2e-12
L_PG3_01|_DFF_P0|B3 _PG3_01|_DFF_P0|11 _PG3_01|_DFF_P0|13  2e-12
L_PG3_01|_DFF_P0|B4 _PG3_01|_DFF_P0|16 _PG3_01|_DFF_P0|14  2e-12
L_PG3_01|_DFF_P0|1 IP2_0_TO3 _PG3_01|_DFF_P0|1  2.059e-12
L_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|1 _PG3_01|_DFF_P0|4  4.123e-12
L_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|8  6.873e-12
L_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|10 _PG3_01|_DFF_P0|11  5.195e-12
L_PG3_01|_DFF_P0|5 T07 _PG3_01|_DFF_P0|11  2.071e-12
L_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|8 _PG3_01|_DFF_P0|14  3.287e-12
L_PG3_01|_DFF_P0|7 _PG3_01|_DFF_P0|14 _PG3_01|P0_SYNC  2.066e-12
L_PG3_01|_DFF_P0|P1 _PG3_01|_DFF_P0|2 0  5.042e-13
L_PG3_01|_DFF_P0|P3 _PG3_01|_DFF_P0|6 0  5.799e-13
L_PG3_01|_DFF_P0|P4 _PG3_01|_DFF_P0|9 0  5.733e-13
L_PG3_01|_DFF_P0|P6 _PG3_01|_DFF_P0|12 0  4.605e-13
L_PG3_01|_DFF_P0|P7 _PG3_01|_DFF_P0|15 0  4.961e-13
R_PG3_01|_DFF_P0|B1 _PG3_01|_DFF_P0|1 _PG3_01|_DFF_P0|101  2.7439617672
L_PG3_01|_DFF_P0|RB1 _PG3_01|_DFF_P0|101 0  1.550338398468e-12
R_PG3_01|_DFF_P0|B2 _PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|104  4.260810197515528
L_PG3_01|_DFF_P0|RB2 _PG3_01|_DFF_P0|104 _PG3_01|_DFF_P0|5  2.407357761596273e-12
R_PG3_01|_DFF_P0|B3 _PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|105  4.454483388311688
L_PG3_01|_DFF_P0|RB3 _PG3_01|_DFF_P0|105 0  2.516783114396104e-12
R_PG3_01|_DFF_P0|B4 _PG3_01|_DFF_P0|8 _PG3_01|_DFF_P0|108  4.059115040236686
L_PG3_01|_DFF_P0|RB4 _PG3_01|_DFF_P0|108 0  2.2933999977337278e-12
R_PG3_01|_DFF_P0|B5 _PG3_01|_DFF_P0|10 _PG3_01|_DFF_P0|110  4.970945230434783
L_PG3_01|_DFF_P0|RB5 _PG3_01|_DFF_P0|110 _PG3_01|_DFF_P0|8  2.8085840551956523e-12
R_PG3_01|_DFF_P0|B6 _PG3_01|_DFF_P0|11 _PG3_01|_DFF_P0|111  2.7439617672
L_PG3_01|_DFF_P0|RB6 _PG3_01|_DFF_P0|111 0  1.550338398468e-12
R_PG3_01|_DFF_P0|B7 _PG3_01|_DFF_P0|14 _PG3_01|_DFF_P0|114  2.7439617672
L_PG3_01|_DFF_P0|RB7 _PG3_01|_DFF_P0|114 0  1.550338398468e-12
B_PG3_01|_DFF_P1|1 _PG3_01|_DFF_P1|1 _PG3_01|_DFF_P1|2 JJMIT AREA=2.5
B_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|5 JJMIT AREA=1.61
B_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|6 JJMIT AREA=1.54
B_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|8 _PG3_01|_DFF_P1|9 JJMIT AREA=1.69
B_PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|10 _PG3_01|_DFF_P1|8 JJMIT AREA=1.38
B_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|11 _PG3_01|_DFF_P1|12 JJMIT AREA=2.5
B_PG3_01|_DFF_P1|7 _PG3_01|_DFF_P1|14 _PG3_01|_DFF_P1|15 JJMIT AREA=2.5
I_PG3_01|_DFF_P1|B1 0 _PG3_01|_DFF_P1|3  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_P1|B2 0 _PG3_01|_DFF_P1|7  PWL(0 0 5e-12 0.000173)
I_PG3_01|_DFF_P1|B3 0 _PG3_01|_DFF_P1|13  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_P1|B4 0 _PG3_01|_DFF_P1|16  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|B1 _PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|1  2e-12
L_PG3_01|_DFF_P1|B2 _PG3_01|_DFF_P1|7 _PG3_01|_DFF_P1|5  2e-12
L_PG3_01|_DFF_P1|B3 _PG3_01|_DFF_P1|11 _PG3_01|_DFF_P1|13  2e-12
L_PG3_01|_DFF_P1|B4 _PG3_01|_DFF_P1|16 _PG3_01|_DFF_P1|14  2e-12
L_PG3_01|_DFF_P1|1 _PG3_01|P1_COPY_2 _PG3_01|_DFF_P1|1  2.059e-12
L_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|1 _PG3_01|_DFF_P1|4  4.123e-12
L_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|8  6.873e-12
L_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|10 _PG3_01|_DFF_P1|11  5.195e-12
L_PG3_01|_DFF_P1|5 T07 _PG3_01|_DFF_P1|11  2.071e-12
L_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|8 _PG3_01|_DFF_P1|14  3.287e-12
L_PG3_01|_DFF_P1|7 _PG3_01|_DFF_P1|14 _PG3_01|P1_SYNC  2.066e-12
L_PG3_01|_DFF_P1|P1 _PG3_01|_DFF_P1|2 0  5.042e-13
L_PG3_01|_DFF_P1|P3 _PG3_01|_DFF_P1|6 0  5.799e-13
L_PG3_01|_DFF_P1|P4 _PG3_01|_DFF_P1|9 0  5.733e-13
L_PG3_01|_DFF_P1|P6 _PG3_01|_DFF_P1|12 0  4.605e-13
L_PG3_01|_DFF_P1|P7 _PG3_01|_DFF_P1|15 0  4.961e-13
R_PG3_01|_DFF_P1|B1 _PG3_01|_DFF_P1|1 _PG3_01|_DFF_P1|101  2.7439617672
L_PG3_01|_DFF_P1|RB1 _PG3_01|_DFF_P1|101 0  1.550338398468e-12
R_PG3_01|_DFF_P1|B2 _PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|104  4.260810197515528
L_PG3_01|_DFF_P1|RB2 _PG3_01|_DFF_P1|104 _PG3_01|_DFF_P1|5  2.407357761596273e-12
R_PG3_01|_DFF_P1|B3 _PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|105  4.454483388311688
L_PG3_01|_DFF_P1|RB3 _PG3_01|_DFF_P1|105 0  2.516783114396104e-12
R_PG3_01|_DFF_P1|B4 _PG3_01|_DFF_P1|8 _PG3_01|_DFF_P1|108  4.059115040236686
L_PG3_01|_DFF_P1|RB4 _PG3_01|_DFF_P1|108 0  2.2933999977337278e-12
R_PG3_01|_DFF_P1|B5 _PG3_01|_DFF_P1|10 _PG3_01|_DFF_P1|110  4.970945230434783
L_PG3_01|_DFF_P1|RB5 _PG3_01|_DFF_P1|110 _PG3_01|_DFF_P1|8  2.8085840551956523e-12
R_PG3_01|_DFF_P1|B6 _PG3_01|_DFF_P1|11 _PG3_01|_DFF_P1|111  2.7439617672
L_PG3_01|_DFF_P1|RB6 _PG3_01|_DFF_P1|111 0  1.550338398468e-12
R_PG3_01|_DFF_P1|B7 _PG3_01|_DFF_P1|14 _PG3_01|_DFF_P1|114  2.7439617672
L_PG3_01|_DFF_P1|RB7 _PG3_01|_DFF_P1|114 0  1.550338398468e-12
B_PG3_01|_DFF_PG|1 _PG3_01|_DFF_PG|1 _PG3_01|_DFF_PG|2 JJMIT AREA=2.5
B_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|5 JJMIT AREA=1.61
B_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|6 JJMIT AREA=1.54
B_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|8 _PG3_01|_DFF_PG|9 JJMIT AREA=1.69
B_PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|10 _PG3_01|_DFF_PG|8 JJMIT AREA=1.38
B_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|11 _PG3_01|_DFF_PG|12 JJMIT AREA=2.5
B_PG3_01|_DFF_PG|7 _PG3_01|_DFF_PG|14 _PG3_01|_DFF_PG|15 JJMIT AREA=2.5
I_PG3_01|_DFF_PG|B1 0 _PG3_01|_DFF_PG|3  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_PG|B2 0 _PG3_01|_DFF_PG|7  PWL(0 0 5e-12 0.000173)
I_PG3_01|_DFF_PG|B3 0 _PG3_01|_DFF_PG|13  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_PG|B4 0 _PG3_01|_DFF_PG|16  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|B1 _PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|1  2e-12
L_PG3_01|_DFF_PG|B2 _PG3_01|_DFF_PG|7 _PG3_01|_DFF_PG|5  2e-12
L_PG3_01|_DFF_PG|B3 _PG3_01|_DFF_PG|11 _PG3_01|_DFF_PG|13  2e-12
L_PG3_01|_DFF_PG|B4 _PG3_01|_DFF_PG|16 _PG3_01|_DFF_PG|14  2e-12
L_PG3_01|_DFF_PG|1 _PG3_01|PG _PG3_01|_DFF_PG|1  2.059e-12
L_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|1 _PG3_01|_DFF_PG|4  4.123e-12
L_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|8  6.873e-12
L_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|10 _PG3_01|_DFF_PG|11  5.195e-12
L_PG3_01|_DFF_PG|5 T07 _PG3_01|_DFF_PG|11  2.071e-12
L_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|8 _PG3_01|_DFF_PG|14  3.287e-12
L_PG3_01|_DFF_PG|7 _PG3_01|_DFF_PG|14 _PG3_01|PG_SYNC  2.066e-12
L_PG3_01|_DFF_PG|P1 _PG3_01|_DFF_PG|2 0  5.042e-13
L_PG3_01|_DFF_PG|P3 _PG3_01|_DFF_PG|6 0  5.799e-13
L_PG3_01|_DFF_PG|P4 _PG3_01|_DFF_PG|9 0  5.733e-13
L_PG3_01|_DFF_PG|P6 _PG3_01|_DFF_PG|12 0  4.605e-13
L_PG3_01|_DFF_PG|P7 _PG3_01|_DFF_PG|15 0  4.961e-13
R_PG3_01|_DFF_PG|B1 _PG3_01|_DFF_PG|1 _PG3_01|_DFF_PG|101  2.7439617672
L_PG3_01|_DFF_PG|RB1 _PG3_01|_DFF_PG|101 0  1.550338398468e-12
R_PG3_01|_DFF_PG|B2 _PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|104  4.260810197515528
L_PG3_01|_DFF_PG|RB2 _PG3_01|_DFF_PG|104 _PG3_01|_DFF_PG|5  2.407357761596273e-12
R_PG3_01|_DFF_PG|B3 _PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|105  4.454483388311688
L_PG3_01|_DFF_PG|RB3 _PG3_01|_DFF_PG|105 0  2.516783114396104e-12
R_PG3_01|_DFF_PG|B4 _PG3_01|_DFF_PG|8 _PG3_01|_DFF_PG|108  4.059115040236686
L_PG3_01|_DFF_PG|RB4 _PG3_01|_DFF_PG|108 0  2.2933999977337278e-12
R_PG3_01|_DFF_PG|B5 _PG3_01|_DFF_PG|10 _PG3_01|_DFF_PG|110  4.970945230434783
L_PG3_01|_DFF_PG|RB5 _PG3_01|_DFF_PG|110 _PG3_01|_DFF_PG|8  2.8085840551956523e-12
R_PG3_01|_DFF_PG|B6 _PG3_01|_DFF_PG|11 _PG3_01|_DFF_PG|111  2.7439617672
L_PG3_01|_DFF_PG|RB6 _PG3_01|_DFF_PG|111 0  1.550338398468e-12
R_PG3_01|_DFF_PG|B7 _PG3_01|_DFF_PG|14 _PG3_01|_DFF_PG|114  2.7439617672
L_PG3_01|_DFF_PG|RB7 _PG3_01|_DFF_PG|114 0  1.550338398468e-12
B_PG3_01|_DFF_GG|1 _PG3_01|_DFF_GG|1 _PG3_01|_DFF_GG|2 JJMIT AREA=2.5
B_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|5 JJMIT AREA=1.61
B_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|6 JJMIT AREA=1.54
B_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|8 _PG3_01|_DFF_GG|9 JJMIT AREA=1.69
B_PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|10 _PG3_01|_DFF_GG|8 JJMIT AREA=1.38
B_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|11 _PG3_01|_DFF_GG|12 JJMIT AREA=2.5
B_PG3_01|_DFF_GG|7 _PG3_01|_DFF_GG|14 _PG3_01|_DFF_GG|15 JJMIT AREA=2.5
I_PG3_01|_DFF_GG|B1 0 _PG3_01|_DFF_GG|3  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_GG|B2 0 _PG3_01|_DFF_GG|7  PWL(0 0 5e-12 0.000173)
I_PG3_01|_DFF_GG|B3 0 _PG3_01|_DFF_GG|13  PWL(0 0 5e-12 0.000175)
I_PG3_01|_DFF_GG|B4 0 _PG3_01|_DFF_GG|16  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|B1 _PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|1  2e-12
L_PG3_01|_DFF_GG|B2 _PG3_01|_DFF_GG|7 _PG3_01|_DFF_GG|5  2e-12
L_PG3_01|_DFF_GG|B3 _PG3_01|_DFF_GG|11 _PG3_01|_DFF_GG|13  2e-12
L_PG3_01|_DFF_GG|B4 _PG3_01|_DFF_GG|16 _PG3_01|_DFF_GG|14  2e-12
L_PG3_01|_DFF_GG|1 _PG3_01|GG _PG3_01|_DFF_GG|1  2.059e-12
L_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|1 _PG3_01|_DFF_GG|4  4.123e-12
L_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|8  6.873e-12
L_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|10 _PG3_01|_DFF_GG|11  5.195e-12
L_PG3_01|_DFF_GG|5 T07 _PG3_01|_DFF_GG|11  2.071e-12
L_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|8 _PG3_01|_DFF_GG|14  3.287e-12
L_PG3_01|_DFF_GG|7 _PG3_01|_DFF_GG|14 _PG3_01|GG_SYNC  2.066e-12
L_PG3_01|_DFF_GG|P1 _PG3_01|_DFF_GG|2 0  5.042e-13
L_PG3_01|_DFF_GG|P3 _PG3_01|_DFF_GG|6 0  5.799e-13
L_PG3_01|_DFF_GG|P4 _PG3_01|_DFF_GG|9 0  5.733e-13
L_PG3_01|_DFF_GG|P6 _PG3_01|_DFF_GG|12 0  4.605e-13
L_PG3_01|_DFF_GG|P7 _PG3_01|_DFF_GG|15 0  4.961e-13
R_PG3_01|_DFF_GG|B1 _PG3_01|_DFF_GG|1 _PG3_01|_DFF_GG|101  2.7439617672
L_PG3_01|_DFF_GG|RB1 _PG3_01|_DFF_GG|101 0  1.550338398468e-12
R_PG3_01|_DFF_GG|B2 _PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|104  4.260810197515528
L_PG3_01|_DFF_GG|RB2 _PG3_01|_DFF_GG|104 _PG3_01|_DFF_GG|5  2.407357761596273e-12
R_PG3_01|_DFF_GG|B3 _PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|105  4.454483388311688
L_PG3_01|_DFF_GG|RB3 _PG3_01|_DFF_GG|105 0  2.516783114396104e-12
R_PG3_01|_DFF_GG|B4 _PG3_01|_DFF_GG|8 _PG3_01|_DFF_GG|108  4.059115040236686
L_PG3_01|_DFF_GG|RB4 _PG3_01|_DFF_GG|108 0  2.2933999977337278e-12
R_PG3_01|_DFF_GG|B5 _PG3_01|_DFF_GG|10 _PG3_01|_DFF_GG|110  4.970945230434783
L_PG3_01|_DFF_GG|RB5 _PG3_01|_DFF_GG|110 _PG3_01|_DFF_GG|8  2.8085840551956523e-12
R_PG3_01|_DFF_GG|B6 _PG3_01|_DFF_GG|11 _PG3_01|_DFF_GG|111  2.7439617672
L_PG3_01|_DFF_GG|RB6 _PG3_01|_DFF_GG|111 0  1.550338398468e-12
R_PG3_01|_DFF_GG|B7 _PG3_01|_DFF_GG|14 _PG3_01|_DFF_GG|114  2.7439617672
L_PG3_01|_DFF_GG|RB7 _PG3_01|_DFF_GG|114 0  1.550338398468e-12
L_PG3_01|_AND_G|A1 _PG3_01|PG_SYNC _PG3_01|_AND_G|A1  2.067833848e-12
L_PG3_01|_AND_G|A2 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A2  4.135667696e-12
L_PG3_01|_AND_G|A3 _PG3_01|_AND_G|A3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|B1 _PG3_01|GG_SYNC _PG3_01|_AND_G|B1  2.067833848e-12
L_PG3_01|_AND_G|B2 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B2  4.135667696e-12
L_PG3_01|_AND_G|B3 _PG3_01|_AND_G|B3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q2  4.135667696e-12
L_PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q1  4.135667696e-12
L_PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1 G3_1  2.067833848e-12
L_PG3_01|_AND_P|A1 _PG3_01|P0_SYNC _PG3_01|_AND_P|A1  2.067833848e-12
L_PG3_01|_AND_P|A2 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A2  4.135667696e-12
L_PG3_01|_AND_P|A3 _PG3_01|_AND_P|A3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|B1 _PG3_01|P1_SYNC _PG3_01|_AND_P|B1  2.067833848e-12
L_PG3_01|_AND_P|B2 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B2  4.135667696e-12
L_PG3_01|_AND_P|B3 _PG3_01|_AND_P|B3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q2  4.135667696e-12
L_PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q1  4.135667696e-12
L_PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1 P3_1  2.067833848e-12
B_PTL_P0_1|_TX|1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|2 JJMIT AREA=2.5
B_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|5 JJMIT AREA=2.5
I_PTL_P0_1|_TX|B1 0 _PTL_P0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_1|_TX|B2 0 _PTL_P0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|3  1.684e-12
L_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|6  3.596e-12
L_PTL_P0_1|_TX|1 P0_1 _PTL_P0_1|_TX|1  2.063e-12
L_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|4  4.123e-12
L_PTL_P0_1|_TX|3 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|7  2.193e-12
R_PTL_P0_1|_TX|D _PTL_P0_1|_TX|7 _PTL_P0_1|A_PTL  1.36
L_PTL_P0_1|_TX|P1 _PTL_P0_1|_TX|2 0  5.254e-13
L_PTL_P0_1|_TX|P2 _PTL_P0_1|_TX|5 0  5.141e-13
R_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|101  2.7439617672
R_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|104  2.7439617672
L_PTL_P0_1|_TX|RB1 _PTL_P0_1|_TX|101 0  1.550338398468e-12
L_PTL_P0_1|_TX|RB2 _PTL_P0_1|_TX|104 0  1.550338398468e-12
B_PTL_P0_1|_RX|1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|5 JJMIT AREA=2.0
B_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|8 JJMIT AREA=2.5
I_PTL_P0_1|_RX|B1 0 _PTL_P0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|3  2.777e-12
I_PTL_P0_1|_RX|B2 0 _PTL_P0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|6  2.685e-12
I_PTL_P0_1|_RX|B3 0 _PTL_P0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|9  2.764e-12
L_PTL_P0_1|_RX|1 _PTL_P0_1|A_PTL _PTL_P0_1|_RX|1  1.346e-12
L_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|4  6.348e-12
L_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7  5.197e-12
L_PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7 P0_1_RX  2.058e-12
L_PTL_P0_1|_RX|P1 _PTL_P0_1|_RX|2 0  4.795e-13
L_PTL_P0_1|_RX|P2 _PTL_P0_1|_RX|5 0  5.431e-13
L_PTL_P0_1|_RX|P3 _PTL_P0_1|_RX|8 0  5.339e-13
R_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|101  4.225701121488
R_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|104  3.429952209
R_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|107  2.7439617672
L_PTL_P0_1|_RX|RB1 _PTL_P0_1|_RX|101 0  2.38752113364072e-12
L_PTL_P0_1|_RX|RB2 _PTL_P0_1|_RX|104 0  1.937922998085e-12
L_PTL_P0_1|_RX|RB3 _PTL_P0_1|_RX|107 0  1.550338398468e-12
B_PTL_G0_1|_TX|1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|2 JJMIT AREA=2.5
B_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|5 JJMIT AREA=2.5
I_PTL_G0_1|_TX|B1 0 _PTL_G0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_1|_TX|B2 0 _PTL_G0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|3  1.684e-12
L_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|6  3.596e-12
L_PTL_G0_1|_TX|1 G0_1 _PTL_G0_1|_TX|1  2.063e-12
L_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|4  4.123e-12
L_PTL_G0_1|_TX|3 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|7  2.193e-12
R_PTL_G0_1|_TX|D _PTL_G0_1|_TX|7 _PTL_G0_1|A_PTL  1.36
L_PTL_G0_1|_TX|P1 _PTL_G0_1|_TX|2 0  5.254e-13
L_PTL_G0_1|_TX|P2 _PTL_G0_1|_TX|5 0  5.141e-13
R_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|101  2.7439617672
R_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|104  2.7439617672
L_PTL_G0_1|_TX|RB1 _PTL_G0_1|_TX|101 0  1.550338398468e-12
L_PTL_G0_1|_TX|RB2 _PTL_G0_1|_TX|104 0  1.550338398468e-12
B_PTL_G0_1|_RX|1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|5 JJMIT AREA=2.0
B_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|8 JJMIT AREA=2.5
I_PTL_G0_1|_RX|B1 0 _PTL_G0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|3  2.777e-12
I_PTL_G0_1|_RX|B2 0 _PTL_G0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|6  2.685e-12
I_PTL_G0_1|_RX|B3 0 _PTL_G0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|9  2.764e-12
L_PTL_G0_1|_RX|1 _PTL_G0_1|A_PTL _PTL_G0_1|_RX|1  1.346e-12
L_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|4  6.348e-12
L_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7  5.197e-12
L_PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7 G0_1_RX  2.058e-12
L_PTL_G0_1|_RX|P1 _PTL_G0_1|_RX|2 0  4.795e-13
L_PTL_G0_1|_RX|P2 _PTL_G0_1|_RX|5 0  5.431e-13
L_PTL_G0_1|_RX|P3 _PTL_G0_1|_RX|8 0  5.339e-13
R_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|101  4.225701121488
R_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|104  3.429952209
R_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|107  2.7439617672
L_PTL_G0_1|_RX|RB1 _PTL_G0_1|_RX|101 0  2.38752113364072e-12
L_PTL_G0_1|_RX|RB2 _PTL_G0_1|_RX|104 0  1.937922998085e-12
L_PTL_G0_1|_RX|RB3 _PTL_G0_1|_RX|107 0  1.550338398468e-12
B_PTL_G1_1|_TX|1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|2 JJMIT AREA=2.5
B_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|5 JJMIT AREA=2.5
I_PTL_G1_1|_TX|B1 0 _PTL_G1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_1|_TX|B2 0 _PTL_G1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|3  1.684e-12
L_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|6  3.596e-12
L_PTL_G1_1|_TX|1 G1_1 _PTL_G1_1|_TX|1  2.063e-12
L_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|4  4.123e-12
L_PTL_G1_1|_TX|3 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|7  2.193e-12
R_PTL_G1_1|_TX|D _PTL_G1_1|_TX|7 _PTL_G1_1|A_PTL  1.36
L_PTL_G1_1|_TX|P1 _PTL_G1_1|_TX|2 0  5.254e-13
L_PTL_G1_1|_TX|P2 _PTL_G1_1|_TX|5 0  5.141e-13
R_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|101  2.7439617672
R_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|104  2.7439617672
L_PTL_G1_1|_TX|RB1 _PTL_G1_1|_TX|101 0  1.550338398468e-12
L_PTL_G1_1|_TX|RB2 _PTL_G1_1|_TX|104 0  1.550338398468e-12
B_PTL_G1_1|_RX|1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|5 JJMIT AREA=2.0
B_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|8 JJMIT AREA=2.5
I_PTL_G1_1|_RX|B1 0 _PTL_G1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|3  2.777e-12
I_PTL_G1_1|_RX|B2 0 _PTL_G1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|6  2.685e-12
I_PTL_G1_1|_RX|B3 0 _PTL_G1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|9  2.764e-12
L_PTL_G1_1|_RX|1 _PTL_G1_1|A_PTL _PTL_G1_1|_RX|1  1.346e-12
L_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|4  6.348e-12
L_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7  5.197e-12
L_PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7 G1_1_RX  2.058e-12
L_PTL_G1_1|_RX|P1 _PTL_G1_1|_RX|2 0  4.795e-13
L_PTL_G1_1|_RX|P2 _PTL_G1_1|_RX|5 0  5.431e-13
L_PTL_G1_1|_RX|P3 _PTL_G1_1|_RX|8 0  5.339e-13
R_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|101  4.225701121488
R_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|104  3.429952209
R_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|107  2.7439617672
L_PTL_G1_1|_RX|RB1 _PTL_G1_1|_RX|101 0  2.38752113364072e-12
L_PTL_G1_1|_RX|RB2 _PTL_G1_1|_RX|104 0  1.937922998085e-12
L_PTL_G1_1|_RX|RB3 _PTL_G1_1|_RX|107 0  1.550338398468e-12
B_PTL_P2_1|_TX|1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|2 JJMIT AREA=2.5
B_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|5 JJMIT AREA=2.5
I_PTL_P2_1|_TX|B1 0 _PTL_P2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P2_1|_TX|B2 0 _PTL_P2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|3  1.684e-12
L_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|6  3.596e-12
L_PTL_P2_1|_TX|1 P2_1 _PTL_P2_1|_TX|1  2.063e-12
L_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|4  4.123e-12
L_PTL_P2_1|_TX|3 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|7  2.193e-12
R_PTL_P2_1|_TX|D _PTL_P2_1|_TX|7 _PTL_P2_1|A_PTL  1.36
L_PTL_P2_1|_TX|P1 _PTL_P2_1|_TX|2 0  5.254e-13
L_PTL_P2_1|_TX|P2 _PTL_P2_1|_TX|5 0  5.141e-13
R_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|101  2.7439617672
R_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|104  2.7439617672
L_PTL_P2_1|_TX|RB1 _PTL_P2_1|_TX|101 0  1.550338398468e-12
L_PTL_P2_1|_TX|RB2 _PTL_P2_1|_TX|104 0  1.550338398468e-12
B_PTL_P2_1|_RX|1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|5 JJMIT AREA=2.0
B_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|8 JJMIT AREA=2.5
I_PTL_P2_1|_RX|B1 0 _PTL_P2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|3  2.777e-12
I_PTL_P2_1|_RX|B2 0 _PTL_P2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|6  2.685e-12
I_PTL_P2_1|_RX|B3 0 _PTL_P2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|9  2.764e-12
L_PTL_P2_1|_RX|1 _PTL_P2_1|A_PTL _PTL_P2_1|_RX|1  1.346e-12
L_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|4  6.348e-12
L_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7  5.197e-12
L_PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7 P2_1_RX  2.058e-12
L_PTL_P2_1|_RX|P1 _PTL_P2_1|_RX|2 0  4.795e-13
L_PTL_P2_1|_RX|P2 _PTL_P2_1|_RX|5 0  5.431e-13
L_PTL_P2_1|_RX|P3 _PTL_P2_1|_RX|8 0  5.339e-13
R_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|101  4.225701121488
R_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|104  3.429952209
R_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|107  2.7439617672
L_PTL_P2_1|_RX|RB1 _PTL_P2_1|_RX|101 0  2.38752113364072e-12
L_PTL_P2_1|_RX|RB2 _PTL_P2_1|_RX|104 0  1.937922998085e-12
L_PTL_P2_1|_RX|RB3 _PTL_P2_1|_RX|107 0  1.550338398468e-12
B_PTL_G2_1|_TX|1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|2 JJMIT AREA=2.5
B_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|5 JJMIT AREA=2.5
I_PTL_G2_1|_TX|B1 0 _PTL_G2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_1|_TX|B2 0 _PTL_G2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|3  1.684e-12
L_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|6  3.596e-12
L_PTL_G2_1|_TX|1 G2_1 _PTL_G2_1|_TX|1  2.063e-12
L_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|4  4.123e-12
L_PTL_G2_1|_TX|3 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|7  2.193e-12
R_PTL_G2_1|_TX|D _PTL_G2_1|_TX|7 _PTL_G2_1|A_PTL  1.36
L_PTL_G2_1|_TX|P1 _PTL_G2_1|_TX|2 0  5.254e-13
L_PTL_G2_1|_TX|P2 _PTL_G2_1|_TX|5 0  5.141e-13
R_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|101  2.7439617672
R_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|104  2.7439617672
L_PTL_G2_1|_TX|RB1 _PTL_G2_1|_TX|101 0  1.550338398468e-12
L_PTL_G2_1|_TX|RB2 _PTL_G2_1|_TX|104 0  1.550338398468e-12
B_PTL_G2_1|_RX|1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|5 JJMIT AREA=2.0
B_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|8 JJMIT AREA=2.5
I_PTL_G2_1|_RX|B1 0 _PTL_G2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|3  2.777e-12
I_PTL_G2_1|_RX|B2 0 _PTL_G2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|6  2.685e-12
I_PTL_G2_1|_RX|B3 0 _PTL_G2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|9  2.764e-12
L_PTL_G2_1|_RX|1 _PTL_G2_1|A_PTL _PTL_G2_1|_RX|1  1.346e-12
L_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|4  6.348e-12
L_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7  5.197e-12
L_PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7 G2_1_RX  2.058e-12
L_PTL_G2_1|_RX|P1 _PTL_G2_1|_RX|2 0  4.795e-13
L_PTL_G2_1|_RX|P2 _PTL_G2_1|_RX|5 0  5.431e-13
L_PTL_G2_1|_RX|P3 _PTL_G2_1|_RX|8 0  5.339e-13
R_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|101  4.225701121488
R_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|104  3.429952209
R_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|107  2.7439617672
L_PTL_G2_1|_RX|RB1 _PTL_G2_1|_RX|101 0  2.38752113364072e-12
L_PTL_G2_1|_RX|RB2 _PTL_G2_1|_RX|104 0  1.937922998085e-12
L_PTL_G2_1|_RX|RB3 _PTL_G2_1|_RX|107 0  1.550338398468e-12
B_PTL_P3_1|_TX|1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|2 JJMIT AREA=2.5
B_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|5 JJMIT AREA=2.5
I_PTL_P3_1|_TX|B1 0 _PTL_P3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P3_1|_TX|B2 0 _PTL_P3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|3  1.684e-12
L_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|6  3.596e-12
L_PTL_P3_1|_TX|1 P3_1 _PTL_P3_1|_TX|1  2.063e-12
L_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|4  4.123e-12
L_PTL_P3_1|_TX|3 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|7  2.193e-12
R_PTL_P3_1|_TX|D _PTL_P3_1|_TX|7 _PTL_P3_1|A_PTL  1.36
L_PTL_P3_1|_TX|P1 _PTL_P3_1|_TX|2 0  5.254e-13
L_PTL_P3_1|_TX|P2 _PTL_P3_1|_TX|5 0  5.141e-13
R_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|101  2.7439617672
R_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|104  2.7439617672
L_PTL_P3_1|_TX|RB1 _PTL_P3_1|_TX|101 0  1.550338398468e-12
L_PTL_P3_1|_TX|RB2 _PTL_P3_1|_TX|104 0  1.550338398468e-12
B_PTL_P3_1|_RX|1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|5 JJMIT AREA=2.0
B_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|8 JJMIT AREA=2.5
I_PTL_P3_1|_RX|B1 0 _PTL_P3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|3  2.777e-12
I_PTL_P3_1|_RX|B2 0 _PTL_P3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|6  2.685e-12
I_PTL_P3_1|_RX|B3 0 _PTL_P3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|9  2.764e-12
L_PTL_P3_1|_RX|1 _PTL_P3_1|A_PTL _PTL_P3_1|_RX|1  1.346e-12
L_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|4  6.348e-12
L_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7  5.197e-12
L_PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7 P3_1_RX  2.058e-12
L_PTL_P3_1|_RX|P1 _PTL_P3_1|_RX|2 0  4.795e-13
L_PTL_P3_1|_RX|P2 _PTL_P3_1|_RX|5 0  5.431e-13
L_PTL_P3_1|_RX|P3 _PTL_P3_1|_RX|8 0  5.339e-13
R_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|101  4.225701121488
R_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|104  3.429952209
R_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|107  2.7439617672
L_PTL_P3_1|_RX|RB1 _PTL_P3_1|_RX|101 0  2.38752113364072e-12
L_PTL_P3_1|_RX|RB2 _PTL_P3_1|_RX|104 0  1.937922998085e-12
L_PTL_P3_1|_RX|RB3 _PTL_P3_1|_RX|107 0  1.550338398468e-12
B_PTL_G3_1|_TX|1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|2 JJMIT AREA=2.5
B_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|5 JJMIT AREA=2.5
I_PTL_G3_1|_TX|B1 0 _PTL_G3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_1|_TX|B2 0 _PTL_G3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|3  1.684e-12
L_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|6  3.596e-12
L_PTL_G3_1|_TX|1 G3_1 _PTL_G3_1|_TX|1  2.063e-12
L_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|4  4.123e-12
L_PTL_G3_1|_TX|3 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|7  2.193e-12
R_PTL_G3_1|_TX|D _PTL_G3_1|_TX|7 _PTL_G3_1|A_PTL  1.36
L_PTL_G3_1|_TX|P1 _PTL_G3_1|_TX|2 0  5.254e-13
L_PTL_G3_1|_TX|P2 _PTL_G3_1|_TX|5 0  5.141e-13
R_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|101  2.7439617672
R_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|104  2.7439617672
L_PTL_G3_1|_TX|RB1 _PTL_G3_1|_TX|101 0  1.550338398468e-12
L_PTL_G3_1|_TX|RB2 _PTL_G3_1|_TX|104 0  1.550338398468e-12
B_PTL_G3_1|_RX|1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|5 JJMIT AREA=2.0
B_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|8 JJMIT AREA=2.5
I_PTL_G3_1|_RX|B1 0 _PTL_G3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|3  2.777e-12
I_PTL_G3_1|_RX|B2 0 _PTL_G3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|6  2.685e-12
I_PTL_G3_1|_RX|B3 0 _PTL_G3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|9  2.764e-12
L_PTL_G3_1|_RX|1 _PTL_G3_1|A_PTL _PTL_G3_1|_RX|1  1.346e-12
L_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|4  6.348e-12
L_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7  5.197e-12
L_PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7 G3_1_RX  2.058e-12
L_PTL_G3_1|_RX|P1 _PTL_G3_1|_RX|2 0  4.795e-13
L_PTL_G3_1|_RX|P2 _PTL_G3_1|_RX|5 0  5.431e-13
L_PTL_G3_1|_RX|P3 _PTL_G3_1|_RX|8 0  5.339e-13
R_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|101  4.225701121488
R_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|104  3.429952209
R_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|107  2.7439617672
L_PTL_G3_1|_RX|RB1 _PTL_G3_1|_RX|101 0  2.38752113364072e-12
L_PTL_G3_1|_RX|RB2 _PTL_G3_1|_RX|104 0  1.937922998085e-12
L_PTL_G3_1|_RX|RB3 _PTL_G3_1|_RX|107 0  1.550338398468e-12
B_PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_1|_TX|B1 0 _PTL_IP1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_1|_TX|B2 0 _PTL_IP1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|3  1.684e-12
L_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|6  3.596e-12
L_PTL_IP1_1|_TX|1 IP1_1_OUT _PTL_IP1_1|_TX|1  2.063e-12
L_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|4  4.123e-12
L_PTL_IP1_1|_TX|3 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|7  2.193e-12
R_PTL_IP1_1|_TX|D _PTL_IP1_1|_TX|7 _PTL_IP1_1|A_PTL  1.36
L_PTL_IP1_1|_TX|P1 _PTL_IP1_1|_TX|2 0  5.254e-13
L_PTL_IP1_1|_TX|P2 _PTL_IP1_1|_TX|5 0  5.141e-13
R_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|101  2.7439617672
R_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|104  2.7439617672
L_PTL_IP1_1|_TX|RB1 _PTL_IP1_1|_TX|101 0  1.550338398468e-12
L_PTL_IP1_1|_TX|RB2 _PTL_IP1_1|_TX|104 0  1.550338398468e-12
B_PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_1|_RX|B1 0 _PTL_IP1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|3  2.777e-12
I_PTL_IP1_1|_RX|B2 0 _PTL_IP1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|6  2.685e-12
I_PTL_IP1_1|_RX|B3 0 _PTL_IP1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|9  2.764e-12
L_PTL_IP1_1|_RX|1 _PTL_IP1_1|A_PTL _PTL_IP1_1|_RX|1  1.346e-12
L_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|4  6.348e-12
L_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7  5.197e-12
L_PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7 IP1_1_OUT_RX  2.058e-12
L_PTL_IP1_1|_RX|P1 _PTL_IP1_1|_RX|2 0  4.795e-13
L_PTL_IP1_1|_RX|P2 _PTL_IP1_1|_RX|5 0  5.431e-13
L_PTL_IP1_1|_RX|P3 _PTL_IP1_1|_RX|8 0  5.339e-13
R_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|101  4.225701121488
R_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|104  3.429952209
R_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|107  2.7439617672
L_PTL_IP1_1|_RX|RB1 _PTL_IP1_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_1|_RX|RB2 _PTL_IP1_1|_RX|104 0  1.937922998085e-12
L_PTL_IP1_1|_RX|RB3 _PTL_IP1_1|_RX|107 0  1.550338398468e-12
B_PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_1|_TX|B1 0 _PTL_IP2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_1|_TX|B2 0 _PTL_IP2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|3  1.684e-12
L_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|6  3.596e-12
L_PTL_IP2_1|_TX|1 IP2_1_OUT _PTL_IP2_1|_TX|1  2.063e-12
L_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|4  4.123e-12
L_PTL_IP2_1|_TX|3 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|7  2.193e-12
R_PTL_IP2_1|_TX|D _PTL_IP2_1|_TX|7 _PTL_IP2_1|A_PTL  1.36
L_PTL_IP2_1|_TX|P1 _PTL_IP2_1|_TX|2 0  5.254e-13
L_PTL_IP2_1|_TX|P2 _PTL_IP2_1|_TX|5 0  5.141e-13
R_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|101  2.7439617672
R_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|104  2.7439617672
L_PTL_IP2_1|_TX|RB1 _PTL_IP2_1|_TX|101 0  1.550338398468e-12
L_PTL_IP2_1|_TX|RB2 _PTL_IP2_1|_TX|104 0  1.550338398468e-12
B_PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_1|_RX|B1 0 _PTL_IP2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|3  2.777e-12
I_PTL_IP2_1|_RX|B2 0 _PTL_IP2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|6  2.685e-12
I_PTL_IP2_1|_RX|B3 0 _PTL_IP2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|9  2.764e-12
L_PTL_IP2_1|_RX|1 _PTL_IP2_1|A_PTL _PTL_IP2_1|_RX|1  1.346e-12
L_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|4  6.348e-12
L_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7  5.197e-12
L_PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7 IP2_1_OUT_RX  2.058e-12
L_PTL_IP2_1|_RX|P1 _PTL_IP2_1|_RX|2 0  4.795e-13
L_PTL_IP2_1|_RX|P2 _PTL_IP2_1|_RX|5 0  5.431e-13
L_PTL_IP2_1|_RX|P3 _PTL_IP2_1|_RX|8 0  5.339e-13
R_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|101  4.225701121488
R_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|104  3.429952209
R_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|107  2.7439617672
L_PTL_IP2_1|_RX|RB1 _PTL_IP2_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_1|_RX|RB2 _PTL_IP2_1|_RX|104 0  1.937922998085e-12
L_PTL_IP2_1|_RX|RB3 _PTL_IP2_1|_RX|107 0  1.550338398468e-12
B_PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_1|_TX|B1 0 _PTL_IP3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_1|_TX|B2 0 _PTL_IP3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|3  1.684e-12
L_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|6  3.596e-12
L_PTL_IP3_1|_TX|1 IP3_1_OUT _PTL_IP3_1|_TX|1  2.063e-12
L_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|4  4.123e-12
L_PTL_IP3_1|_TX|3 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|7  2.193e-12
R_PTL_IP3_1|_TX|D _PTL_IP3_1|_TX|7 _PTL_IP3_1|A_PTL  1.36
L_PTL_IP3_1|_TX|P1 _PTL_IP3_1|_TX|2 0  5.254e-13
L_PTL_IP3_1|_TX|P2 _PTL_IP3_1|_TX|5 0  5.141e-13
R_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|101  2.7439617672
R_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|104  2.7439617672
L_PTL_IP3_1|_TX|RB1 _PTL_IP3_1|_TX|101 0  1.550338398468e-12
L_PTL_IP3_1|_TX|RB2 _PTL_IP3_1|_TX|104 0  1.550338398468e-12
B_PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_1|_RX|B1 0 _PTL_IP3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|3  2.777e-12
I_PTL_IP3_1|_RX|B2 0 _PTL_IP3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|6  2.685e-12
I_PTL_IP3_1|_RX|B3 0 _PTL_IP3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|9  2.764e-12
L_PTL_IP3_1|_RX|1 _PTL_IP3_1|A_PTL _PTL_IP3_1|_RX|1  1.346e-12
L_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|4  6.348e-12
L_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7  5.197e-12
L_PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7 IP3_1_OUT_RX  2.058e-12
L_PTL_IP3_1|_RX|P1 _PTL_IP3_1|_RX|2 0  4.795e-13
L_PTL_IP3_1|_RX|P2 _PTL_IP3_1|_RX|5 0  5.431e-13
L_PTL_IP3_1|_RX|P3 _PTL_IP3_1|_RX|8 0  5.339e-13
R_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|101  4.225701121488
R_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|104  3.429952209
R_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|107  2.7439617672
L_PTL_IP3_1|_RX|RB1 _PTL_IP3_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_1|_RX|RB2 _PTL_IP3_1|_RX|104 0  1.937922998085e-12
L_PTL_IP3_1|_RX|RB3 _PTL_IP3_1|_RX|107 0  1.550338398468e-12
LSPL_G1_1|SPL1|1 G1_1_RX SPL_G1_1|SPL1|D1  2e-12
LSPL_G1_1|SPL1|2 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|D2  4.135667696e-12
LSPL_G1_1|SPL1|3 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|JCT  9.84682784761905e-13
LSPL_G1_1|SPL1|4 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QA1  9.84682784761905e-13
LSPL_G1_1|SPL1|5 SPL_G1_1|SPL1|QA1 G1_1_TO1  2e-12
LSPL_G1_1|SPL1|6 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QB1  9.84682784761905e-13
LSPL_G1_1|SPL1|7 SPL_G1_1|SPL1|QB1 SPL_G1_1|QTMP  2e-12
LSPL_G1_1|SPL2|1 SPL_G1_1|QTMP SPL_G1_1|SPL2|D1  2e-12
LSPL_G1_1|SPL2|2 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|D2  4.135667696e-12
LSPL_G1_1|SPL2|3 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|JCT  9.84682784761905e-13
LSPL_G1_1|SPL2|4 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QA1  9.84682784761905e-13
LSPL_G1_1|SPL2|5 SPL_G1_1|SPL2|QA1 G1_1_TO2  2e-12
LSPL_G1_1|SPL2|6 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QB1  9.84682784761905e-13
LSPL_G1_1|SPL2|7 SPL_G1_1|SPL2|QB1 G1_1_TO3  2e-12
B_PG0_12|P|1 _PG0_12|P|1 _PG0_12|P|2 JJMIT AREA=2.5
B_PG0_12|P|2 _PG0_12|P|4 _PG0_12|P|5 JJMIT AREA=1.61
B_PG0_12|P|3 _PG0_12|P|5 _PG0_12|P|6 JJMIT AREA=1.54
B_PG0_12|P|4 _PG0_12|P|8 _PG0_12|P|9 JJMIT AREA=1.69
B_PG0_12|P|5 _PG0_12|P|10 _PG0_12|P|8 JJMIT AREA=1.38
B_PG0_12|P|6 _PG0_12|P|11 _PG0_12|P|12 JJMIT AREA=2.5
B_PG0_12|P|7 _PG0_12|P|14 _PG0_12|P|15 JJMIT AREA=2.5
I_PG0_12|P|B1 0 _PG0_12|P|3  PWL(0 0 5e-12 0.000175)
I_PG0_12|P|B2 0 _PG0_12|P|7  PWL(0 0 5e-12 0.000173)
I_PG0_12|P|B3 0 _PG0_12|P|13  PWL(0 0 5e-12 0.000175)
I_PG0_12|P|B4 0 _PG0_12|P|16  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|B1 _PG0_12|P|3 _PG0_12|P|1  2e-12
L_PG0_12|P|B2 _PG0_12|P|7 _PG0_12|P|5  2e-12
L_PG0_12|P|B3 _PG0_12|P|11 _PG0_12|P|13  2e-12
L_PG0_12|P|B4 _PG0_12|P|16 _PG0_12|P|14  2e-12
L_PG0_12|P|1 P0_1_RX _PG0_12|P|1  2.059e-12
L_PG0_12|P|2 _PG0_12|P|1 _PG0_12|P|4  4.123e-12
L_PG0_12|P|3 _PG0_12|P|5 _PG0_12|P|8  6.873e-12
L_PG0_12|P|4 _PG0_12|P|10 _PG0_12|P|11  5.195e-12
L_PG0_12|P|5 T08 _PG0_12|P|11  2.071e-12
L_PG0_12|P|6 _PG0_12|P|8 _PG0_12|P|14  3.287e-12
L_PG0_12|P|7 _PG0_12|P|14 P0_2  2.066e-12
L_PG0_12|P|P1 _PG0_12|P|2 0  5.042e-13
L_PG0_12|P|P3 _PG0_12|P|6 0  5.799e-13
L_PG0_12|P|P4 _PG0_12|P|9 0  5.733e-13
L_PG0_12|P|P6 _PG0_12|P|12 0  4.605e-13
L_PG0_12|P|P7 _PG0_12|P|15 0  4.961e-13
R_PG0_12|P|B1 _PG0_12|P|1 _PG0_12|P|101  2.7439617672
L_PG0_12|P|RB1 _PG0_12|P|101 0  1.550338398468e-12
R_PG0_12|P|B2 _PG0_12|P|4 _PG0_12|P|104  4.260810197515528
L_PG0_12|P|RB2 _PG0_12|P|104 _PG0_12|P|5  2.407357761596273e-12
R_PG0_12|P|B3 _PG0_12|P|5 _PG0_12|P|105  4.454483388311688
L_PG0_12|P|RB3 _PG0_12|P|105 0  2.516783114396104e-12
R_PG0_12|P|B4 _PG0_12|P|8 _PG0_12|P|108  4.059115040236686
L_PG0_12|P|RB4 _PG0_12|P|108 0  2.2933999977337278e-12
R_PG0_12|P|B5 _PG0_12|P|10 _PG0_12|P|110  4.970945230434783
L_PG0_12|P|RB5 _PG0_12|P|110 _PG0_12|P|8  2.8085840551956523e-12
R_PG0_12|P|B6 _PG0_12|P|11 _PG0_12|P|111  2.7439617672
L_PG0_12|P|RB6 _PG0_12|P|111 0  1.550338398468e-12
R_PG0_12|P|B7 _PG0_12|P|14 _PG0_12|P|114  2.7439617672
L_PG0_12|P|RB7 _PG0_12|P|114 0  1.550338398468e-12
B_PG0_12|G|1 _PG0_12|G|1 _PG0_12|G|2 JJMIT AREA=2.5
B_PG0_12|G|2 _PG0_12|G|4 _PG0_12|G|5 JJMIT AREA=1.61
B_PG0_12|G|3 _PG0_12|G|5 _PG0_12|G|6 JJMIT AREA=1.54
B_PG0_12|G|4 _PG0_12|G|8 _PG0_12|G|9 JJMIT AREA=1.69
B_PG0_12|G|5 _PG0_12|G|10 _PG0_12|G|8 JJMIT AREA=1.38
B_PG0_12|G|6 _PG0_12|G|11 _PG0_12|G|12 JJMIT AREA=2.5
B_PG0_12|G|7 _PG0_12|G|14 _PG0_12|G|15 JJMIT AREA=2.5
I_PG0_12|G|B1 0 _PG0_12|G|3  PWL(0 0 5e-12 0.000175)
I_PG0_12|G|B2 0 _PG0_12|G|7  PWL(0 0 5e-12 0.000173)
I_PG0_12|G|B3 0 _PG0_12|G|13  PWL(0 0 5e-12 0.000175)
I_PG0_12|G|B4 0 _PG0_12|G|16  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|B1 _PG0_12|G|3 _PG0_12|G|1  2e-12
L_PG0_12|G|B2 _PG0_12|G|7 _PG0_12|G|5  2e-12
L_PG0_12|G|B3 _PG0_12|G|11 _PG0_12|G|13  2e-12
L_PG0_12|G|B4 _PG0_12|G|16 _PG0_12|G|14  2e-12
L_PG0_12|G|1 G0_1_RX _PG0_12|G|1  2.059e-12
L_PG0_12|G|2 _PG0_12|G|1 _PG0_12|G|4  4.123e-12
L_PG0_12|G|3 _PG0_12|G|5 _PG0_12|G|8  6.873e-12
L_PG0_12|G|4 _PG0_12|G|10 _PG0_12|G|11  5.195e-12
L_PG0_12|G|5 T08 _PG0_12|G|11  2.071e-12
L_PG0_12|G|6 _PG0_12|G|8 _PG0_12|G|14  3.287e-12
L_PG0_12|G|7 _PG0_12|G|14 G0_2  2.066e-12
L_PG0_12|G|P1 _PG0_12|G|2 0  5.042e-13
L_PG0_12|G|P3 _PG0_12|G|6 0  5.799e-13
L_PG0_12|G|P4 _PG0_12|G|9 0  5.733e-13
L_PG0_12|G|P6 _PG0_12|G|12 0  4.605e-13
L_PG0_12|G|P7 _PG0_12|G|15 0  4.961e-13
R_PG0_12|G|B1 _PG0_12|G|1 _PG0_12|G|101  2.7439617672
L_PG0_12|G|RB1 _PG0_12|G|101 0  1.550338398468e-12
R_PG0_12|G|B2 _PG0_12|G|4 _PG0_12|G|104  4.260810197515528
L_PG0_12|G|RB2 _PG0_12|G|104 _PG0_12|G|5  2.407357761596273e-12
R_PG0_12|G|B3 _PG0_12|G|5 _PG0_12|G|105  4.454483388311688
L_PG0_12|G|RB3 _PG0_12|G|105 0  2.516783114396104e-12
R_PG0_12|G|B4 _PG0_12|G|8 _PG0_12|G|108  4.059115040236686
L_PG0_12|G|RB4 _PG0_12|G|108 0  2.2933999977337278e-12
R_PG0_12|G|B5 _PG0_12|G|10 _PG0_12|G|110  4.970945230434783
L_PG0_12|G|RB5 _PG0_12|G|110 _PG0_12|G|8  2.8085840551956523e-12
R_PG0_12|G|B6 _PG0_12|G|11 _PG0_12|G|111  2.7439617672
L_PG0_12|G|RB6 _PG0_12|G|111 0  1.550338398468e-12
R_PG0_12|G|B7 _PG0_12|G|14 _PG0_12|G|114  2.7439617672
L_PG0_12|G|RB7 _PG0_12|G|114 0  1.550338398468e-12
I_PG2_12|_SPL_G1|B1 0 _PG2_12|_SPL_G1|3  PWL(0 0 5e-12 0.000175)
I_PG2_12|_SPL_G1|B2 0 _PG2_12|_SPL_G1|6  PWL(0 0 5e-12 0.00028)
I_PG2_12|_SPL_G1|B3 0 _PG2_12|_SPL_G1|10  PWL(0 0 5e-12 0.000175)
I_PG2_12|_SPL_G1|B4 0 _PG2_12|_SPL_G1|13  PWL(0 0 5e-12 0.000175)
L_PG2_12|_SPL_G1|B1 _PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|1  9.175e-13
L_PG2_12|_SPL_G1|B2 _PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|4  7.666e-13
L_PG2_12|_SPL_G1|B3 _PG2_12|_SPL_G1|10 _PG2_12|_SPL_G1|8  1.928e-12
L_PG2_12|_SPL_G1|B4 _PG2_12|_SPL_G1|13 _PG2_12|_SPL_G1|11  8.786e-13
B_PG2_12|_SPL_G1|1 _PG2_12|_SPL_G1|1 _PG2_12|_SPL_G1|2 JJMIT AREA=2.5
B_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|5 JJMIT AREA=3.0
B_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|8 _PG2_12|_SPL_G1|9 JJMIT AREA=2.5
B_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|11 _PG2_12|_SPL_G1|12 JJMIT AREA=2.5
L_PG2_12|_SPL_G1|1 G2_1_RX _PG2_12|_SPL_G1|1  2.063e-12
L_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|1 _PG2_12|_SPL_G1|4  3.637e-12
L_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|7  1.278e-12
L_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|8  1.305e-12
L_PG2_12|_SPL_G1|5 _PG2_12|_SPL_G1|8 _PG2_12|G1_COPY_1  2.05e-12
L_PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|11  1.315e-12
L_PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|11 _PG2_12|G1_COPY_2  2.06e-12
L_PG2_12|_SPL_G1|P1 _PG2_12|_SPL_G1|2 0  4.676e-13
L_PG2_12|_SPL_G1|P2 _PG2_12|_SPL_G1|5 0  4.498e-13
L_PG2_12|_SPL_G1|P3 _PG2_12|_SPL_G1|9 0  5.183e-13
L_PG2_12|_SPL_G1|P4 _PG2_12|_SPL_G1|12 0  4.639e-13
R_PG2_12|_SPL_G1|B1 _PG2_12|_SPL_G1|1 _PG2_12|_SPL_G1|101  2.7439617672
L_PG2_12|_SPL_G1|RB1 _PG2_12|_SPL_G1|101 0  1.550338398468e-12
R_PG2_12|_SPL_G1|B2 _PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|104  2.286634806
L_PG2_12|_SPL_G1|RB2 _PG2_12|_SPL_G1|104 0  1.29194866539e-12
R_PG2_12|_SPL_G1|B3 _PG2_12|_SPL_G1|8 _PG2_12|_SPL_G1|108  2.7439617672
L_PG2_12|_SPL_G1|RB3 _PG2_12|_SPL_G1|108 0  1.550338398468e-12
R_PG2_12|_SPL_G1|B4 _PG2_12|_SPL_G1|11 _PG2_12|_SPL_G1|111  2.7439617672
L_PG2_12|_SPL_G1|RB4 _PG2_12|_SPL_G1|111 0  1.550338398468e-12
L_PG2_12|_PG|A1 P2_1_RX _PG2_12|_PG|A1  2.067833848e-12
L_PG2_12|_PG|A2 _PG2_12|_PG|A1 _PG2_12|_PG|A2  4.135667696e-12
L_PG2_12|_PG|A3 _PG2_12|_PG|A3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|B1 _PG2_12|G1_COPY_1 _PG2_12|_PG|B1  2.067833848e-12
L_PG2_12|_PG|B2 _PG2_12|_PG|B1 _PG2_12|_PG|B2  4.135667696e-12
L_PG2_12|_PG|B3 _PG2_12|_PG|B3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|Q3 _PG2_12|_PG|Q3 _PG2_12|_PG|Q2  4.135667696e-12
L_PG2_12|_PG|Q2 _PG2_12|_PG|Q2 _PG2_12|_PG|Q1  4.135667696e-12
L_PG2_12|_PG|Q1 _PG2_12|_PG|Q1 _PG2_12|PG  2.067833848e-12
L_PG2_12|_GG|A1 G1_1_TO2 _PG2_12|_GG|A1  2.067833848e-12
L_PG2_12|_GG|A2 _PG2_12|_GG|A1 _PG2_12|_GG|A2  4.135667696e-12
L_PG2_12|_GG|A3 _PG2_12|_GG|A3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|B1 _PG2_12|G1_COPY_2 _PG2_12|_GG|B1  2.067833848e-12
L_PG2_12|_GG|B2 _PG2_12|_GG|B1 _PG2_12|_GG|B2  4.135667696e-12
L_PG2_12|_GG|B3 _PG2_12|_GG|B3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|Q3 _PG2_12|_GG|Q3 _PG2_12|_GG|Q2  4.135667696e-12
L_PG2_12|_GG|Q2 _PG2_12|_GG|Q2 _PG2_12|_GG|Q1  4.135667696e-12
L_PG2_12|_GG|Q1 _PG2_12|_GG|Q1 _PG2_12|GG  2.067833848e-12
B_PG2_12|_DFF_PG|1 _PG2_12|_DFF_PG|1 _PG2_12|_DFF_PG|2 JJMIT AREA=2.5
B_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|5 JJMIT AREA=1.61
B_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|6 JJMIT AREA=1.54
B_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|8 _PG2_12|_DFF_PG|9 JJMIT AREA=1.69
B_PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|10 _PG2_12|_DFF_PG|8 JJMIT AREA=1.38
B_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|11 _PG2_12|_DFF_PG|12 JJMIT AREA=2.5
B_PG2_12|_DFF_PG|7 _PG2_12|_DFF_PG|14 _PG2_12|_DFF_PG|15 JJMIT AREA=2.5
I_PG2_12|_DFF_PG|B1 0 _PG2_12|_DFF_PG|3  PWL(0 0 5e-12 0.000175)
I_PG2_12|_DFF_PG|B2 0 _PG2_12|_DFF_PG|7  PWL(0 0 5e-12 0.000173)
I_PG2_12|_DFF_PG|B3 0 _PG2_12|_DFF_PG|13  PWL(0 0 5e-12 0.000175)
I_PG2_12|_DFF_PG|B4 0 _PG2_12|_DFF_PG|16  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|B1 _PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|1  2e-12
L_PG2_12|_DFF_PG|B2 _PG2_12|_DFF_PG|7 _PG2_12|_DFF_PG|5  2e-12
L_PG2_12|_DFF_PG|B3 _PG2_12|_DFF_PG|11 _PG2_12|_DFF_PG|13  2e-12
L_PG2_12|_DFF_PG|B4 _PG2_12|_DFF_PG|16 _PG2_12|_DFF_PG|14  2e-12
L_PG2_12|_DFF_PG|1 _PG2_12|PG _PG2_12|_DFF_PG|1  2.059e-12
L_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|1 _PG2_12|_DFF_PG|4  4.123e-12
L_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|8  6.873e-12
L_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|10 _PG2_12|_DFF_PG|11  5.195e-12
L_PG2_12|_DFF_PG|5 T10 _PG2_12|_DFF_PG|11  2.071e-12
L_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|8 _PG2_12|_DFF_PG|14  3.287e-12
L_PG2_12|_DFF_PG|7 _PG2_12|_DFF_PG|14 _PG2_12|PG_SYNC  2.066e-12
L_PG2_12|_DFF_PG|P1 _PG2_12|_DFF_PG|2 0  5.042e-13
L_PG2_12|_DFF_PG|P3 _PG2_12|_DFF_PG|6 0  5.799e-13
L_PG2_12|_DFF_PG|P4 _PG2_12|_DFF_PG|9 0  5.733e-13
L_PG2_12|_DFF_PG|P6 _PG2_12|_DFF_PG|12 0  4.605e-13
L_PG2_12|_DFF_PG|P7 _PG2_12|_DFF_PG|15 0  4.961e-13
R_PG2_12|_DFF_PG|B1 _PG2_12|_DFF_PG|1 _PG2_12|_DFF_PG|101  2.7439617672
L_PG2_12|_DFF_PG|RB1 _PG2_12|_DFF_PG|101 0  1.550338398468e-12
R_PG2_12|_DFF_PG|B2 _PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|104  4.260810197515528
L_PG2_12|_DFF_PG|RB2 _PG2_12|_DFF_PG|104 _PG2_12|_DFF_PG|5  2.407357761596273e-12
R_PG2_12|_DFF_PG|B3 _PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|105  4.454483388311688
L_PG2_12|_DFF_PG|RB3 _PG2_12|_DFF_PG|105 0  2.516783114396104e-12
R_PG2_12|_DFF_PG|B4 _PG2_12|_DFF_PG|8 _PG2_12|_DFF_PG|108  4.059115040236686
L_PG2_12|_DFF_PG|RB4 _PG2_12|_DFF_PG|108 0  2.2933999977337278e-12
R_PG2_12|_DFF_PG|B5 _PG2_12|_DFF_PG|10 _PG2_12|_DFF_PG|110  4.970945230434783
L_PG2_12|_DFF_PG|RB5 _PG2_12|_DFF_PG|110 _PG2_12|_DFF_PG|8  2.8085840551956523e-12
R_PG2_12|_DFF_PG|B6 _PG2_12|_DFF_PG|11 _PG2_12|_DFF_PG|111  2.7439617672
L_PG2_12|_DFF_PG|RB6 _PG2_12|_DFF_PG|111 0  1.550338398468e-12
R_PG2_12|_DFF_PG|B7 _PG2_12|_DFF_PG|14 _PG2_12|_DFF_PG|114  2.7439617672
L_PG2_12|_DFF_PG|RB7 _PG2_12|_DFF_PG|114 0  1.550338398468e-12
B_PG2_12|_DFF_GG|1 _PG2_12|_DFF_GG|1 _PG2_12|_DFF_GG|2 JJMIT AREA=2.5
B_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|5 JJMIT AREA=1.61
B_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|6 JJMIT AREA=1.54
B_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|8 _PG2_12|_DFF_GG|9 JJMIT AREA=1.69
B_PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|10 _PG2_12|_DFF_GG|8 JJMIT AREA=1.38
B_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|11 _PG2_12|_DFF_GG|12 JJMIT AREA=2.5
B_PG2_12|_DFF_GG|7 _PG2_12|_DFF_GG|14 _PG2_12|_DFF_GG|15 JJMIT AREA=2.5
I_PG2_12|_DFF_GG|B1 0 _PG2_12|_DFF_GG|3  PWL(0 0 5e-12 0.000175)
I_PG2_12|_DFF_GG|B2 0 _PG2_12|_DFF_GG|7  PWL(0 0 5e-12 0.000173)
I_PG2_12|_DFF_GG|B3 0 _PG2_12|_DFF_GG|13  PWL(0 0 5e-12 0.000175)
I_PG2_12|_DFF_GG|B4 0 _PG2_12|_DFF_GG|16  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|B1 _PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|1  2e-12
L_PG2_12|_DFF_GG|B2 _PG2_12|_DFF_GG|7 _PG2_12|_DFF_GG|5  2e-12
L_PG2_12|_DFF_GG|B3 _PG2_12|_DFF_GG|11 _PG2_12|_DFF_GG|13  2e-12
L_PG2_12|_DFF_GG|B4 _PG2_12|_DFF_GG|16 _PG2_12|_DFF_GG|14  2e-12
L_PG2_12|_DFF_GG|1 _PG2_12|GG _PG2_12|_DFF_GG|1  2.059e-12
L_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|1 _PG2_12|_DFF_GG|4  4.123e-12
L_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|8  6.873e-12
L_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|10 _PG2_12|_DFF_GG|11  5.195e-12
L_PG2_12|_DFF_GG|5 T10 _PG2_12|_DFF_GG|11  2.071e-12
L_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|8 _PG2_12|_DFF_GG|14  3.287e-12
L_PG2_12|_DFF_GG|7 _PG2_12|_DFF_GG|14 _PG2_12|GG_SYNC  2.066e-12
L_PG2_12|_DFF_GG|P1 _PG2_12|_DFF_GG|2 0  5.042e-13
L_PG2_12|_DFF_GG|P3 _PG2_12|_DFF_GG|6 0  5.799e-13
L_PG2_12|_DFF_GG|P4 _PG2_12|_DFF_GG|9 0  5.733e-13
L_PG2_12|_DFF_GG|P6 _PG2_12|_DFF_GG|12 0  4.605e-13
L_PG2_12|_DFF_GG|P7 _PG2_12|_DFF_GG|15 0  4.961e-13
R_PG2_12|_DFF_GG|B1 _PG2_12|_DFF_GG|1 _PG2_12|_DFF_GG|101  2.7439617672
L_PG2_12|_DFF_GG|RB1 _PG2_12|_DFF_GG|101 0  1.550338398468e-12
R_PG2_12|_DFF_GG|B2 _PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|104  4.260810197515528
L_PG2_12|_DFF_GG|RB2 _PG2_12|_DFF_GG|104 _PG2_12|_DFF_GG|5  2.407357761596273e-12
R_PG2_12|_DFF_GG|B3 _PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|105  4.454483388311688
L_PG2_12|_DFF_GG|RB3 _PG2_12|_DFF_GG|105 0  2.516783114396104e-12
R_PG2_12|_DFF_GG|B4 _PG2_12|_DFF_GG|8 _PG2_12|_DFF_GG|108  4.059115040236686
L_PG2_12|_DFF_GG|RB4 _PG2_12|_DFF_GG|108 0  2.2933999977337278e-12
R_PG2_12|_DFF_GG|B5 _PG2_12|_DFF_GG|10 _PG2_12|_DFF_GG|110  4.970945230434783
L_PG2_12|_DFF_GG|RB5 _PG2_12|_DFF_GG|110 _PG2_12|_DFF_GG|8  2.8085840551956523e-12
R_PG2_12|_DFF_GG|B6 _PG2_12|_DFF_GG|11 _PG2_12|_DFF_GG|111  2.7439617672
L_PG2_12|_DFF_GG|RB6 _PG2_12|_DFF_GG|111 0  1.550338398468e-12
R_PG2_12|_DFF_GG|B7 _PG2_12|_DFF_GG|14 _PG2_12|_DFF_GG|114  2.7439617672
L_PG2_12|_DFF_GG|RB7 _PG2_12|_DFF_GG|114 0  1.550338398468e-12
L_PG2_12|_AND_G|A1 _PG2_12|PG_SYNC _PG2_12|_AND_G|A1  2.067833848e-12
L_PG2_12|_AND_G|A2 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A2  4.135667696e-12
L_PG2_12|_AND_G|A3 _PG2_12|_AND_G|A3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|B1 _PG2_12|GG_SYNC _PG2_12|_AND_G|B1  2.067833848e-12
L_PG2_12|_AND_G|B2 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B2  4.135667696e-12
L_PG2_12|_AND_G|B3 _PG2_12|_AND_G|B3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q2  4.135667696e-12
L_PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q1  4.135667696e-12
L_PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1 G2_2  2.067833848e-12
I_PG3_12|_SPL_G1|B1 0 _PG3_12|_SPL_G1|3  PWL(0 0 5e-12 0.000175)
I_PG3_12|_SPL_G1|B2 0 _PG3_12|_SPL_G1|6  PWL(0 0 5e-12 0.00028)
I_PG3_12|_SPL_G1|B3 0 _PG3_12|_SPL_G1|10  PWL(0 0 5e-12 0.000175)
I_PG3_12|_SPL_G1|B4 0 _PG3_12|_SPL_G1|13  PWL(0 0 5e-12 0.000175)
L_PG3_12|_SPL_G1|B1 _PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|1  9.175e-13
L_PG3_12|_SPL_G1|B2 _PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|4  7.666e-13
L_PG3_12|_SPL_G1|B3 _PG3_12|_SPL_G1|10 _PG3_12|_SPL_G1|8  1.928e-12
L_PG3_12|_SPL_G1|B4 _PG3_12|_SPL_G1|13 _PG3_12|_SPL_G1|11  8.786e-13
B_PG3_12|_SPL_G1|1 _PG3_12|_SPL_G1|1 _PG3_12|_SPL_G1|2 JJMIT AREA=2.5
B_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|5 JJMIT AREA=3.0
B_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|8 _PG3_12|_SPL_G1|9 JJMIT AREA=2.5
B_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|11 _PG3_12|_SPL_G1|12 JJMIT AREA=2.5
L_PG3_12|_SPL_G1|1 G3_1_RX _PG3_12|_SPL_G1|1  2.063e-12
L_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|1 _PG3_12|_SPL_G1|4  3.637e-12
L_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|7  1.278e-12
L_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|8  1.305e-12
L_PG3_12|_SPL_G1|5 _PG3_12|_SPL_G1|8 _PG3_12|G1_COPY_1  2.05e-12
L_PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|11  1.315e-12
L_PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|11 _PG3_12|G1_COPY_2  2.06e-12
L_PG3_12|_SPL_G1|P1 _PG3_12|_SPL_G1|2 0  4.676e-13
L_PG3_12|_SPL_G1|P2 _PG3_12|_SPL_G1|5 0  4.498e-13
L_PG3_12|_SPL_G1|P3 _PG3_12|_SPL_G1|9 0  5.183e-13
L_PG3_12|_SPL_G1|P4 _PG3_12|_SPL_G1|12 0  4.639e-13
R_PG3_12|_SPL_G1|B1 _PG3_12|_SPL_G1|1 _PG3_12|_SPL_G1|101  2.7439617672
L_PG3_12|_SPL_G1|RB1 _PG3_12|_SPL_G1|101 0  1.550338398468e-12
R_PG3_12|_SPL_G1|B2 _PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|104  2.286634806
L_PG3_12|_SPL_G1|RB2 _PG3_12|_SPL_G1|104 0  1.29194866539e-12
R_PG3_12|_SPL_G1|B3 _PG3_12|_SPL_G1|8 _PG3_12|_SPL_G1|108  2.7439617672
L_PG3_12|_SPL_G1|RB3 _PG3_12|_SPL_G1|108 0  1.550338398468e-12
R_PG3_12|_SPL_G1|B4 _PG3_12|_SPL_G1|11 _PG3_12|_SPL_G1|111  2.7439617672
L_PG3_12|_SPL_G1|RB4 _PG3_12|_SPL_G1|111 0  1.550338398468e-12
L_PG3_12|_PG|A1 P3_1_RX _PG3_12|_PG|A1  2.067833848e-12
L_PG3_12|_PG|A2 _PG3_12|_PG|A1 _PG3_12|_PG|A2  4.135667696e-12
L_PG3_12|_PG|A3 _PG3_12|_PG|A3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|B1 _PG3_12|G1_COPY_1 _PG3_12|_PG|B1  2.067833848e-12
L_PG3_12|_PG|B2 _PG3_12|_PG|B1 _PG3_12|_PG|B2  4.135667696e-12
L_PG3_12|_PG|B3 _PG3_12|_PG|B3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|Q3 _PG3_12|_PG|Q3 _PG3_12|_PG|Q2  4.135667696e-12
L_PG3_12|_PG|Q2 _PG3_12|_PG|Q2 _PG3_12|_PG|Q1  4.135667696e-12
L_PG3_12|_PG|Q1 _PG3_12|_PG|Q1 _PG3_12|PG  2.067833848e-12
L_PG3_12|_GG|A1 G1_1_TO3 _PG3_12|_GG|A1  2.067833848e-12
L_PG3_12|_GG|A2 _PG3_12|_GG|A1 _PG3_12|_GG|A2  4.135667696e-12
L_PG3_12|_GG|A3 _PG3_12|_GG|A3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|B1 _PG3_12|G1_COPY_2 _PG3_12|_GG|B1  2.067833848e-12
L_PG3_12|_GG|B2 _PG3_12|_GG|B1 _PG3_12|_GG|B2  4.135667696e-12
L_PG3_12|_GG|B3 _PG3_12|_GG|B3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|Q3 _PG3_12|_GG|Q3 _PG3_12|_GG|Q2  4.135667696e-12
L_PG3_12|_GG|Q2 _PG3_12|_GG|Q2 _PG3_12|_GG|Q1  4.135667696e-12
L_PG3_12|_GG|Q1 _PG3_12|_GG|Q1 _PG3_12|GG  2.067833848e-12
B_PG3_12|_DFF_PG|1 _PG3_12|_DFF_PG|1 _PG3_12|_DFF_PG|2 JJMIT AREA=2.5
B_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|5 JJMIT AREA=1.61
B_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|6 JJMIT AREA=1.54
B_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|8 _PG3_12|_DFF_PG|9 JJMIT AREA=1.69
B_PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|10 _PG3_12|_DFF_PG|8 JJMIT AREA=1.38
B_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|11 _PG3_12|_DFF_PG|12 JJMIT AREA=2.5
B_PG3_12|_DFF_PG|7 _PG3_12|_DFF_PG|14 _PG3_12|_DFF_PG|15 JJMIT AREA=2.5
I_PG3_12|_DFF_PG|B1 0 _PG3_12|_DFF_PG|3  PWL(0 0 5e-12 0.000175)
I_PG3_12|_DFF_PG|B2 0 _PG3_12|_DFF_PG|7  PWL(0 0 5e-12 0.000173)
I_PG3_12|_DFF_PG|B3 0 _PG3_12|_DFF_PG|13  PWL(0 0 5e-12 0.000175)
I_PG3_12|_DFF_PG|B4 0 _PG3_12|_DFF_PG|16  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|B1 _PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|1  2e-12
L_PG3_12|_DFF_PG|B2 _PG3_12|_DFF_PG|7 _PG3_12|_DFF_PG|5  2e-12
L_PG3_12|_DFF_PG|B3 _PG3_12|_DFF_PG|11 _PG3_12|_DFF_PG|13  2e-12
L_PG3_12|_DFF_PG|B4 _PG3_12|_DFF_PG|16 _PG3_12|_DFF_PG|14  2e-12
L_PG3_12|_DFF_PG|1 _PG3_12|PG _PG3_12|_DFF_PG|1  2.059e-12
L_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|1 _PG3_12|_DFF_PG|4  4.123e-12
L_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|8  6.873e-12
L_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|10 _PG3_12|_DFF_PG|11  5.195e-12
L_PG3_12|_DFF_PG|5 T11 _PG3_12|_DFF_PG|11  2.071e-12
L_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|8 _PG3_12|_DFF_PG|14  3.287e-12
L_PG3_12|_DFF_PG|7 _PG3_12|_DFF_PG|14 _PG3_12|PG_SYNC  2.066e-12
L_PG3_12|_DFF_PG|P1 _PG3_12|_DFF_PG|2 0  5.042e-13
L_PG3_12|_DFF_PG|P3 _PG3_12|_DFF_PG|6 0  5.799e-13
L_PG3_12|_DFF_PG|P4 _PG3_12|_DFF_PG|9 0  5.733e-13
L_PG3_12|_DFF_PG|P6 _PG3_12|_DFF_PG|12 0  4.605e-13
L_PG3_12|_DFF_PG|P7 _PG3_12|_DFF_PG|15 0  4.961e-13
R_PG3_12|_DFF_PG|B1 _PG3_12|_DFF_PG|1 _PG3_12|_DFF_PG|101  2.7439617672
L_PG3_12|_DFF_PG|RB1 _PG3_12|_DFF_PG|101 0  1.550338398468e-12
R_PG3_12|_DFF_PG|B2 _PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|104  4.260810197515528
L_PG3_12|_DFF_PG|RB2 _PG3_12|_DFF_PG|104 _PG3_12|_DFF_PG|5  2.407357761596273e-12
R_PG3_12|_DFF_PG|B3 _PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|105  4.454483388311688
L_PG3_12|_DFF_PG|RB3 _PG3_12|_DFF_PG|105 0  2.516783114396104e-12
R_PG3_12|_DFF_PG|B4 _PG3_12|_DFF_PG|8 _PG3_12|_DFF_PG|108  4.059115040236686
L_PG3_12|_DFF_PG|RB4 _PG3_12|_DFF_PG|108 0  2.2933999977337278e-12
R_PG3_12|_DFF_PG|B5 _PG3_12|_DFF_PG|10 _PG3_12|_DFF_PG|110  4.970945230434783
L_PG3_12|_DFF_PG|RB5 _PG3_12|_DFF_PG|110 _PG3_12|_DFF_PG|8  2.8085840551956523e-12
R_PG3_12|_DFF_PG|B6 _PG3_12|_DFF_PG|11 _PG3_12|_DFF_PG|111  2.7439617672
L_PG3_12|_DFF_PG|RB6 _PG3_12|_DFF_PG|111 0  1.550338398468e-12
R_PG3_12|_DFF_PG|B7 _PG3_12|_DFF_PG|14 _PG3_12|_DFF_PG|114  2.7439617672
L_PG3_12|_DFF_PG|RB7 _PG3_12|_DFF_PG|114 0  1.550338398468e-12
B_PG3_12|_DFF_GG|1 _PG3_12|_DFF_GG|1 _PG3_12|_DFF_GG|2 JJMIT AREA=2.5
B_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|5 JJMIT AREA=1.61
B_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|6 JJMIT AREA=1.54
B_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|8 _PG3_12|_DFF_GG|9 JJMIT AREA=1.69
B_PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|10 _PG3_12|_DFF_GG|8 JJMIT AREA=1.38
B_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|11 _PG3_12|_DFF_GG|12 JJMIT AREA=2.5
B_PG3_12|_DFF_GG|7 _PG3_12|_DFF_GG|14 _PG3_12|_DFF_GG|15 JJMIT AREA=2.5
I_PG3_12|_DFF_GG|B1 0 _PG3_12|_DFF_GG|3  PWL(0 0 5e-12 0.000175)
I_PG3_12|_DFF_GG|B2 0 _PG3_12|_DFF_GG|7  PWL(0 0 5e-12 0.000173)
I_PG3_12|_DFF_GG|B3 0 _PG3_12|_DFF_GG|13  PWL(0 0 5e-12 0.000175)
I_PG3_12|_DFF_GG|B4 0 _PG3_12|_DFF_GG|16  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|B1 _PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|1  2e-12
L_PG3_12|_DFF_GG|B2 _PG3_12|_DFF_GG|7 _PG3_12|_DFF_GG|5  2e-12
L_PG3_12|_DFF_GG|B3 _PG3_12|_DFF_GG|11 _PG3_12|_DFF_GG|13  2e-12
L_PG3_12|_DFF_GG|B4 _PG3_12|_DFF_GG|16 _PG3_12|_DFF_GG|14  2e-12
L_PG3_12|_DFF_GG|1 _PG3_12|GG _PG3_12|_DFF_GG|1  2.059e-12
L_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|1 _PG3_12|_DFF_GG|4  4.123e-12
L_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|8  6.873e-12
L_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|10 _PG3_12|_DFF_GG|11  5.195e-12
L_PG3_12|_DFF_GG|5 T11 _PG3_12|_DFF_GG|11  2.071e-12
L_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|8 _PG3_12|_DFF_GG|14  3.287e-12
L_PG3_12|_DFF_GG|7 _PG3_12|_DFF_GG|14 _PG3_12|GG_SYNC  2.066e-12
L_PG3_12|_DFF_GG|P1 _PG3_12|_DFF_GG|2 0  5.042e-13
L_PG3_12|_DFF_GG|P3 _PG3_12|_DFF_GG|6 0  5.799e-13
L_PG3_12|_DFF_GG|P4 _PG3_12|_DFF_GG|9 0  5.733e-13
L_PG3_12|_DFF_GG|P6 _PG3_12|_DFF_GG|12 0  4.605e-13
L_PG3_12|_DFF_GG|P7 _PG3_12|_DFF_GG|15 0  4.961e-13
R_PG3_12|_DFF_GG|B1 _PG3_12|_DFF_GG|1 _PG3_12|_DFF_GG|101  2.7439617672
L_PG3_12|_DFF_GG|RB1 _PG3_12|_DFF_GG|101 0  1.550338398468e-12
R_PG3_12|_DFF_GG|B2 _PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|104  4.260810197515528
L_PG3_12|_DFF_GG|RB2 _PG3_12|_DFF_GG|104 _PG3_12|_DFF_GG|5  2.407357761596273e-12
R_PG3_12|_DFF_GG|B3 _PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|105  4.454483388311688
L_PG3_12|_DFF_GG|RB3 _PG3_12|_DFF_GG|105 0  2.516783114396104e-12
R_PG3_12|_DFF_GG|B4 _PG3_12|_DFF_GG|8 _PG3_12|_DFF_GG|108  4.059115040236686
L_PG3_12|_DFF_GG|RB4 _PG3_12|_DFF_GG|108 0  2.2933999977337278e-12
R_PG3_12|_DFF_GG|B5 _PG3_12|_DFF_GG|10 _PG3_12|_DFF_GG|110  4.970945230434783
L_PG3_12|_DFF_GG|RB5 _PG3_12|_DFF_GG|110 _PG3_12|_DFF_GG|8  2.8085840551956523e-12
R_PG3_12|_DFF_GG|B6 _PG3_12|_DFF_GG|11 _PG3_12|_DFF_GG|111  2.7439617672
L_PG3_12|_DFF_GG|RB6 _PG3_12|_DFF_GG|111 0  1.550338398468e-12
R_PG3_12|_DFF_GG|B7 _PG3_12|_DFF_GG|14 _PG3_12|_DFF_GG|114  2.7439617672
L_PG3_12|_DFF_GG|RB7 _PG3_12|_DFF_GG|114 0  1.550338398468e-12
L_PG3_12|_AND_G|A1 _PG3_12|PG_SYNC _PG3_12|_AND_G|A1  2.067833848e-12
L_PG3_12|_AND_G|A2 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A2  4.135667696e-12
L_PG3_12|_AND_G|A3 _PG3_12|_AND_G|A3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|B1 _PG3_12|GG_SYNC _PG3_12|_AND_G|B1  2.067833848e-12
L_PG3_12|_AND_G|B2 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B2  4.135667696e-12
L_PG3_12|_AND_G|B3 _PG3_12|_AND_G|B3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q2  4.135667696e-12
L_PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q1  4.135667696e-12
L_PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1 G3_2  2.067833848e-12
B_PTL_P0_2|_TX|1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|2 JJMIT AREA=2.5
B_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|5 JJMIT AREA=2.5
I_PTL_P0_2|_TX|B1 0 _PTL_P0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_2|_TX|B2 0 _PTL_P0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|3  1.684e-12
L_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|6  3.596e-12
L_PTL_P0_2|_TX|1 P0_2 _PTL_P0_2|_TX|1  2.063e-12
L_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|4  4.123e-12
L_PTL_P0_2|_TX|3 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|7  2.193e-12
R_PTL_P0_2|_TX|D _PTL_P0_2|_TX|7 _PTL_P0_2|A_PTL  1.36
L_PTL_P0_2|_TX|P1 _PTL_P0_2|_TX|2 0  5.254e-13
L_PTL_P0_2|_TX|P2 _PTL_P0_2|_TX|5 0  5.141e-13
R_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|101  2.7439617672
R_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|104  2.7439617672
L_PTL_P0_2|_TX|RB1 _PTL_P0_2|_TX|101 0  1.550338398468e-12
L_PTL_P0_2|_TX|RB2 _PTL_P0_2|_TX|104 0  1.550338398468e-12
B_PTL_P0_2|_RX|1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|5 JJMIT AREA=2.0
B_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|8 JJMIT AREA=2.5
I_PTL_P0_2|_RX|B1 0 _PTL_P0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|3  2.777e-12
I_PTL_P0_2|_RX|B2 0 _PTL_P0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|6  2.685e-12
I_PTL_P0_2|_RX|B3 0 _PTL_P0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|9  2.764e-12
L_PTL_P0_2|_RX|1 _PTL_P0_2|A_PTL _PTL_P0_2|_RX|1  1.346e-12
L_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|4  6.348e-12
L_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7  5.197e-12
L_PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7 P0_2_RX  2.058e-12
L_PTL_P0_2|_RX|P1 _PTL_P0_2|_RX|2 0  4.795e-13
L_PTL_P0_2|_RX|P2 _PTL_P0_2|_RX|5 0  5.431e-13
L_PTL_P0_2|_RX|P3 _PTL_P0_2|_RX|8 0  5.339e-13
R_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|101  4.225701121488
R_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|104  3.429952209
R_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|107  2.7439617672
L_PTL_P0_2|_RX|RB1 _PTL_P0_2|_RX|101 0  2.38752113364072e-12
L_PTL_P0_2|_RX|RB2 _PTL_P0_2|_RX|104 0  1.937922998085e-12
L_PTL_P0_2|_RX|RB3 _PTL_P0_2|_RX|107 0  1.550338398468e-12
B_PTL_G0_2|_TX|1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|2 JJMIT AREA=2.5
B_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|5 JJMIT AREA=2.5
I_PTL_G0_2|_TX|B1 0 _PTL_G0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_2|_TX|B2 0 _PTL_G0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|3  1.684e-12
L_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|6  3.596e-12
L_PTL_G0_2|_TX|1 G0_2 _PTL_G0_2|_TX|1  2.063e-12
L_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|4  4.123e-12
L_PTL_G0_2|_TX|3 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|7  2.193e-12
R_PTL_G0_2|_TX|D _PTL_G0_2|_TX|7 _PTL_G0_2|A_PTL  1.36
L_PTL_G0_2|_TX|P1 _PTL_G0_2|_TX|2 0  5.254e-13
L_PTL_G0_2|_TX|P2 _PTL_G0_2|_TX|5 0  5.141e-13
R_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|101  2.7439617672
R_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|104  2.7439617672
L_PTL_G0_2|_TX|RB1 _PTL_G0_2|_TX|101 0  1.550338398468e-12
L_PTL_G0_2|_TX|RB2 _PTL_G0_2|_TX|104 0  1.550338398468e-12
B_PTL_G0_2|_RX|1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|5 JJMIT AREA=2.0
B_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|8 JJMIT AREA=2.5
I_PTL_G0_2|_RX|B1 0 _PTL_G0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|3  2.777e-12
I_PTL_G0_2|_RX|B2 0 _PTL_G0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|6  2.685e-12
I_PTL_G0_2|_RX|B3 0 _PTL_G0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|9  2.764e-12
L_PTL_G0_2|_RX|1 _PTL_G0_2|A_PTL _PTL_G0_2|_RX|1  1.346e-12
L_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|4  6.348e-12
L_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7  5.197e-12
L_PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7 G0_2_RX  2.058e-12
L_PTL_G0_2|_RX|P1 _PTL_G0_2|_RX|2 0  4.795e-13
L_PTL_G0_2|_RX|P2 _PTL_G0_2|_RX|5 0  5.431e-13
L_PTL_G0_2|_RX|P3 _PTL_G0_2|_RX|8 0  5.339e-13
R_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|101  4.225701121488
R_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|104  3.429952209
R_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|107  2.7439617672
L_PTL_G0_2|_RX|RB1 _PTL_G0_2|_RX|101 0  2.38752113364072e-12
L_PTL_G0_2|_RX|RB2 _PTL_G0_2|_RX|104 0  1.937922998085e-12
L_PTL_G0_2|_RX|RB3 _PTL_G0_2|_RX|107 0  1.550338398468e-12
B_PTL_G1_2|_TX|1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|2 JJMIT AREA=2.5
B_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|5 JJMIT AREA=2.5
I_PTL_G1_2|_TX|B1 0 _PTL_G1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_2|_TX|B2 0 _PTL_G1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|3  1.684e-12
L_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|6  3.596e-12
L_PTL_G1_2|_TX|1 G1_2 _PTL_G1_2|_TX|1  2.063e-12
L_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|4  4.123e-12
L_PTL_G1_2|_TX|3 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|7  2.193e-12
R_PTL_G1_2|_TX|D _PTL_G1_2|_TX|7 _PTL_G1_2|A_PTL  1.36
L_PTL_G1_2|_TX|P1 _PTL_G1_2|_TX|2 0  5.254e-13
L_PTL_G1_2|_TX|P2 _PTL_G1_2|_TX|5 0  5.141e-13
R_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|101  2.7439617672
R_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|104  2.7439617672
L_PTL_G1_2|_TX|RB1 _PTL_G1_2|_TX|101 0  1.550338398468e-12
L_PTL_G1_2|_TX|RB2 _PTL_G1_2|_TX|104 0  1.550338398468e-12
B_PTL_G1_2|_RX|1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|5 JJMIT AREA=2.0
B_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|8 JJMIT AREA=2.5
I_PTL_G1_2|_RX|B1 0 _PTL_G1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|3  2.777e-12
I_PTL_G1_2|_RX|B2 0 _PTL_G1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|6  2.685e-12
I_PTL_G1_2|_RX|B3 0 _PTL_G1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|9  2.764e-12
L_PTL_G1_2|_RX|1 _PTL_G1_2|A_PTL _PTL_G1_2|_RX|1  1.346e-12
L_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|4  6.348e-12
L_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7  5.197e-12
L_PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7 G1_2_RX  2.058e-12
L_PTL_G1_2|_RX|P1 _PTL_G1_2|_RX|2 0  4.795e-13
L_PTL_G1_2|_RX|P2 _PTL_G1_2|_RX|5 0  5.431e-13
L_PTL_G1_2|_RX|P3 _PTL_G1_2|_RX|8 0  5.339e-13
R_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|101  4.225701121488
R_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|104  3.429952209
R_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|107  2.7439617672
L_PTL_G1_2|_RX|RB1 _PTL_G1_2|_RX|101 0  2.38752113364072e-12
L_PTL_G1_2|_RX|RB2 _PTL_G1_2|_RX|104 0  1.937922998085e-12
L_PTL_G1_2|_RX|RB3 _PTL_G1_2|_RX|107 0  1.550338398468e-12
B_PTL_G2_2|_TX|1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|2 JJMIT AREA=2.5
B_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|5 JJMIT AREA=2.5
I_PTL_G2_2|_TX|B1 0 _PTL_G2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_2|_TX|B2 0 _PTL_G2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|3  1.684e-12
L_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|6  3.596e-12
L_PTL_G2_2|_TX|1 G2_2 _PTL_G2_2|_TX|1  2.063e-12
L_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|4  4.123e-12
L_PTL_G2_2|_TX|3 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|7  2.193e-12
R_PTL_G2_2|_TX|D _PTL_G2_2|_TX|7 _PTL_G2_2|A_PTL  1.36
L_PTL_G2_2|_TX|P1 _PTL_G2_2|_TX|2 0  5.254e-13
L_PTL_G2_2|_TX|P2 _PTL_G2_2|_TX|5 0  5.141e-13
R_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|101  2.7439617672
R_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|104  2.7439617672
L_PTL_G2_2|_TX|RB1 _PTL_G2_2|_TX|101 0  1.550338398468e-12
L_PTL_G2_2|_TX|RB2 _PTL_G2_2|_TX|104 0  1.550338398468e-12
B_PTL_G2_2|_RX|1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|5 JJMIT AREA=2.0
B_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|8 JJMIT AREA=2.5
I_PTL_G2_2|_RX|B1 0 _PTL_G2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|3  2.777e-12
I_PTL_G2_2|_RX|B2 0 _PTL_G2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|6  2.685e-12
I_PTL_G2_2|_RX|B3 0 _PTL_G2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|9  2.764e-12
L_PTL_G2_2|_RX|1 _PTL_G2_2|A_PTL _PTL_G2_2|_RX|1  1.346e-12
L_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|4  6.348e-12
L_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7  5.197e-12
L_PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7 G2_2_RX  2.058e-12
L_PTL_G2_2|_RX|P1 _PTL_G2_2|_RX|2 0  4.795e-13
L_PTL_G2_2|_RX|P2 _PTL_G2_2|_RX|5 0  5.431e-13
L_PTL_G2_2|_RX|P3 _PTL_G2_2|_RX|8 0  5.339e-13
R_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|101  4.225701121488
R_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|104  3.429952209
R_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|107  2.7439617672
L_PTL_G2_2|_RX|RB1 _PTL_G2_2|_RX|101 0  2.38752113364072e-12
L_PTL_G2_2|_RX|RB2 _PTL_G2_2|_RX|104 0  1.937922998085e-12
L_PTL_G2_2|_RX|RB3 _PTL_G2_2|_RX|107 0  1.550338398468e-12
B_PTL_G3_2|_TX|1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|2 JJMIT AREA=2.5
B_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|5 JJMIT AREA=2.5
I_PTL_G3_2|_TX|B1 0 _PTL_G3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_2|_TX|B2 0 _PTL_G3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|3  1.684e-12
L_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|6  3.596e-12
L_PTL_G3_2|_TX|1 G3_2 _PTL_G3_2|_TX|1  2.063e-12
L_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|4  4.123e-12
L_PTL_G3_2|_TX|3 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|7  2.193e-12
R_PTL_G3_2|_TX|D _PTL_G3_2|_TX|7 _PTL_G3_2|A_PTL  1.36
L_PTL_G3_2|_TX|P1 _PTL_G3_2|_TX|2 0  5.254e-13
L_PTL_G3_2|_TX|P2 _PTL_G3_2|_TX|5 0  5.141e-13
R_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|101  2.7439617672
R_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|104  2.7439617672
L_PTL_G3_2|_TX|RB1 _PTL_G3_2|_TX|101 0  1.550338398468e-12
L_PTL_G3_2|_TX|RB2 _PTL_G3_2|_TX|104 0  1.550338398468e-12
B_PTL_G3_2|_RX|1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|5 JJMIT AREA=2.0
B_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|8 JJMIT AREA=2.5
I_PTL_G3_2|_RX|B1 0 _PTL_G3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|3  2.777e-12
I_PTL_G3_2|_RX|B2 0 _PTL_G3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|6  2.685e-12
I_PTL_G3_2|_RX|B3 0 _PTL_G3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|9  2.764e-12
L_PTL_G3_2|_RX|1 _PTL_G3_2|A_PTL _PTL_G3_2|_RX|1  1.346e-12
L_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|4  6.348e-12
L_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7  5.197e-12
L_PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7 G3_2_RX  2.058e-12
L_PTL_G3_2|_RX|P1 _PTL_G3_2|_RX|2 0  4.795e-13
L_PTL_G3_2|_RX|P2 _PTL_G3_2|_RX|5 0  5.431e-13
L_PTL_G3_2|_RX|P3 _PTL_G3_2|_RX|8 0  5.339e-13
R_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|101  4.225701121488
R_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|104  3.429952209
R_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|107  2.7439617672
L_PTL_G3_2|_RX|RB1 _PTL_G3_2|_RX|101 0  2.38752113364072e-12
L_PTL_G3_2|_RX|RB2 _PTL_G3_2|_RX|104 0  1.937922998085e-12
L_PTL_G3_2|_RX|RB3 _PTL_G3_2|_RX|107 0  1.550338398468e-12
B_PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_2|_TX|B1 0 _PTL_IP1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_2|_TX|B2 0 _PTL_IP1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|3  1.684e-12
L_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|6  3.596e-12
L_PTL_IP1_2|_TX|1 IP1_2_OUT _PTL_IP1_2|_TX|1  2.063e-12
L_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|4  4.123e-12
L_PTL_IP1_2|_TX|3 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|7  2.193e-12
R_PTL_IP1_2|_TX|D _PTL_IP1_2|_TX|7 _PTL_IP1_2|A_PTL  1.36
L_PTL_IP1_2|_TX|P1 _PTL_IP1_2|_TX|2 0  5.254e-13
L_PTL_IP1_2|_TX|P2 _PTL_IP1_2|_TX|5 0  5.141e-13
R_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|101  2.7439617672
R_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|104  2.7439617672
L_PTL_IP1_2|_TX|RB1 _PTL_IP1_2|_TX|101 0  1.550338398468e-12
L_PTL_IP1_2|_TX|RB2 _PTL_IP1_2|_TX|104 0  1.550338398468e-12
B_PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_2|_RX|B1 0 _PTL_IP1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|3  2.777e-12
I_PTL_IP1_2|_RX|B2 0 _PTL_IP1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|6  2.685e-12
I_PTL_IP1_2|_RX|B3 0 _PTL_IP1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|9  2.764e-12
L_PTL_IP1_2|_RX|1 _PTL_IP1_2|A_PTL _PTL_IP1_2|_RX|1  1.346e-12
L_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|4  6.348e-12
L_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7  5.197e-12
L_PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7 IP1_2_OUT_RX  2.058e-12
L_PTL_IP1_2|_RX|P1 _PTL_IP1_2|_RX|2 0  4.795e-13
L_PTL_IP1_2|_RX|P2 _PTL_IP1_2|_RX|5 0  5.431e-13
L_PTL_IP1_2|_RX|P3 _PTL_IP1_2|_RX|8 0  5.339e-13
R_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|101  4.225701121488
R_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|104  3.429952209
R_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|107  2.7439617672
L_PTL_IP1_2|_RX|RB1 _PTL_IP1_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_2|_RX|RB2 _PTL_IP1_2|_RX|104 0  1.937922998085e-12
L_PTL_IP1_2|_RX|RB3 _PTL_IP1_2|_RX|107 0  1.550338398468e-12
B_PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_2|_TX|B1 0 _PTL_IP2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_2|_TX|B2 0 _PTL_IP2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|3  1.684e-12
L_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|6  3.596e-12
L_PTL_IP2_2|_TX|1 IP2_2_OUT _PTL_IP2_2|_TX|1  2.063e-12
L_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|4  4.123e-12
L_PTL_IP2_2|_TX|3 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|7  2.193e-12
R_PTL_IP2_2|_TX|D _PTL_IP2_2|_TX|7 _PTL_IP2_2|A_PTL  1.36
L_PTL_IP2_2|_TX|P1 _PTL_IP2_2|_TX|2 0  5.254e-13
L_PTL_IP2_2|_TX|P2 _PTL_IP2_2|_TX|5 0  5.141e-13
R_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|101  2.7439617672
R_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|104  2.7439617672
L_PTL_IP2_2|_TX|RB1 _PTL_IP2_2|_TX|101 0  1.550338398468e-12
L_PTL_IP2_2|_TX|RB2 _PTL_IP2_2|_TX|104 0  1.550338398468e-12
B_PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_2|_RX|B1 0 _PTL_IP2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|3  2.777e-12
I_PTL_IP2_2|_RX|B2 0 _PTL_IP2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|6  2.685e-12
I_PTL_IP2_2|_RX|B3 0 _PTL_IP2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|9  2.764e-12
L_PTL_IP2_2|_RX|1 _PTL_IP2_2|A_PTL _PTL_IP2_2|_RX|1  1.346e-12
L_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|4  6.348e-12
L_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7  5.197e-12
L_PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7 IP2_2_OUT_RX  2.058e-12
L_PTL_IP2_2|_RX|P1 _PTL_IP2_2|_RX|2 0  4.795e-13
L_PTL_IP2_2|_RX|P2 _PTL_IP2_2|_RX|5 0  5.431e-13
L_PTL_IP2_2|_RX|P3 _PTL_IP2_2|_RX|8 0  5.339e-13
R_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|101  4.225701121488
R_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|104  3.429952209
R_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|107  2.7439617672
L_PTL_IP2_2|_RX|RB1 _PTL_IP2_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_2|_RX|RB2 _PTL_IP2_2|_RX|104 0  1.937922998085e-12
L_PTL_IP2_2|_RX|RB3 _PTL_IP2_2|_RX|107 0  1.550338398468e-12
B_PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_2|_TX|B1 0 _PTL_IP3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_2|_TX|B2 0 _PTL_IP3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|3  1.684e-12
L_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|6  3.596e-12
L_PTL_IP3_2|_TX|1 IP3_2_OUT _PTL_IP3_2|_TX|1  2.063e-12
L_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|4  4.123e-12
L_PTL_IP3_2|_TX|3 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|7  2.193e-12
R_PTL_IP3_2|_TX|D _PTL_IP3_2|_TX|7 _PTL_IP3_2|A_PTL  1.36
L_PTL_IP3_2|_TX|P1 _PTL_IP3_2|_TX|2 0  5.254e-13
L_PTL_IP3_2|_TX|P2 _PTL_IP3_2|_TX|5 0  5.141e-13
R_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|101  2.7439617672
R_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|104  2.7439617672
L_PTL_IP3_2|_TX|RB1 _PTL_IP3_2|_TX|101 0  1.550338398468e-12
L_PTL_IP3_2|_TX|RB2 _PTL_IP3_2|_TX|104 0  1.550338398468e-12
B_PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_2|_RX|B1 0 _PTL_IP3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|3  2.777e-12
I_PTL_IP3_2|_RX|B2 0 _PTL_IP3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|6  2.685e-12
I_PTL_IP3_2|_RX|B3 0 _PTL_IP3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|9  2.764e-12
L_PTL_IP3_2|_RX|1 _PTL_IP3_2|A_PTL _PTL_IP3_2|_RX|1  1.346e-12
L_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|4  6.348e-12
L_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7  5.197e-12
L_PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7 IP3_2_OUT_RX  2.058e-12
L_PTL_IP3_2|_RX|P1 _PTL_IP3_2|_RX|2 0  4.795e-13
L_PTL_IP3_2|_RX|P2 _PTL_IP3_2|_RX|5 0  5.431e-13
L_PTL_IP3_2|_RX|P3 _PTL_IP3_2|_RX|8 0  5.339e-13
R_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|101  4.225701121488
R_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|104  3.429952209
R_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|107  2.7439617672
L_PTL_IP3_2|_RX|RB1 _PTL_IP3_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_2|_RX|RB2 _PTL_IP3_2|_RX|104 0  1.937922998085e-12
L_PTL_IP3_2|_RX|RB3 _PTL_IP3_2|_RX|107 0  1.550338398468e-12
LI0|_AND|I_A1|B I0|_AND|A1 I0|_AND|I_A1|MID  2e-12
II0|_AND|I_A1|B 0 I0|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_B1|B I0|_AND|B1 I0|_AND|I_B1|MID  2e-12
II0|_AND|I_B1|B 0 I0|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q3|B I0|_AND|Q3 I0|_AND|I_Q3|MID  2e-12
II0|_AND|I_Q3|B 0 I0|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0|_AND|I_Q2|B I0|_AND|Q2 I0|_AND|I_Q2|MID  2e-12
II0|_AND|I_Q2|B 0 I0|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q1|B I0|_AND|Q1 I0|_AND|I_Q1|MID  2e-12
II0|_AND|I_Q1|B 0 I0|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_AND|A1|1 I0|_AND|A1 I0|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A1|P I0|_AND|A1|MID_SERIES 0  2e-13
RI0|_AND|A1|B I0|_AND|A1 I0|_AND|A1|MID_SHUNT  2.7439617672
LI0|_AND|A1|RB I0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A2|1 I0|_AND|A2 I0|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A2|P I0|_AND|A2|MID_SERIES 0  2e-13
RI0|_AND|A2|B I0|_AND|A2 I0|_AND|A2|MID_SHUNT  2.7439617672
LI0|_AND|A2|RB I0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A12|1 I0|_AND|A2 I0|_AND|A3 JJMIT AREA=1.7857142857142858
RI0|_AND|A12|B I0|_AND|A2 I0|_AND|A12|MID_SHUNT  3.84154647408
LI0|_AND|A12|RB I0|_AND|A12|MID_SHUNT I0|_AND|A3  2.1704737578552e-12
BI0|_AND|B1|1 I0|_AND|B1 I0|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B1|P I0|_AND|B1|MID_SERIES 0  2e-13
RI0|_AND|B1|B I0|_AND|B1 I0|_AND|B1|MID_SHUNT  2.7439617672
LI0|_AND|B1|RB I0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B2|1 I0|_AND|B2 I0|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B2|P I0|_AND|B2|MID_SERIES 0  2e-13
RI0|_AND|B2|B I0|_AND|B2 I0|_AND|B2|MID_SHUNT  2.7439617672
LI0|_AND|B2|RB I0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B12|1 I0|_AND|B2 I0|_AND|B3 JJMIT AREA=1.7857142857142858
RI0|_AND|B12|B I0|_AND|B2 I0|_AND|B12|MID_SHUNT  3.84154647408
LI0|_AND|B12|RB I0|_AND|B12|MID_SHUNT I0|_AND|B3  2.1704737578552e-12
BI0|_AND|Q2|1 I0|_AND|Q2 I0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q2|P I0|_AND|Q2|MID_SERIES 0  2e-13
RI0|_AND|Q2|B I0|_AND|Q2 I0|_AND|Q2|MID_SHUNT  2.7439617672
LI0|_AND|Q2|RB I0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|Q1|1 I0|_AND|Q1 I0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q1|P I0|_AND|Q1|MID_SERIES 0  2e-13
RI0|_AND|Q1|B I0|_AND|Q1 I0|_AND|Q1|MID_SHUNT  2.7439617672
LI0|_AND|Q1|RB I0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1|_AND|I_A1|B I1|_AND|A1 I1|_AND|I_A1|MID  2e-12
II1|_AND|I_A1|B 0 I1|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_B1|B I1|_AND|B1 I1|_AND|I_B1|MID  2e-12
II1|_AND|I_B1|B 0 I1|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q3|B I1|_AND|Q3 I1|_AND|I_Q3|MID  2e-12
II1|_AND|I_Q3|B 0 I1|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1|_AND|I_Q2|B I1|_AND|Q2 I1|_AND|I_Q2|MID  2e-12
II1|_AND|I_Q2|B 0 I1|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q1|B I1|_AND|Q1 I1|_AND|I_Q1|MID  2e-12
II1|_AND|I_Q1|B 0 I1|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_AND|A1|1 I1|_AND|A1 I1|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A1|P I1|_AND|A1|MID_SERIES 0  2e-13
RI1|_AND|A1|B I1|_AND|A1 I1|_AND|A1|MID_SHUNT  2.7439617672
LI1|_AND|A1|RB I1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A2|1 I1|_AND|A2 I1|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A2|P I1|_AND|A2|MID_SERIES 0  2e-13
RI1|_AND|A2|B I1|_AND|A2 I1|_AND|A2|MID_SHUNT  2.7439617672
LI1|_AND|A2|RB I1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A12|1 I1|_AND|A2 I1|_AND|A3 JJMIT AREA=1.7857142857142858
RI1|_AND|A12|B I1|_AND|A2 I1|_AND|A12|MID_SHUNT  3.84154647408
LI1|_AND|A12|RB I1|_AND|A12|MID_SHUNT I1|_AND|A3  2.1704737578552e-12
BI1|_AND|B1|1 I1|_AND|B1 I1|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B1|P I1|_AND|B1|MID_SERIES 0  2e-13
RI1|_AND|B1|B I1|_AND|B1 I1|_AND|B1|MID_SHUNT  2.7439617672
LI1|_AND|B1|RB I1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B2|1 I1|_AND|B2 I1|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B2|P I1|_AND|B2|MID_SERIES 0  2e-13
RI1|_AND|B2|B I1|_AND|B2 I1|_AND|B2|MID_SHUNT  2.7439617672
LI1|_AND|B2|RB I1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B12|1 I1|_AND|B2 I1|_AND|B3 JJMIT AREA=1.7857142857142858
RI1|_AND|B12|B I1|_AND|B2 I1|_AND|B12|MID_SHUNT  3.84154647408
LI1|_AND|B12|RB I1|_AND|B12|MID_SHUNT I1|_AND|B3  2.1704737578552e-12
BI1|_AND|Q2|1 I1|_AND|Q2 I1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q2|P I1|_AND|Q2|MID_SERIES 0  2e-13
RI1|_AND|Q2|B I1|_AND|Q2 I1|_AND|Q2|MID_SHUNT  2.7439617672
LI1|_AND|Q2|RB I1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|Q1|1 I1|_AND|Q1 I1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q1|P I1|_AND|Q1|MID_SERIES 0  2e-13
RI1|_AND|Q1|B I1|_AND|Q1 I1|_AND|Q1|MID_SHUNT  2.7439617672
LI1|_AND|Q1|RB I1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2|_AND|I_A1|B I2|_AND|A1 I2|_AND|I_A1|MID  2e-12
II2|_AND|I_A1|B 0 I2|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_B1|B I2|_AND|B1 I2|_AND|I_B1|MID  2e-12
II2|_AND|I_B1|B 0 I2|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q3|B I2|_AND|Q3 I2|_AND|I_Q3|MID  2e-12
II2|_AND|I_Q3|B 0 I2|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2|_AND|I_Q2|B I2|_AND|Q2 I2|_AND|I_Q2|MID  2e-12
II2|_AND|I_Q2|B 0 I2|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q1|B I2|_AND|Q1 I2|_AND|I_Q1|MID  2e-12
II2|_AND|I_Q1|B 0 I2|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_AND|A1|1 I2|_AND|A1 I2|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A1|P I2|_AND|A1|MID_SERIES 0  2e-13
RI2|_AND|A1|B I2|_AND|A1 I2|_AND|A1|MID_SHUNT  2.7439617672
LI2|_AND|A1|RB I2|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A2|1 I2|_AND|A2 I2|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A2|P I2|_AND|A2|MID_SERIES 0  2e-13
RI2|_AND|A2|B I2|_AND|A2 I2|_AND|A2|MID_SHUNT  2.7439617672
LI2|_AND|A2|RB I2|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A12|1 I2|_AND|A2 I2|_AND|A3 JJMIT AREA=1.7857142857142858
RI2|_AND|A12|B I2|_AND|A2 I2|_AND|A12|MID_SHUNT  3.84154647408
LI2|_AND|A12|RB I2|_AND|A12|MID_SHUNT I2|_AND|A3  2.1704737578552e-12
BI2|_AND|B1|1 I2|_AND|B1 I2|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B1|P I2|_AND|B1|MID_SERIES 0  2e-13
RI2|_AND|B1|B I2|_AND|B1 I2|_AND|B1|MID_SHUNT  2.7439617672
LI2|_AND|B1|RB I2|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B2|1 I2|_AND|B2 I2|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B2|P I2|_AND|B2|MID_SERIES 0  2e-13
RI2|_AND|B2|B I2|_AND|B2 I2|_AND|B2|MID_SHUNT  2.7439617672
LI2|_AND|B2|RB I2|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B12|1 I2|_AND|B2 I2|_AND|B3 JJMIT AREA=1.7857142857142858
RI2|_AND|B12|B I2|_AND|B2 I2|_AND|B12|MID_SHUNT  3.84154647408
LI2|_AND|B12|RB I2|_AND|B12|MID_SHUNT I2|_AND|B3  2.1704737578552e-12
BI2|_AND|Q2|1 I2|_AND|Q2 I2|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q2|P I2|_AND|Q2|MID_SERIES 0  2e-13
RI2|_AND|Q2|B I2|_AND|Q2 I2|_AND|Q2|MID_SHUNT  2.7439617672
LI2|_AND|Q2|RB I2|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|Q1|1 I2|_AND|Q1 I2|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q1|P I2|_AND|Q1|MID_SERIES 0  2e-13
RI2|_AND|Q1|B I2|_AND|Q1 I2|_AND|Q1|MID_SHUNT  2.7439617672
LI2|_AND|Q1|RB I2|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3|_AND|I_A1|B I3|_AND|A1 I3|_AND|I_A1|MID  2e-12
II3|_AND|I_A1|B 0 I3|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_B1|B I3|_AND|B1 I3|_AND|I_B1|MID  2e-12
II3|_AND|I_B1|B 0 I3|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q3|B I3|_AND|Q3 I3|_AND|I_Q3|MID  2e-12
II3|_AND|I_Q3|B 0 I3|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3|_AND|I_Q2|B I3|_AND|Q2 I3|_AND|I_Q2|MID  2e-12
II3|_AND|I_Q2|B 0 I3|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q1|B I3|_AND|Q1 I3|_AND|I_Q1|MID  2e-12
II3|_AND|I_Q1|B 0 I3|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_AND|A1|1 I3|_AND|A1 I3|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A1|P I3|_AND|A1|MID_SERIES 0  2e-13
RI3|_AND|A1|B I3|_AND|A1 I3|_AND|A1|MID_SHUNT  2.7439617672
LI3|_AND|A1|RB I3|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A2|1 I3|_AND|A2 I3|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A2|P I3|_AND|A2|MID_SERIES 0  2e-13
RI3|_AND|A2|B I3|_AND|A2 I3|_AND|A2|MID_SHUNT  2.7439617672
LI3|_AND|A2|RB I3|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A12|1 I3|_AND|A2 I3|_AND|A3 JJMIT AREA=1.7857142857142858
RI3|_AND|A12|B I3|_AND|A2 I3|_AND|A12|MID_SHUNT  3.84154647408
LI3|_AND|A12|RB I3|_AND|A12|MID_SHUNT I3|_AND|A3  2.1704737578552e-12
BI3|_AND|B1|1 I3|_AND|B1 I3|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B1|P I3|_AND|B1|MID_SERIES 0  2e-13
RI3|_AND|B1|B I3|_AND|B1 I3|_AND|B1|MID_SHUNT  2.7439617672
LI3|_AND|B1|RB I3|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B2|1 I3|_AND|B2 I3|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B2|P I3|_AND|B2|MID_SERIES 0  2e-13
RI3|_AND|B2|B I3|_AND|B2 I3|_AND|B2|MID_SHUNT  2.7439617672
LI3|_AND|B2|RB I3|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B12|1 I3|_AND|B2 I3|_AND|B3 JJMIT AREA=1.7857142857142858
RI3|_AND|B12|B I3|_AND|B2 I3|_AND|B12|MID_SHUNT  3.84154647408
LI3|_AND|B12|RB I3|_AND|B12|MID_SHUNT I3|_AND|B3  2.1704737578552e-12
BI3|_AND|Q2|1 I3|_AND|Q2 I3|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q2|P I3|_AND|Q2|MID_SERIES 0  2e-13
RI3|_AND|Q2|B I3|_AND|Q2 I3|_AND|Q2|MID_SHUNT  2.7439617672
LI3|_AND|Q2|RB I3|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|Q1|1 I3|_AND|Q1 I3|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q1|P I3|_AND|Q1|MID_SERIES 0  2e-13
RI3|_AND|Q1|B I3|_AND|Q1 I3|_AND|Q1|MID_SHUNT  2.7439617672
LI3|_AND|Q1|RB I3|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|I_D1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|I_D1|MID  2e-12
ISPL_IP2_0|SPL1|I_D1|B 0 SPL_IP2_0|SPL1|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0|SPL1|I_D2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|I_D2|MID  2e-12
ISPL_IP2_0|SPL1|I_D2|B 0 SPL_IP2_0|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IP2_0|SPL1|I_Q1|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|I_Q1|MID  2e-12
ISPL_IP2_0|SPL1|I_Q1|B 0 SPL_IP2_0|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0|SPL1|I_Q2|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|I_Q2|MID  2e-12
ISPL_IP2_0|SPL1|I_Q2|B 0 SPL_IP2_0|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IP2_0|SPL1|1|1 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|1|P SPL_IP2_0|SPL1|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|1|RB SPL_IP2_0|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|2|1 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|2|P SPL_IP2_0|SPL1|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|2|RB SPL_IP2_0|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|A|1 SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|A|P SPL_IP2_0|SPL1|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|A|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|A|RB SPL_IP2_0|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|B|1 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|B|P SPL_IP2_0|SPL1|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|B|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|B|RB SPL_IP2_0|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL2|I_D1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|I_D1|MID  2e-12
ISPL_IP2_0|SPL2|I_D1|B 0 SPL_IP2_0|SPL2|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0|SPL2|I_D2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|I_D2|MID  2e-12
ISPL_IP2_0|SPL2|I_D2|B 0 SPL_IP2_0|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IP2_0|SPL2|I_Q1|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|I_Q1|MID  2e-12
ISPL_IP2_0|SPL2|I_Q1|B 0 SPL_IP2_0|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0|SPL2|I_Q2|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|I_Q2|MID  2e-12
ISPL_IP2_0|SPL2|I_Q2|B 0 SPL_IP2_0|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IP2_0|SPL2|1|1 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|1|P SPL_IP2_0|SPL2|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|1|RB SPL_IP2_0|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|2|1 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|2|P SPL_IP2_0|SPL2|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|2|RB SPL_IP2_0|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|A|1 SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|A|P SPL_IP2_0|SPL2|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|A|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|A|RB SPL_IP2_0|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|B|1 SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|B|P SPL_IP2_0|SPL2|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|B|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|B|RB SPL_IP2_0|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_PG|I_A1|B _PG1_01|_PG|A1 _PG1_01|_PG|I_A1|MID  2e-12
I_PG1_01|_PG|I_A1|B 0 _PG1_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_B1|B _PG1_01|_PG|B1 _PG1_01|_PG|I_B1|MID  2e-12
I_PG1_01|_PG|I_B1|B 0 _PG1_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q3|B _PG1_01|_PG|Q3 _PG1_01|_PG|I_Q3|MID  2e-12
I_PG1_01|_PG|I_Q3|B 0 _PG1_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_PG|I_Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|I_Q2|MID  2e-12
I_PG1_01|_PG|I_Q2|B 0 _PG1_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|I_Q1|MID  2e-12
I_PG1_01|_PG|I_Q1|B 0 _PG1_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_PG|A1|1 _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A1|P _PG1_01|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01|_PG|A1|B _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A1|RB _PG1_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A2|1 _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A2|P _PG1_01|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01|_PG|A2|B _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A2|RB _PG1_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A12|1 _PG1_01|_PG|A2 _PG1_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|A12|B _PG1_01|_PG|A2 _PG1_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|A12|RB _PG1_01|_PG|A12|MID_SHUNT _PG1_01|_PG|A3  2.1704737578552e-12
B_PG1_01|_PG|B1|1 _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B1|P _PG1_01|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01|_PG|B1|B _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B1|RB _PG1_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B2|1 _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B2|P _PG1_01|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01|_PG|B2|B _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B2|RB _PG1_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B12|1 _PG1_01|_PG|B2 _PG1_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|B12|B _PG1_01|_PG|B2 _PG1_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|B12|RB _PG1_01|_PG|B12|MID_SHUNT _PG1_01|_PG|B3  2.1704737578552e-12
B_PG1_01|_PG|Q2|1 _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q2|P _PG1_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q2|RB _PG1_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|Q1|1 _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q1|P _PG1_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q1|RB _PG1_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_GG|I_A1|B _PG1_01|_GG|A1 _PG1_01|_GG|I_A1|MID  2e-12
I_PG1_01|_GG|I_A1|B 0 _PG1_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_B1|B _PG1_01|_GG|B1 _PG1_01|_GG|I_B1|MID  2e-12
I_PG1_01|_GG|I_B1|B 0 _PG1_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q3|B _PG1_01|_GG|Q3 _PG1_01|_GG|I_Q3|MID  2e-12
I_PG1_01|_GG|I_Q3|B 0 _PG1_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_GG|I_Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|I_Q2|MID  2e-12
I_PG1_01|_GG|I_Q2|B 0 _PG1_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|I_Q1|MID  2e-12
I_PG1_01|_GG|I_Q1|B 0 _PG1_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_GG|A1|1 _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A1|P _PG1_01|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01|_GG|A1|B _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A1|RB _PG1_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A2|1 _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A2|P _PG1_01|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01|_GG|A2|B _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A2|RB _PG1_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A12|1 _PG1_01|_GG|A2 _PG1_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|A12|B _PG1_01|_GG|A2 _PG1_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|A12|RB _PG1_01|_GG|A12|MID_SHUNT _PG1_01|_GG|A3  2.1704737578552e-12
B_PG1_01|_GG|B1|1 _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B1|P _PG1_01|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01|_GG|B1|B _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B1|RB _PG1_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B2|1 _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B2|P _PG1_01|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01|_GG|B2|B _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B2|RB _PG1_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B12|1 _PG1_01|_GG|B2 _PG1_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|B12|B _PG1_01|_GG|B2 _PG1_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|B12|RB _PG1_01|_GG|B12|MID_SHUNT _PG1_01|_GG|B3  2.1704737578552e-12
B_PG1_01|_GG|Q2|1 _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q2|P _PG1_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q2|RB _PG1_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|Q1|1 _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q1|P _PG1_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q1|RB _PG1_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_G|I_A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|I_A1|MID  2e-12
I_PG1_01|_AND_G|I_A1|B 0 _PG1_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|I_B1|MID  2e-12
I_PG1_01|_AND_G|I_B1|B 0 _PG1_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q3|B _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|I_Q3|MID  2e-12
I_PG1_01|_AND_G|I_Q3|B 0 _PG1_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_G|I_Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|I_Q2|MID  2e-12
I_PG1_01|_AND_G|I_Q2|B 0 _PG1_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|I_Q1|MID  2e-12
I_PG1_01|_AND_G|I_Q1|B 0 _PG1_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_G|A1|1 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A1|P _PG1_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A1|RB _PG1_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A2|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A2|P _PG1_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A2|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A2|RB _PG1_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A12|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|A12|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|A12|RB _PG1_01|_AND_G|A12|MID_SHUNT _PG1_01|_AND_G|A3  2.1704737578552e-12
B_PG1_01|_AND_G|B1|1 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B1|P _PG1_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B1|RB _PG1_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B2|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B2|P _PG1_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B2|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B2|RB _PG1_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B12|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|B12|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|B12|RB _PG1_01|_AND_G|B12|MID_SHUNT _PG1_01|_AND_G|B3  2.1704737578552e-12
B_PG1_01|_AND_G|Q2|1 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q2|P _PG1_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q2|RB _PG1_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|Q1|1 _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q1|P _PG1_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q1|RB _PG1_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_PG|I_A1|B _PG3_01|_PG|A1 _PG3_01|_PG|I_A1|MID  2e-12
I_PG3_01|_PG|I_A1|B 0 _PG3_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_B1|B _PG3_01|_PG|B1 _PG3_01|_PG|I_B1|MID  2e-12
I_PG3_01|_PG|I_B1|B 0 _PG3_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q3|B _PG3_01|_PG|Q3 _PG3_01|_PG|I_Q3|MID  2e-12
I_PG3_01|_PG|I_Q3|B 0 _PG3_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_PG|I_Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|I_Q2|MID  2e-12
I_PG3_01|_PG|I_Q2|B 0 _PG3_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|I_Q1|MID  2e-12
I_PG3_01|_PG|I_Q1|B 0 _PG3_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_PG|A1|1 _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A1|P _PG3_01|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01|_PG|A1|B _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A1|RB _PG3_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A2|1 _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A2|P _PG3_01|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01|_PG|A2|B _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A2|RB _PG3_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A12|1 _PG3_01|_PG|A2 _PG3_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|A12|B _PG3_01|_PG|A2 _PG3_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|A12|RB _PG3_01|_PG|A12|MID_SHUNT _PG3_01|_PG|A3  2.1704737578552e-12
B_PG3_01|_PG|B1|1 _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B1|P _PG3_01|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01|_PG|B1|B _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B1|RB _PG3_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B2|1 _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B2|P _PG3_01|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01|_PG|B2|B _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B2|RB _PG3_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B12|1 _PG3_01|_PG|B2 _PG3_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|B12|B _PG3_01|_PG|B2 _PG3_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|B12|RB _PG3_01|_PG|B12|MID_SHUNT _PG3_01|_PG|B3  2.1704737578552e-12
B_PG3_01|_PG|Q2|1 _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q2|P _PG3_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q2|RB _PG3_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|Q1|1 _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q1|P _PG3_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q1|RB _PG3_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_GG|I_A1|B _PG3_01|_GG|A1 _PG3_01|_GG|I_A1|MID  2e-12
I_PG3_01|_GG|I_A1|B 0 _PG3_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_B1|B _PG3_01|_GG|B1 _PG3_01|_GG|I_B1|MID  2e-12
I_PG3_01|_GG|I_B1|B 0 _PG3_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q3|B _PG3_01|_GG|Q3 _PG3_01|_GG|I_Q3|MID  2e-12
I_PG3_01|_GG|I_Q3|B 0 _PG3_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_GG|I_Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|I_Q2|MID  2e-12
I_PG3_01|_GG|I_Q2|B 0 _PG3_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|I_Q1|MID  2e-12
I_PG3_01|_GG|I_Q1|B 0 _PG3_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_GG|A1|1 _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A1|P _PG3_01|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01|_GG|A1|B _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A1|RB _PG3_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A2|1 _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A2|P _PG3_01|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01|_GG|A2|B _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A2|RB _PG3_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A12|1 _PG3_01|_GG|A2 _PG3_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|A12|B _PG3_01|_GG|A2 _PG3_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|A12|RB _PG3_01|_GG|A12|MID_SHUNT _PG3_01|_GG|A3  2.1704737578552e-12
B_PG3_01|_GG|B1|1 _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B1|P _PG3_01|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01|_GG|B1|B _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B1|RB _PG3_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B2|1 _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B2|P _PG3_01|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01|_GG|B2|B _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B2|RB _PG3_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B12|1 _PG3_01|_GG|B2 _PG3_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|B12|B _PG3_01|_GG|B2 _PG3_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|B12|RB _PG3_01|_GG|B12|MID_SHUNT _PG3_01|_GG|B3  2.1704737578552e-12
B_PG3_01|_GG|Q2|1 _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q2|P _PG3_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q2|RB _PG3_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|Q1|1 _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q1|P _PG3_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q1|RB _PG3_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_G|I_A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|I_A1|MID  2e-12
I_PG3_01|_AND_G|I_A1|B 0 _PG3_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|I_B1|MID  2e-12
I_PG3_01|_AND_G|I_B1|B 0 _PG3_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q3|B _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|I_Q3|MID  2e-12
I_PG3_01|_AND_G|I_Q3|B 0 _PG3_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_G|I_Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|I_Q2|MID  2e-12
I_PG3_01|_AND_G|I_Q2|B 0 _PG3_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|I_Q1|MID  2e-12
I_PG3_01|_AND_G|I_Q1|B 0 _PG3_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_G|A1|1 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A1|P _PG3_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A1|RB _PG3_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A2|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A2|P _PG3_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A2|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A2|RB _PG3_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A12|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|A12|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|A12|RB _PG3_01|_AND_G|A12|MID_SHUNT _PG3_01|_AND_G|A3  2.1704737578552e-12
B_PG3_01|_AND_G|B1|1 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B1|P _PG3_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B1|RB _PG3_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B2|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B2|P _PG3_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B2|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B2|RB _PG3_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B12|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|B12|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|B12|RB _PG3_01|_AND_G|B12|MID_SHUNT _PG3_01|_AND_G|B3  2.1704737578552e-12
B_PG3_01|_AND_G|Q2|1 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q2|P _PG3_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q2|RB _PG3_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|Q1|1 _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q1|P _PG3_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q1|RB _PG3_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_P|I_A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|I_A1|MID  2e-12
I_PG3_01|_AND_P|I_A1|B 0 _PG3_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|I_B1|MID  2e-12
I_PG3_01|_AND_P|I_B1|B 0 _PG3_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q3|B _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|I_Q3|MID  2e-12
I_PG3_01|_AND_P|I_Q3|B 0 _PG3_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_P|I_Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|I_Q2|MID  2e-12
I_PG3_01|_AND_P|I_Q2|B 0 _PG3_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|I_Q1|MID  2e-12
I_PG3_01|_AND_P|I_Q1|B 0 _PG3_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_P|A1|1 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A1|P _PG3_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A1|RB _PG3_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A2|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A2|P _PG3_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A2|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A2|RB _PG3_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A12|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|A12|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|A12|RB _PG3_01|_AND_P|A12|MID_SHUNT _PG3_01|_AND_P|A3  2.1704737578552e-12
B_PG3_01|_AND_P|B1|1 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B1|P _PG3_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B1|RB _PG3_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B2|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B2|P _PG3_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B2|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B2|RB _PG3_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B12|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|B12|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|B12|RB _PG3_01|_AND_P|B12|MID_SHUNT _PG3_01|_AND_P|B3  2.1704737578552e-12
B_PG3_01|_AND_P|Q2|1 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q2|P _PG3_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q2|RB _PG3_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|Q1|1 _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q1|P _PG3_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q1|RB _PG3_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL1|I_D1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|I_D1|MID  2e-12
ISPL_G1_1|SPL1|I_D1|B 0 SPL_G1_1|SPL1|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1|SPL1|I_D2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|I_D2|MID  2e-12
ISPL_G1_1|SPL1|I_D2|B 0 SPL_G1_1|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_G1_1|SPL1|I_Q1|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|I_Q1|MID  2e-12
ISPL_G1_1|SPL1|I_Q1|B 0 SPL_G1_1|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1|SPL1|I_Q2|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|I_Q2|MID  2e-12
ISPL_G1_1|SPL1|I_Q2|B 0 SPL_G1_1|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_G1_1|SPL1|1|1 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|1|P SPL_G1_1|SPL1|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|1|RB SPL_G1_1|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|2|1 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|2|P SPL_G1_1|SPL1|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|2|RB SPL_G1_1|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|A|1 SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|A|P SPL_G1_1|SPL1|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|A|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|A|RB SPL_G1_1|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|B|1 SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|B|P SPL_G1_1|SPL1|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|B|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|B|RB SPL_G1_1|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL2|I_D1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|I_D1|MID  2e-12
ISPL_G1_1|SPL2|I_D1|B 0 SPL_G1_1|SPL2|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1|SPL2|I_D2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|I_D2|MID  2e-12
ISPL_G1_1|SPL2|I_D2|B 0 SPL_G1_1|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_G1_1|SPL2|I_Q1|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|I_Q1|MID  2e-12
ISPL_G1_1|SPL2|I_Q1|B 0 SPL_G1_1|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1|SPL2|I_Q2|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|I_Q2|MID  2e-12
ISPL_G1_1|SPL2|I_Q2|B 0 SPL_G1_1|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_G1_1|SPL2|1|1 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|1|P SPL_G1_1|SPL2|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|1|RB SPL_G1_1|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|2|1 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|2|P SPL_G1_1|SPL2|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|2|RB SPL_G1_1|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|A|1 SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|A|P SPL_G1_1|SPL2|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|A|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|A|RB SPL_G1_1|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|B|1 SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|B|P SPL_G1_1|SPL2|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|B|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|B|RB SPL_G1_1|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_PG|I_A1|B _PG2_12|_PG|A1 _PG2_12|_PG|I_A1|MID  2e-12
I_PG2_12|_PG|I_A1|B 0 _PG2_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_B1|B _PG2_12|_PG|B1 _PG2_12|_PG|I_B1|MID  2e-12
I_PG2_12|_PG|I_B1|B 0 _PG2_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q3|B _PG2_12|_PG|Q3 _PG2_12|_PG|I_Q3|MID  2e-12
I_PG2_12|_PG|I_Q3|B 0 _PG2_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_PG|I_Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|I_Q2|MID  2e-12
I_PG2_12|_PG|I_Q2|B 0 _PG2_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|I_Q1|MID  2e-12
I_PG2_12|_PG|I_Q1|B 0 _PG2_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_PG|A1|1 _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A1|P _PG2_12|_PG|A1|MID_SERIES 0  2e-13
R_PG2_12|_PG|A1|B _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A1|RB _PG2_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A2|1 _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A2|P _PG2_12|_PG|A2|MID_SERIES 0  2e-13
R_PG2_12|_PG|A2|B _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A2|RB _PG2_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A12|1 _PG2_12|_PG|A2 _PG2_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|A12|B _PG2_12|_PG|A2 _PG2_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|A12|RB _PG2_12|_PG|A12|MID_SHUNT _PG2_12|_PG|A3  2.1704737578552e-12
B_PG2_12|_PG|B1|1 _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B1|P _PG2_12|_PG|B1|MID_SERIES 0  2e-13
R_PG2_12|_PG|B1|B _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B1|RB _PG2_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B2|1 _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B2|P _PG2_12|_PG|B2|MID_SERIES 0  2e-13
R_PG2_12|_PG|B2|B _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B2|RB _PG2_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B12|1 _PG2_12|_PG|B2 _PG2_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|B12|B _PG2_12|_PG|B2 _PG2_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|B12|RB _PG2_12|_PG|B12|MID_SHUNT _PG2_12|_PG|B3  2.1704737578552e-12
B_PG2_12|_PG|Q2|1 _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q2|P _PG2_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q2|RB _PG2_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|Q1|1 _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q1|P _PG2_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q1|RB _PG2_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_GG|I_A1|B _PG2_12|_GG|A1 _PG2_12|_GG|I_A1|MID  2e-12
I_PG2_12|_GG|I_A1|B 0 _PG2_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_B1|B _PG2_12|_GG|B1 _PG2_12|_GG|I_B1|MID  2e-12
I_PG2_12|_GG|I_B1|B 0 _PG2_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q3|B _PG2_12|_GG|Q3 _PG2_12|_GG|I_Q3|MID  2e-12
I_PG2_12|_GG|I_Q3|B 0 _PG2_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_GG|I_Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|I_Q2|MID  2e-12
I_PG2_12|_GG|I_Q2|B 0 _PG2_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|I_Q1|MID  2e-12
I_PG2_12|_GG|I_Q1|B 0 _PG2_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_GG|A1|1 _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A1|P _PG2_12|_GG|A1|MID_SERIES 0  2e-13
R_PG2_12|_GG|A1|B _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A1|RB _PG2_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A2|1 _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A2|P _PG2_12|_GG|A2|MID_SERIES 0  2e-13
R_PG2_12|_GG|A2|B _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A2|RB _PG2_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A12|1 _PG2_12|_GG|A2 _PG2_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|A12|B _PG2_12|_GG|A2 _PG2_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|A12|RB _PG2_12|_GG|A12|MID_SHUNT _PG2_12|_GG|A3  2.1704737578552e-12
B_PG2_12|_GG|B1|1 _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B1|P _PG2_12|_GG|B1|MID_SERIES 0  2e-13
R_PG2_12|_GG|B1|B _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B1|RB _PG2_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B2|1 _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B2|P _PG2_12|_GG|B2|MID_SERIES 0  2e-13
R_PG2_12|_GG|B2|B _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B2|RB _PG2_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B12|1 _PG2_12|_GG|B2 _PG2_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|B12|B _PG2_12|_GG|B2 _PG2_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|B12|RB _PG2_12|_GG|B12|MID_SHUNT _PG2_12|_GG|B3  2.1704737578552e-12
B_PG2_12|_GG|Q2|1 _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q2|P _PG2_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q2|RB _PG2_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|Q1|1 _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q1|P _PG2_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q1|RB _PG2_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_G|I_A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|I_A1|MID  2e-12
I_PG2_12|_AND_G|I_A1|B 0 _PG2_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|I_B1|MID  2e-12
I_PG2_12|_AND_G|I_B1|B 0 _PG2_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q3|B _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|I_Q3|MID  2e-12
I_PG2_12|_AND_G|I_Q3|B 0 _PG2_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_G|I_Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|I_Q2|MID  2e-12
I_PG2_12|_AND_G|I_Q2|B 0 _PG2_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|I_Q1|MID  2e-12
I_PG2_12|_AND_G|I_Q1|B 0 _PG2_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_G|A1|1 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A1|P _PG2_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A1|RB _PG2_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A2|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A2|P _PG2_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A2|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A2|RB _PG2_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A12|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|A12|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|A12|RB _PG2_12|_AND_G|A12|MID_SHUNT _PG2_12|_AND_G|A3  2.1704737578552e-12
B_PG2_12|_AND_G|B1|1 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B1|P _PG2_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B1|RB _PG2_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B2|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B2|P _PG2_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B2|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B2|RB _PG2_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B12|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|B12|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|B12|RB _PG2_12|_AND_G|B12|MID_SHUNT _PG2_12|_AND_G|B3  2.1704737578552e-12
B_PG2_12|_AND_G|Q2|1 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q2|P _PG2_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q2|RB _PG2_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|Q1|1 _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q1|P _PG2_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q1|RB _PG2_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_PG|I_A1|B _PG3_12|_PG|A1 _PG3_12|_PG|I_A1|MID  2e-12
I_PG3_12|_PG|I_A1|B 0 _PG3_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_B1|B _PG3_12|_PG|B1 _PG3_12|_PG|I_B1|MID  2e-12
I_PG3_12|_PG|I_B1|B 0 _PG3_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q3|B _PG3_12|_PG|Q3 _PG3_12|_PG|I_Q3|MID  2e-12
I_PG3_12|_PG|I_Q3|B 0 _PG3_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_PG|I_Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|I_Q2|MID  2e-12
I_PG3_12|_PG|I_Q2|B 0 _PG3_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|I_Q1|MID  2e-12
I_PG3_12|_PG|I_Q1|B 0 _PG3_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_PG|A1|1 _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A1|P _PG3_12|_PG|A1|MID_SERIES 0  2e-13
R_PG3_12|_PG|A1|B _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A1|RB _PG3_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A2|1 _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A2|P _PG3_12|_PG|A2|MID_SERIES 0  2e-13
R_PG3_12|_PG|A2|B _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A2|RB _PG3_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A12|1 _PG3_12|_PG|A2 _PG3_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|A12|B _PG3_12|_PG|A2 _PG3_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|A12|RB _PG3_12|_PG|A12|MID_SHUNT _PG3_12|_PG|A3  2.1704737578552e-12
B_PG3_12|_PG|B1|1 _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B1|P _PG3_12|_PG|B1|MID_SERIES 0  2e-13
R_PG3_12|_PG|B1|B _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B1|RB _PG3_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B2|1 _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B2|P _PG3_12|_PG|B2|MID_SERIES 0  2e-13
R_PG3_12|_PG|B2|B _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B2|RB _PG3_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B12|1 _PG3_12|_PG|B2 _PG3_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|B12|B _PG3_12|_PG|B2 _PG3_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|B12|RB _PG3_12|_PG|B12|MID_SHUNT _PG3_12|_PG|B3  2.1704737578552e-12
B_PG3_12|_PG|Q2|1 _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q2|P _PG3_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q2|RB _PG3_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|Q1|1 _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q1|P _PG3_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q1|RB _PG3_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_GG|I_A1|B _PG3_12|_GG|A1 _PG3_12|_GG|I_A1|MID  2e-12
I_PG3_12|_GG|I_A1|B 0 _PG3_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_B1|B _PG3_12|_GG|B1 _PG3_12|_GG|I_B1|MID  2e-12
I_PG3_12|_GG|I_B1|B 0 _PG3_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q3|B _PG3_12|_GG|Q3 _PG3_12|_GG|I_Q3|MID  2e-12
I_PG3_12|_GG|I_Q3|B 0 _PG3_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_GG|I_Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|I_Q2|MID  2e-12
I_PG3_12|_GG|I_Q2|B 0 _PG3_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|I_Q1|MID  2e-12
I_PG3_12|_GG|I_Q1|B 0 _PG3_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_GG|A1|1 _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A1|P _PG3_12|_GG|A1|MID_SERIES 0  2e-13
R_PG3_12|_GG|A1|B _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A1|RB _PG3_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A2|1 _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A2|P _PG3_12|_GG|A2|MID_SERIES 0  2e-13
R_PG3_12|_GG|A2|B _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A2|RB _PG3_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A12|1 _PG3_12|_GG|A2 _PG3_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|A12|B _PG3_12|_GG|A2 _PG3_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|A12|RB _PG3_12|_GG|A12|MID_SHUNT _PG3_12|_GG|A3  2.1704737578552e-12
B_PG3_12|_GG|B1|1 _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B1|P _PG3_12|_GG|B1|MID_SERIES 0  2e-13
R_PG3_12|_GG|B1|B _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B1|RB _PG3_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B2|1 _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B2|P _PG3_12|_GG|B2|MID_SERIES 0  2e-13
R_PG3_12|_GG|B2|B _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B2|RB _PG3_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B12|1 _PG3_12|_GG|B2 _PG3_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|B12|B _PG3_12|_GG|B2 _PG3_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|B12|RB _PG3_12|_GG|B12|MID_SHUNT _PG3_12|_GG|B3  2.1704737578552e-12
B_PG3_12|_GG|Q2|1 _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q2|P _PG3_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q2|RB _PG3_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|Q1|1 _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q1|P _PG3_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q1|RB _PG3_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_G|I_A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|I_A1|MID  2e-12
I_PG3_12|_AND_G|I_A1|B 0 _PG3_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|I_B1|MID  2e-12
I_PG3_12|_AND_G|I_B1|B 0 _PG3_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q3|B _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|I_Q3|MID  2e-12
I_PG3_12|_AND_G|I_Q3|B 0 _PG3_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_G|I_Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|I_Q2|MID  2e-12
I_PG3_12|_AND_G|I_Q2|B 0 _PG3_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|I_Q1|MID  2e-12
I_PG3_12|_AND_G|I_Q1|B 0 _PG3_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_G|A1|1 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A1|P _PG3_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A1|RB _PG3_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A2|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A2|P _PG3_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A2|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A2|RB _PG3_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A12|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|A12|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|A12|RB _PG3_12|_AND_G|A12|MID_SHUNT _PG3_12|_AND_G|A3  2.1704737578552e-12
B_PG3_12|_AND_G|B1|1 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B1|P _PG3_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B1|RB _PG3_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B2|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B2|P _PG3_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B2|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B2|RB _PG3_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B12|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|B12|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|B12|RB _PG3_12|_AND_G|B12|MID_SHUNT _PG3_12|_AND_G|B3  2.1704737578552e-12
B_PG3_12|_AND_G|Q2|1 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q2|P _PG3_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q2|RB _PG3_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|Q1|1 _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q1|P _PG3_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q1|RB _PG3_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_S0
.print DEVI R_S1
.print DEVI R_S2
.print DEVI R_S3
.print DEVI R_S4
.print V P0_2
.print V IG0_0_TO1
.print V D01
.print V IG2_0
.print V IP1_0
.print V T16
.print V P3_1
.print V P2_1
.print V IG2_0_RX
.print V IP2_0_OUT
.print V IG3_0_RX
.print V S3
.print V IP1_0_RX
.print V IG0_0_RX
.print V T01
.print V IP3_2_OUT_RX
.print V T13
.print V IP2_0_TO2
.print V P0_1_RX
.print V G1_1_TO3
.print V P0_2_RX
.print V S2
.print V G1_1
.print V S0
.print V A1
.print V IP2_0
.print V G0_2_RX
.print V G2_2_RX
.print V IP2_2_OUT
.print V T02
.print V G1_1_RX
.print V IP2_1_OUT
.print V T04
.print V IP0_0
.print V S1
.print V IP3_0_OUT
.print V IP1_1_OUT
.print V G3_2_RX
.print V IG1_0
.print V IP0_0_RX
.print V IP3_0_TO1
.print V IP2_0_RX
.print V IP3_2_OUT
.print V IP3_1_OUT_RX
.print V G1_2_RX
.print V IP2_0_TO3
.print V G0_1_RX
.print V IP1_2_OUT
.print V IP1_1_OUT_RX
.print V IP1_0_OUT
.print V D13
.print V IP3_0
.print V G1_1_TO1
.print V T12
.print V IP1_2_OUT_RX
.print V T07
.print V G2_1_RX
.print V D11
.print V G1_1_TO2
.print V S4
.print V IP2_2_OUT_RX
.print V B1
.print V B3
.print V IG2_0_TO2
.print V B0
.print V G2_2
.print V IP3_0_RX
.print V T06
.print V T14
.print V G3_1
.print V IP2_1_OUT_RX
.print V G0_2
.print V IP1_0_TO1
.print V IG0_0_TO0
.print V T09
.print V D02
.print V IG0_0
.print V T10
.print V T11
.print V T00
.print V D03
.print V G0_1
.print V A3
.print V IG2_0_TO3
.print V G3_1_RX
.print V T15
.print V IG3_0
.print V T08
.print V IP3_1_OUT
.print V A0
.print V P0_1
.print V P3_1_RX
.print V P2_1_RX
.print V T05
.print V G1_2
.print V D12
.print V T03
.print V B2
.print V IG1_0_RX
.print V G3_2
.print V G2_1
.print V A2
