*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM IU=1.25e-05
.PARAM VU=0.0006857
.PARAM LU=2.632e-12
.PARAM JCRIT=0.0001
.PARAM OFFSET1=5e-11
.PARAM TCLOCK=2.5e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT_ADJ JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1.25E-12 2.6E-9
LDRO CLK0 CLK1  PHI0/(4*IC*IC0)
LSUM SUM0 SUM1  PHI0/(4*IC*IC0)
RSUM SUM 0  1
LCARRY CARRY0 CARRY1  PHI0/(4*IC*IC0)
RCARRY CARRY 0  1
RCBAR CBAR 0  1
IDATA|H 0 A  PWL(0 0 -1.55e-11 0 -1.25e-11 0 -9.5e-12 0 4.7e-11 0 5e-11 0 5.3e-11 0 1.095e-10 0 1.125e-10 0 1.155e-10 0 1.72e-10 0 1.75e-10 0 1.78e-10 0 2.345e-10 0 2.375e-10 0 2.405e-10 0 2.97e-10 0 3e-10 0 3.03e-10 0 3.595e-10 0 3.625e-10 0 3.655e-10 0 4.22e-10 0 4.25e-10 0 4.28e-10 0 4.845e-10 0 4.875e-10 0.0007 4.905e-10 0 5.47e-10 0 5.5e-10 0 5.53e-10 0 6.095e-10 0 6.125e-10 0 6.155e-10 0 6.72e-10 0 6.75e-10 0.0007 6.78e-10 0 7.345e-10 0 7.375e-10 0 7.405e-10 0 7.97e-10 0 8e-10 0 8.03e-10 0 8.595e-10 0 8.625e-10 0.0007 8.655e-10 0 9.22e-10 0 9.25e-10 0 9.28e-10 0 9.845e-10 0 9.875e-10 0 9.905e-10 0 1.047e-09 0 1.05e-09 0 1.053e-09 0 1.1095e-09 0 1.1125e-09 0 1.1155e-09 0 1.172e-09 0 1.175e-09 0.0007 1.178e-09 0 1.2345e-09 0 1.2375e-09 0.0007 1.2405e-09 0 1.297e-09 0 1.3e-09 0 1.303e-09 0 1.3595e-09 0 1.3625e-09 0.0007 1.3655e-09 0 1.422e-09 0 1.425e-09 0 1.428e-09 0 1.4845e-09 0 1.4875e-09 0.0007 1.4905e-09 0 1.547e-09 0 1.55e-09 0 1.553e-09 0 1.6095e-09 0 1.6125e-09 0.0007 1.6155e-09 0 1.672e-09 0 1.675e-09 0.0007 1.678e-09 0 1.7345e-09 0 1.7375e-09 0 1.7405e-09 0 1.797e-09 0 1.8e-09 0 1.803e-09 0 1.8595e-09 0 1.8625e-09 0.0007 1.8655e-09 0 1.922e-09 0 1.925e-09 0.0007 1.928e-09 0 1.9845e-09 0 1.9875e-09 0.0007 1.9905e-09 0 2.047e-09 0 2.05e-09 0 2.053e-09 0 2.1095e-09 0 2.1125e-09 0 2.1155e-09 0 2.172e-09 0 2.175e-09 0.0007 2.178e-09 0 2.2345e-09 0 2.2375e-09 0 2.2405e-09 0 2.297e-09 0 2.3e-09 0 2.303e-09 0 2.3595e-09 0 2.3625e-09 0 2.3655e-09 0 2.422e-09 0 2.425e-09 0.0007 2.428e-09 0 2.4845e-09 0 2.4875e-09 0 2.4905e-09 0 2.547e-09 0 2.55e-09 0 2.553e-09 0 2.6095e-09 0 2.6125e-09 0 2.6155e-09 0 2.672e-09 0 2.675e-09 0 2.678e-09 0 2.7345e-09 0 2.7375e-09 0 2.7405e-09 0 2.797e-09 0 2.8e-09 0 2.803e-09 0 2.8595e-09 0 2.8625e-09 0 2.8655e-09 0 2.922e-09 0 2.925e-09 0 2.928e-09 0 2.9845e-09 0 2.9875e-09 0 2.9905e-09 0 3.047e-09 0 3.05e-09 0 3.053e-09 0 3.1095e-09 0 3.1125e-09 0 3.1155e-09 0 3.172e-09 0 3.175e-09 0 3.178e-09 0 3.2345e-09 0 3.2375e-09 0 3.2405e-09 0 3.297e-09 0 3.3e-09 0 3.303e-09 0 3.3595e-09 0 3.3625e-09 0 3.3655e-09 0 3.422e-09 0 3.425e-09 0 3.428e-09 0 3.4845e-09 0 3.4875e-09 0 3.4905e-09 0 3.547e-09 0 3.55e-09 0 3.553e-09 0 3.6095e-09 0 3.6125e-09 0 3.6155e-09 0 3.672e-09 0 3.675e-09 0 3.678e-09 0 3.7345e-09 0 3.7375e-09 0 3.7405e-09 0 3.797e-09 0 3.8e-09 0 3.803e-09 0 3.8595e-09 0 3.8625e-09 0 3.8655e-09 0 3.922e-09 0 3.925e-09 0 3.928e-09 0 3.9845e-09 0 3.9875e-09 0 3.9905e-09 0 4.047e-09 0 4.05e-09 0 4.053e-09 0 4.1095e-09 0 4.1125e-09 0 4.1155e-09 0 4.172e-09 0 4.175e-09 0 4.178e-09 0 4.2345e-09 0 4.2375e-09 0 4.2405e-09 0 4.297e-09 0 4.3e-09 0 4.303e-09 0 4.3595e-09 0 4.3625e-09 0 4.3655e-09 0 4.422e-09 0 4.425e-09 0 4.428e-09 0 4.4845e-09 0 4.4875e-09 0 4.4905e-09 0 4.547e-09 0 4.55e-09 0 4.553e-09 0 4.6095e-09 0 4.6125e-09 0 4.6155e-09 0 4.672e-09 0 4.675e-09 0 4.678e-09 0 4.7345e-09 0 4.7375e-09 0 4.7405e-09 0 4.797e-09 0 4.8e-09 0 4.803e-09 0 4.8595e-09 0 4.8625e-09 0 4.8655e-09 0 4.922e-09 0 4.925e-09 0 4.928e-09 0 4.9845e-09 0 4.9875e-09 0 4.9905e-09 0 5.047e-09 0 5.05e-09 0 5.053e-09 0 5.1095e-09 0 5.1125e-09 0 5.1155e-09 0 5.172e-09 0 5.175e-09 0 5.178e-09 0 5.2345e-09 0 5.2375e-09 0 5.2405e-09 0 5.297e-09 0 5.3e-09 0 5.303e-09 0 5.3595e-09 0 5.3625e-09 0 5.3655e-09 0 5.422e-09 0 5.425e-09 0 5.428e-09 0 5.4845e-09 0 5.4875e-09 0 5.4905e-09 0 5.547e-09 0 5.55e-09 0 5.553e-09 0 5.6095e-09 0 5.6125e-09 0 5.6155e-09 0 5.672e-09 0 5.675e-09 0 5.678e-09 0 5.7345e-09 0 5.7375e-09 0 5.7405e-09 0 5.797e-09 0 5.8e-09 0 5.803e-09 0 5.8595e-09 0 5.8625e-09 0 5.8655e-09 0 5.922e-09 0 5.925e-09 0 5.928e-09 0 5.9845e-09 0 5.9875e-09 0 5.9905e-09 0 6.047e-09 0 6.05e-09 0 6.053e-09 0 6.1095e-09 0 6.1125e-09 0 6.1155e-09 0 6.172e-09 0 6.175e-09 0 6.178e-09 0 6.2345e-09 0 6.2375e-09 0 6.2405e-09 0 6.297e-09 0 6.3e-09 0 6.303e-09 0 6.3595e-09 0 6.3625e-09 0 6.3655e-09 0 6.422e-09 0 6.425e-09 0 6.428e-09 0 6.4845e-09 0 6.4875e-09 0 6.4905e-09 0 6.547e-09 0 6.55e-09 0 6.553e-09 0 6.6095e-09 0 6.6125e-09 0 6.6155e-09 0 6.672e-09 0 6.675e-09 0 6.678e-09 0 6.7345e-09 0 6.7375e-09 0 6.7405e-09 0 6.797e-09 0 6.8e-09 0 6.803e-09 0 6.8595e-09 0 6.8625e-09 0 6.8655e-09 0 6.922e-09 0 6.925e-09 0 6.928e-09 0 6.9845e-09 0 6.9875e-09 0 6.9905e-09 0 7.047e-09 0 7.05e-09 0 7.053e-09 0 7.1095e-09 0 7.1125e-09 0 7.1155e-09 0 7.172e-09 0 7.175e-09 0 7.178e-09 0 7.2345e-09 0 7.2375e-09 0 7.2405e-09 0 7.297e-09 0 7.3e-09 0 7.303e-09 0 7.3595e-09 0 7.3625e-09 0 7.3655e-09 0 7.422e-09 0 7.425e-09 0 7.428e-09 0 7.4845e-09 0 7.4875e-09 0 7.4905e-09 0 7.547e-09 0 7.55e-09 0 7.553e-09 0 7.6095e-09 0 7.6125e-09 0 7.6155e-09 0 7.672e-09 0 7.675e-09 0 7.678e-09 0 7.7345e-09 0 7.7375e-09 0 7.7405e-09 0 7.797e-09 0 7.8e-09 0 7.803e-09 0 7.8595e-09 0 7.8625e-09 0 7.8655e-09 0 7.922e-09 0 7.925e-09 0 7.928e-09 0 7.9845e-09 0 7.9875e-09 0 7.9905e-09 0)
IT1|T 0 CLK0  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.97e-10 0 3e-10 0.0007 3.03e-10 0 5.47e-10 0 5.5e-10 0.0007 5.53e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.297e-09 0 1.3e-09 0.0007 1.303e-09 0 1.547e-09 0 1.55e-09 0.0007 1.553e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.297e-09 0 2.3e-09 0.0007 2.303e-09 0 2.547e-09 0 2.55e-09 0.0007 2.553e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.297e-09 0 3.3e-09 0.0007 3.303e-09 0 3.547e-09 0 3.55e-09 0.0007 3.553e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.297e-09 0 4.3e-09 0.0007 4.303e-09 0 4.547e-09 0 4.55e-09 0.0007 4.553e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.297e-09 0 5.3e-09 0.0007 5.303e-09 0 5.547e-09 0 5.55e-09 0.0007 5.553e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.297e-09 0 6.3e-09 0.0007 6.303e-09 0 6.547e-09 0 6.55e-09 0.0007 6.553e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.297e-09 0 7.3e-09 0.0007 7.303e-09 0 7.547e-09 0 7.55e-09 0.0007 7.553e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.297e-09 0 8.3e-09 0.0007 8.303e-09 0 8.547e-09 0 8.55e-09 0.0007 8.553e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.297e-09 0 9.3e-09 0.0007 9.303e-09 0 9.547e-09 0 9.55e-09 0.0007 9.553e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0297e-08 0 1.03e-08 0.0007 1.0303e-08 0 1.0547e-08 0 1.055e-08 0.0007 1.0553e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1297e-08 0 1.13e-08 0.0007 1.1303e-08 0 1.1547e-08 0 1.155e-08 0.0007 1.1553e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2297e-08 0 1.23e-08 0.0007 1.2303e-08 0 1.2547e-08 0 1.255e-08 0.0007 1.2553e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3297e-08 0 1.33e-08 0.0007 1.3303e-08 0 1.3547e-08 0 1.355e-08 0.0007 1.3553e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4297e-08 0 1.43e-08 0.0007 1.4303e-08 0 1.4547e-08 0 1.455e-08 0.0007 1.4553e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5297e-08 0 1.53e-08 0.0007 1.5303e-08 0 1.5547e-08 0 1.555e-08 0.0007 1.5553e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6297e-08 0 1.63e-08 0.0007 1.6303e-08 0 1.6547e-08 0 1.655e-08 0.0007 1.6553e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7297e-08 0 1.73e-08 0.0007 1.7303e-08 0 1.7547e-08 0 1.755e-08 0.0007 1.7553e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8297e-08 0 1.83e-08 0.0007 1.8303e-08 0 1.8547e-08 0 1.855e-08 0.0007 1.8553e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9297e-08 0 1.93e-08 0.0007 1.9303e-08 0 1.9547e-08 0 1.955e-08 0.0007 1.9553e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0297e-08 0 2.03e-08 0.0007 2.0303e-08 0 2.0547e-08 0 2.055e-08 0.0007 2.0553e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1297e-08 0 2.13e-08 0.0007 2.1303e-08 0 2.1547e-08 0 2.155e-08 0.0007 2.1553e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2297e-08 0 2.23e-08 0.0007 2.2303e-08 0 2.2547e-08 0 2.255e-08 0.0007 2.2553e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3297e-08 0 2.33e-08 0.0007 2.3303e-08 0 2.3547e-08 0 2.355e-08 0.0007 2.3553e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4297e-08 0 2.43e-08 0.0007 2.4303e-08 0 2.4547e-08 0 2.455e-08 0.0007 2.4553e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5297e-08 0 2.53e-08 0.0007 2.5303e-08 0 2.5547e-08 0 2.555e-08 0.0007 2.5553e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6297e-08 0 2.63e-08 0.0007 2.6303e-08 0 2.6547e-08 0 2.655e-08 0.0007 2.6553e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7297e-08 0 2.73e-08 0.0007 2.7303e-08 0 2.7547e-08 0 2.755e-08 0.0007 2.7553e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8297e-08 0 2.83e-08 0.0007 2.8303e-08 0 2.8547e-08 0 2.855e-08 0.0007 2.8553e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9297e-08 0 2.93e-08 0.0007 2.9303e-08 0 2.9547e-08 0 2.955e-08 0.0007 2.9553e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0297e-08 0 3.03e-08 0.0007 3.0303e-08 0 3.0547e-08 0 3.055e-08 0.0007 3.0553e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1297e-08 0 3.13e-08 0.0007 3.1303e-08 0 3.1547e-08 0 3.155e-08 0.0007 3.1553e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2297e-08 0 3.23e-08 0.0007 3.2303e-08 0 3.2547e-08 0 3.255e-08 0.0007 3.2553e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3297e-08 0 3.33e-08 0.0007 3.3303e-08 0 3.3547e-08 0 3.355e-08 0.0007 3.3553e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4297e-08 0 3.43e-08 0.0007 3.4303e-08 0 3.4547e-08 0 3.455e-08 0.0007 3.4553e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5297e-08 0 3.53e-08 0.0007 3.5303e-08 0 3.5547e-08 0 3.555e-08 0.0007 3.5553e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6297e-08 0 3.63e-08 0.0007 3.6303e-08 0 3.6547e-08 0 3.655e-08 0.0007 3.6553e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7297e-08 0 3.73e-08 0.0007 3.7303e-08 0 3.7547e-08 0 3.755e-08 0.0007 3.7553e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8297e-08 0 3.83e-08 0.0007 3.8303e-08 0 3.8547e-08 0 3.855e-08 0.0007 3.8553e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9297e-08 0 3.93e-08 0.0007 3.9303e-08 0 3.9547e-08 0 3.955e-08 0.0007 3.9553e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0297e-08 0 4.03e-08 0.0007 4.0303e-08 0 4.0547e-08 0 4.055e-08 0.0007 4.0553e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1297e-08 0 4.13e-08 0.0007 4.1303e-08 0 4.1547e-08 0 4.155e-08 0.0007 4.1553e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2297e-08 0 4.23e-08 0.0007 4.2303e-08 0 4.2547e-08 0 4.255e-08 0.0007 4.2553e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3297e-08 0 4.33e-08 0.0007 4.3303e-08 0 4.3547e-08 0 4.355e-08 0.0007 4.3553e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4297e-08 0 4.43e-08 0.0007 4.4303e-08 0 4.4547e-08 0 4.455e-08 0.0007 4.4553e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5297e-08 0 4.53e-08 0.0007 4.5303e-08 0 4.5547e-08 0 4.555e-08 0.0007 4.5553e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6297e-08 0 4.63e-08 0.0007 4.6303e-08 0 4.6547e-08 0 4.655e-08 0.0007 4.6553e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7297e-08 0 4.73e-08 0.0007 4.7303e-08 0 4.7547e-08 0 4.755e-08 0.0007 4.7553e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8297e-08 0 4.83e-08 0.0007 4.8303e-08 0 4.8547e-08 0 4.855e-08 0.0007 4.8553e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9297e-08 0 4.93e-08 0.0007 4.9303e-08 0 4.9547e-08 0 4.955e-08 0.0007 4.9553e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0297e-08 0 5.03e-08 0.0007 5.0303e-08 0 5.0547e-08 0 5.055e-08 0.0007 5.0553e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1297e-08 0 5.13e-08 0.0007 5.1303e-08 0 5.1547e-08 0 5.155e-08 0.0007 5.1553e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2297e-08 0 5.23e-08 0.0007 5.2303e-08 0 5.2547e-08 0 5.255e-08 0.0007 5.2553e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3297e-08 0 5.33e-08 0.0007 5.3303e-08 0 5.3547e-08 0 5.355e-08 0.0007 5.3553e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4297e-08 0 5.43e-08 0.0007 5.4303e-08 0 5.4547e-08 0 5.455e-08 0.0007 5.4553e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5297e-08 0 5.53e-08 0.0007 5.5303e-08 0 5.5547e-08 0 5.555e-08 0.0007 5.5553e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6297e-08 0 5.63e-08 0.0007 5.6303e-08 0 5.6547e-08 0 5.655e-08 0.0007 5.6553e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7297e-08 0 5.73e-08 0.0007 5.7303e-08 0 5.7547e-08 0 5.755e-08 0.0007 5.7553e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8297e-08 0 5.83e-08 0.0007 5.8303e-08 0 5.8547e-08 0 5.855e-08 0.0007 5.8553e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9297e-08 0 5.93e-08 0.0007 5.9303e-08 0 5.9547e-08 0 5.955e-08 0.0007 5.9553e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0297e-08 0 6.03e-08 0.0007 6.0303e-08 0 6.0547e-08 0 6.055e-08 0.0007 6.0553e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1297e-08 0 6.13e-08 0.0007 6.1303e-08 0 6.1547e-08 0 6.155e-08 0.0007 6.1553e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2297e-08 0 6.23e-08 0.0007 6.2303e-08 0 6.2547e-08 0 6.255e-08 0.0007 6.2553e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3297e-08 0 6.33e-08 0.0007 6.3303e-08 0 6.3547e-08 0 6.355e-08 0.0007 6.3553e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4297e-08 0 6.43e-08 0.0007 6.4303e-08 0 6.4547e-08 0 6.455e-08 0.0007 6.4553e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5297e-08 0 6.53e-08 0.0007 6.5303e-08 0 6.5547e-08 0 6.555e-08 0.0007 6.5553e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6297e-08 0 6.63e-08 0.0007 6.6303e-08 0 6.6547e-08 0 6.655e-08 0.0007 6.6553e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7297e-08 0 6.73e-08 0.0007 6.7303e-08 0 6.7547e-08 0 6.755e-08 0.0007 6.7553e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8297e-08 0 6.83e-08 0.0007 6.8303e-08 0 6.8547e-08 0 6.855e-08 0.0007 6.8553e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9297e-08 0 6.93e-08 0.0007 6.9303e-08 0 6.9547e-08 0 6.955e-08 0.0007 6.9553e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0297e-08 0 7.03e-08 0.0007 7.0303e-08 0 7.0547e-08 0 7.055e-08 0.0007 7.0553e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1297e-08 0 7.13e-08 0.0007 7.1303e-08 0 7.1547e-08 0 7.155e-08 0.0007 7.1553e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2297e-08 0 7.23e-08 0.0007 7.2303e-08 0 7.2547e-08 0 7.255e-08 0.0007 7.2553e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3297e-08 0 7.33e-08 0.0007 7.3303e-08 0 7.3547e-08 0 7.355e-08 0.0007 7.3553e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4297e-08 0 7.43e-08 0.0007 7.4303e-08 0 7.4547e-08 0 7.455e-08 0.0007 7.4553e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5297e-08 0 7.53e-08 0.0007 7.5303e-08 0 7.5547e-08 0 7.555e-08 0.0007 7.5553e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6297e-08 0 7.63e-08 0.0007 7.6303e-08 0 7.6547e-08 0 7.655e-08 0.0007 7.6553e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7297e-08 0 7.73e-08 0.0007 7.7303e-08 0 7.7547e-08 0 7.755e-08 0.0007 7.7553e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8297e-08 0 7.83e-08 0.0007 7.8303e-08 0 7.8547e-08 0 7.855e-08 0.0007 7.8553e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9297e-08 0 7.93e-08 0.0007 7.9303e-08 0 7.9547e-08 0 7.955e-08 0.0007 7.9553e-08 0 7.9797e-08 0 7.98e-08 0.0007 7.9803e-08 0 8.0047e-08 0 8.005e-08 0.0007 8.0053e-08 0 8.0297e-08 0 8.03e-08 0.0007 8.0303e-08 0 8.0547e-08 0 8.055e-08 0.0007 8.0553e-08 0 8.0797e-08 0 8.08e-08 0.0007 8.0803e-08 0 8.1047e-08 0 8.105e-08 0.0007 8.1053e-08 0 8.1297e-08 0 8.13e-08 0.0007 8.1303e-08 0 8.1547e-08 0 8.155e-08 0.0007 8.1553e-08 0 8.1797e-08 0 8.18e-08 0.0007 8.1803e-08 0 8.2047e-08 0 8.205e-08 0.0007 8.2053e-08 0 8.2297e-08 0 8.23e-08 0.0007 8.2303e-08 0 8.2547e-08 0 8.255e-08 0.0007 8.2553e-08 0 8.2797e-08 0 8.28e-08 0.0007 8.2803e-08 0 8.3047e-08 0 8.305e-08 0.0007 8.3053e-08 0 8.3297e-08 0 8.33e-08 0.0007 8.3303e-08 0 8.3547e-08 0 8.355e-08 0.0007 8.3553e-08 0 8.3797e-08 0 8.38e-08 0.0007 8.3803e-08 0 8.4047e-08 0 8.405e-08 0.0007 8.4053e-08 0 8.4297e-08 0 8.43e-08 0.0007 8.4303e-08 0 8.4547e-08 0 8.455e-08 0.0007 8.4553e-08 0 8.4797e-08 0 8.48e-08 0.0007 8.4803e-08 0 8.5047e-08 0 8.505e-08 0.0007 8.5053e-08 0 8.5297e-08 0 8.53e-08 0.0007 8.5303e-08 0 8.5547e-08 0 8.555e-08 0.0007 8.5553e-08 0 8.5797e-08 0 8.58e-08 0.0007 8.5803e-08 0 8.6047e-08 0 8.605e-08 0.0007 8.6053e-08 0 8.6297e-08 0 8.63e-08 0.0007 8.6303e-08 0 8.6547e-08 0 8.655e-08 0.0007 8.6553e-08 0 8.6797e-08 0 8.68e-08 0.0007 8.6803e-08 0 8.7047e-08 0 8.705e-08 0.0007 8.7053e-08 0 8.7297e-08 0 8.73e-08 0.0007 8.7303e-08 0 8.7547e-08 0 8.755e-08 0.0007 8.7553e-08 0 8.7797e-08 0 8.78e-08 0.0007 8.7803e-08 0 8.8047e-08 0 8.805e-08 0.0007 8.8053e-08 0 8.8297e-08 0 8.83e-08 0.0007 8.8303e-08 0 8.8547e-08 0 8.855e-08 0.0007 8.8553e-08 0 8.8797e-08 0 8.88e-08 0.0007 8.8803e-08 0 8.9047e-08 0 8.905e-08 0.0007 8.9053e-08 0 8.9297e-08 0 8.93e-08 0.0007 8.9303e-08 0 8.9547e-08 0 8.955e-08 0.0007 8.9553e-08 0 8.9797e-08 0 8.98e-08 0.0007 8.9803e-08 0 9.0047e-08 0 9.005e-08 0.0007 9.0053e-08 0 9.0297e-08 0 9.03e-08 0.0007 9.0303e-08 0 9.0547e-08 0 9.055e-08 0.0007 9.0553e-08 0 9.0797e-08 0 9.08e-08 0.0007 9.0803e-08 0 9.1047e-08 0 9.105e-08 0.0007 9.1053e-08 0 9.1297e-08 0 9.13e-08 0.0007 9.1303e-08 0 9.1547e-08 0 9.155e-08 0.0007 9.1553e-08 0 9.1797e-08 0 9.18e-08 0.0007 9.1803e-08 0 9.2047e-08 0 9.205e-08 0.0007 9.2053e-08 0 9.2297e-08 0 9.23e-08 0.0007 9.2303e-08 0 9.2547e-08 0 9.255e-08 0.0007 9.2553e-08 0 9.2797e-08 0 9.28e-08 0.0007 9.2803e-08 0 9.3047e-08 0 9.305e-08 0.0007 9.3053e-08 0 9.3297e-08 0 9.33e-08 0.0007 9.3303e-08 0 9.3547e-08 0 9.355e-08 0.0007 9.3553e-08 0 9.3797e-08 0 9.38e-08 0.0007 9.3803e-08 0 9.4047e-08 0 9.405e-08 0.0007 9.4053e-08 0 9.4297e-08 0 9.43e-08 0.0007 9.4303e-08 0 9.4547e-08 0 9.455e-08 0.0007 9.4553e-08 0 9.4797e-08 0 9.48e-08 0.0007 9.4803e-08 0 9.5047e-08 0 9.505e-08 0.0007 9.5053e-08 0 9.5297e-08 0 9.53e-08 0.0007 9.5303e-08 0 9.5547e-08 0 9.555e-08 0.0007 9.5553e-08 0 9.5797e-08 0 9.58e-08 0.0007 9.5803e-08 0 9.6047e-08 0 9.605e-08 0.0007 9.6053e-08 0 9.6297e-08 0 9.63e-08 0.0007 9.6303e-08 0 9.6547e-08 0 9.655e-08 0.0007 9.6553e-08 0 9.6797e-08 0 9.68e-08 0.0007 9.6803e-08 0 9.7047e-08 0 9.705e-08 0.0007 9.7053e-08 0 9.7297e-08 0 9.73e-08 0.0007 9.7303e-08 0 9.7547e-08 0 9.755e-08 0.0007 9.7553e-08 0 9.7797e-08 0 9.78e-08 0.0007 9.7803e-08 0 9.8047e-08 0 9.805e-08 0.0007 9.8053e-08 0 9.8297e-08 0 9.83e-08 0.0007 9.8303e-08 0 9.8547e-08 0 9.855e-08 0.0007 9.8553e-08 0 9.8797e-08 0 9.88e-08 0.0007 9.8803e-08 0 9.9047e-08 0 9.905e-08 0.0007 9.9053e-08 0 9.9297e-08 0 9.93e-08 0.0007 9.9303e-08 0 9.9547e-08 0 9.955e-08 0.0007 9.9553e-08 0)
BT_PTL|1 T_PTL|1 T_PTL|2 JJMIT AREA=2.5
BT_PTL|2 T_PTL|4 T_PTL|5 JJMIT AREA=2.5
BT_PTL|3 T_PTL|7 T_PTL|8 JJMIT AREA=2.5
BT_PTL|4 T_PTL|10 T_PTL|11 JJMIT AREA=2.5
IT_PTL|B1 0 T_PTL|3  PWL(0 0 5e-12 0.000175)
IT_PTL|B2 0 T_PTL|6  PWL(0 0 5e-12 0.0002375)
IT_PTL|B3 0 T_PTL|9  PWL(0 0 5e-12 0.0002375)
IT_PTL|B4 0 T_PTL|12  PWL(0 0 5e-12 0.000175)
LT_PTL|1 CLK1 T_PTL|1  2.067833848e-12
LT_PTL|2 T_PTL|1 T_PTL|4  4.135667696e-12
LT_PTL|3 T_PTL|4 T_PTL|7  4.135667696e-12
LT_PTL|4 T_PTL|7 T_PTL|10  4.135667696e-12
LT_PTL|5 T_PTL|10 CLK  2.067833848e-12
LT_PTL|P1 T_PTL|2 0  5e-13
LT_PTL|P2 T_PTL|5 0  5e-13
LT_PTL|P3 T_PTL|8 0  5e-13
LT_PTL|P4 T_PTL|11 0  5e-13
LT_PTL|B1 T_PTL|1 T_PTL|3  2e-12
LT_PTL|B2 T_PTL|4 T_PTL|6  2e-12
LT_PTL|B3 T_PTL|7 T_PTL|9  2e-12
LT_PTL|B4 T_PTL|10 T_PTL|12  2e-12
RT_PTL|B1 T_PTL|1 T_PTL|101  2.7439617672
RT_PTL|B2 T_PTL|4 T_PTL|104  2.7439617672
RT_PTL|B3 T_PTL|7 T_PTL|107  2.7439617672
RT_PTL|B4 T_PTL|10 T_PTL|110  2.7439617672
LT_PTL|RB1 T_PTL|101 0  2.050338398468e-12
LT_PTL|RB2 T_PTL|104 0  2.050338398468e-12
LT_PTL|RB3 T_PTL|107 0  2.050338398468e-12
LT_PTL|RB4 T_PTL|110 0  2.050338398468e-12
L_TFF|6 CLK _TFF|1  2.63e-12
B_TFF|11 _TFF|1 _TFF|2 JJMIT_ADJ AREA=2.2
B_TFF|10 _TFF|2 0 JJMIT_ADJ AREA=2.9999999999999996
L_TFF|8 _TFF|2 SUM0  5.26e-12
B_TFF|12 _TFF|2 _TFF|4 JJMIT_ADJ AREA=1.25
B_TFF|6 _TFF|4 _TFF|6 JJMIT_ADJ AREA=1.9
L_TFF|1 _TFF|3 _TFF|4  5.26e-12
L_TFF|3 _TFF|3 CBAR  5.26e-12
B_TFF|1 _TFF|3 0 JJMIT_ADJ AREA=2.5
B_TFF|2 _TFF|3 _TFF|5 JJMIT_ADJ AREA=2.5
B_TFF|5 _TFF|5 _TFF|6 JJMIT_ADJ AREA=1.25
L_TFF|4 _TFF|6 CARRY0  5.26e-12
B_TFF|4 _TFF|6 0 JJMIT_ADJ AREA=1.25
L_TFF|2 _TFF|5 _TFF|7  1.3e-12
B_TFF|3 _TFF|7 0 JJMIT_ADJ AREA=2.5
L_TFF|7 _TFF|7 A  3.9e-12
BSUM|1 SUM|1 SUM|2 JJMIT AREA=2.5
BSUM|2 SUM|4 SUM|5 JJMIT AREA=2.5
BSUM|3 SUM|7 SUM|8 JJMIT AREA=2.5
BSUM|4 SUM|10 SUM|11 JJMIT AREA=2.5
ISUM|B1 0 SUM|3  PWL(0 0 5e-12 0.000175)
ISUM|B2 0 SUM|6  PWL(0 0 5e-12 0.0002375)
ISUM|B3 0 SUM|9  PWL(0 0 5e-12 0.0002375)
ISUM|B4 0 SUM|12  PWL(0 0 5e-12 0.000175)
LSUM|1 SUM1 SUM|1  2.067833848e-12
LSUM|2 SUM|1 SUM|4  4.135667696e-12
LSUM|3 SUM|4 SUM|7  4.135667696e-12
LSUM|4 SUM|7 SUM|10  4.135667696e-12
LSUM|5 SUM|10 SUM  2.067833848e-12
LSUM|P1 SUM|2 0  5e-13
LSUM|P2 SUM|5 0  5e-13
LSUM|P3 SUM|8 0  5e-13
LSUM|P4 SUM|11 0  5e-13
LSUM|B1 SUM|1 SUM|3  2e-12
LSUM|B2 SUM|4 SUM|6  2e-12
LSUM|B3 SUM|7 SUM|9  2e-12
LSUM|B4 SUM|10 SUM|12  2e-12
RSUM|B1 SUM|1 SUM|101  2.7439617672
RSUM|B2 SUM|4 SUM|104  2.7439617672
RSUM|B3 SUM|7 SUM|107  2.7439617672
RSUM|B4 SUM|10 SUM|110  2.7439617672
LSUM|RB1 SUM|101 0  2.050338398468e-12
LSUM|RB2 SUM|104 0  2.050338398468e-12
LSUM|RB3 SUM|107 0  2.050338398468e-12
LSUM|RB4 SUM|110 0  2.050338398468e-12
BQ|1 Q|1 Q|2 JJMIT AREA=2.5
BQ|2 Q|4 Q|5 JJMIT AREA=2.5
BQ|3 Q|7 Q|8 JJMIT AREA=2.5
BQ|4 Q|10 Q|11 JJMIT AREA=2.5
IQ|B1 0 Q|3  PWL(0 0 5e-12 0.000175)
IQ|B2 0 Q|6  PWL(0 0 5e-12 0.0002375)
IQ|B3 0 Q|9  PWL(0 0 5e-12 0.0002375)
IQ|B4 0 Q|12  PWL(0 0 5e-12 0.000175)
LQ|1 CARRY1 Q|1  2.067833848e-12
LQ|2 Q|1 Q|4  4.135667696e-12
LQ|3 Q|4 Q|7  4.135667696e-12
LQ|4 Q|7 Q|10  4.135667696e-12
LQ|5 Q|10 CARRY  2.067833848e-12
LQ|P1 Q|2 0  5e-13
LQ|P2 Q|5 0  5e-13
LQ|P3 Q|8 0  5e-13
LQ|P4 Q|11 0  5e-13
LQ|B1 Q|1 Q|3  2e-12
LQ|B2 Q|4 Q|6  2e-12
LQ|B3 Q|7 Q|9  2e-12
LQ|B4 Q|10 Q|12  2e-12
RQ|B1 Q|1 Q|101  2.7439617672
RQ|B2 Q|4 Q|104  2.7439617672
RQ|B3 Q|7 Q|107  2.7439617672
RQ|B4 Q|10 Q|110  2.7439617672
LQ|RB1 Q|101 0  2.050338398468e-12
LQ|RB2 Q|104 0  2.050338398468e-12
LQ|RB3 Q|107 0  2.050338398468e-12
LQ|RB4 Q|110 0  2.050338398468e-12
L_TFF|I1|B _TFF|3 _TFF|I1|MID  2e-12
I_TFF|I1|B 0 _TFF|I1|MID  PWL(0 0 5e-12 0.00019)
L_TFF|I2|B _TFF|7 _TFF|I2|MID  2e-12
I_TFF|I2|B 0 _TFF|I2|MID  PWL(0 0 5e-12 0.00019)
.print DEVI LDRO
.print DEVI LSUM
.print DEVI RSUM
.print DEVI LCARRY
.print DEVI RCARRY
.print DEVI RCBAR
.print DEVI IDATA|H
.print DEVI IT1|T
.print DEVI BT_PTL|1
.print DEVI BT_PTL|2
.print DEVI BT_PTL|3
.print DEVI BT_PTL|4
.print DEVI IT_PTL|B1
.print DEVI IT_PTL|B2
.print DEVI IT_PTL|B3
.print DEVI IT_PTL|B4
.print DEVI LT_PTL|1
.print DEVI LT_PTL|2
.print DEVI LT_PTL|3
.print DEVI LT_PTL|4
.print DEVI LT_PTL|5
.print DEVI LT_PTL|P1
.print DEVI LT_PTL|P2
.print DEVI LT_PTL|P3
.print DEVI LT_PTL|P4
.print DEVI LT_PTL|B1
.print DEVI LT_PTL|B2
.print DEVI LT_PTL|B3
.print DEVI LT_PTL|B4
.print DEVI RT_PTL|B1
.print DEVI RT_PTL|B2
.print DEVI RT_PTL|B3
.print DEVI RT_PTL|B4
.print DEVI LT_PTL|RB1
.print DEVI LT_PTL|RB2
.print DEVI LT_PTL|RB3
.print DEVI LT_PTL|RB4
.print DEVI L_TFF|6
.print DEVI B_TFF|11
.print DEVI B_TFF|10
.print DEVI L_TFF|8
.print DEVI B_TFF|12
.print DEVI B_TFF|6
.print DEVI L_TFF|1
.print DEVI L_TFF|3
.print DEVI B_TFF|1
.print DEVI B_TFF|2
.print DEVI B_TFF|5
.print DEVI L_TFF|4
.print DEVI B_TFF|4
.print DEVI L_TFF|2
.print DEVI B_TFF|3
.print DEVI L_TFF|7
.print DEVI BSUM|1
.print DEVI BSUM|2
.print DEVI BSUM|3
.print DEVI BSUM|4
.print DEVI ISUM|B1
.print DEVI ISUM|B2
.print DEVI ISUM|B3
.print DEVI ISUM|B4
.print DEVI LSUM|1
.print DEVI LSUM|2
.print DEVI LSUM|3
.print DEVI LSUM|4
.print DEVI LSUM|5
.print DEVI LSUM|P1
.print DEVI LSUM|P2
.print DEVI LSUM|P3
.print DEVI LSUM|P4
.print DEVI LSUM|B1
.print DEVI LSUM|B2
.print DEVI LSUM|B3
.print DEVI LSUM|B4
.print DEVI RSUM|B1
.print DEVI RSUM|B2
.print DEVI RSUM|B3
.print DEVI RSUM|B4
.print DEVI LSUM|RB1
.print DEVI LSUM|RB2
.print DEVI LSUM|RB3
.print DEVI LSUM|RB4
.print DEVI BQ|1
.print DEVI BQ|2
.print DEVI BQ|3
.print DEVI BQ|4
.print DEVI IQ|B1
.print DEVI IQ|B2
.print DEVI IQ|B3
.print DEVI IQ|B4
.print DEVI LQ|1
.print DEVI LQ|2
.print DEVI LQ|3
.print DEVI LQ|4
.print DEVI LQ|5
.print DEVI LQ|P1
.print DEVI LQ|P2
.print DEVI LQ|P3
.print DEVI LQ|P4
.print DEVI LQ|B1
.print DEVI LQ|B2
.print DEVI LQ|B3
.print DEVI LQ|B4
.print DEVI RQ|B1
.print DEVI RQ|B2
.print DEVI RQ|B3
.print DEVI RQ|B4
.print DEVI LQ|RB1
.print DEVI LQ|RB2
.print DEVI LQ|RB3
.print DEVI LQ|RB4
.print V T_PTL|1
.print V SUM1
.print V _TFF|1
.print V Q|5
.print V T_PTL|107
.print V T_PTL|11
.print V _TFF|3
.print V SUM|10
.print V SUM|6
.print V T_PTL|104
.print V _TFF|7
.print V Q|11
.print V Q|104
.print V CLK1
.print V T_PTL|9
.print V Q|10
.print V SUM|8
.print V SUM|9
.print V Q|101
.print V CARRY
.print V SUM|2
.print V SUM|101
.print V SUM|110
.print V Q|1
.print V T_PTL|4
.print V CARRY0
.print V T_PTL|8
.print V SUM|12
.print V SUM|107
.print V Q|6
.print V _TFF|6
.print V SUM|7
.print V _TFF|4
.print V CLK
.print V Q|110
.print V SUM
.print V T_PTL|3
.print V CBAR
.print V CARRY1
.print V T_PTL|12
.print V _TFF|5
.print V Q|3
.print V Q|107
.print V Q|7
.print V T_PTL|10
.print V A
.print V SUM|1
.print V T_PTL|6
.print V Q|8
.print V SUM|3
.print V Q|9
.print V SUM|11
.print V T_PTL|101
.print V SUM|5
.print V SUM|4
.print V T_PTL|2
.print V T_PTL|110
.print V _TFF|2
.print V Q|2
.print V Q|4
.print V T_PTL|5
.print V CLK0
.print V SUM|104
.print V Q|12
.print V T_PTL|7
.print V SUM0
.print DEVP BT_PTL|1
.print DEVP BT_PTL|2
.print DEVP BT_PTL|3
.print DEVP BT_PTL|4
.print DEVP B_TFF|11
.print DEVP B_TFF|10
.print DEVP B_TFF|12
.print DEVP B_TFF|6
.print DEVP B_TFF|1
.print DEVP B_TFF|2
.print DEVP B_TFF|5
.print DEVP B_TFF|4
.print DEVP B_TFF|3
.print DEVP BSUM|1
.print DEVP BSUM|2
.print DEVP BSUM|3
.print DEVP BSUM|4
.print DEVP BQ|1
.print DEVP BQ|2
.print DEVP BQ|3
.print DEVP BQ|4
