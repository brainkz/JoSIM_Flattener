


*
.include /Users/brainkz/Documents/GitHub/SFQ_gate_Exploration/jj_library.cir
.include /Users/brainkz/Documents/GitHub/SFQ/sunmagnetics_library.cir
* .include /Users/brainkz/Documents/GitHub/SFQ_gate_Exploration/pulses.cir

.param offset1=5e-11
.param tclock=10e-11

Xt1       clk  clk_sig    clk_offset=offset1 factor=1    Tck=tclock

X_tff clk q0 tff

L1 q0 q1 Phi0/(4*IC*Ic0) 
X_buf q1 q LSMITLL_BUFF

ROUT q  0  1  

.tran 0.1e-12 1e-09

.end
