*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=1e-11
.PARAM TCLOCK=2e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 2.5E-12 48E-10
RS0 S0 0  1
RS1 S1 0  1
RS2 S2 0  1
IT2|T 0 CLK2  PWL(0 0 7e-12 0 1e-11 0.005 1.3e-11 0 2.07e-10 0 2.1e-10 0.005 2.13e-10 0 4.07e-10 0 4.1e-10 0.005 4.13e-10 0 6.07e-10 0 6.1e-10 0.005 6.13e-10 0 8.07e-10 0 8.1e-10 0.005 8.13e-10 0 1.007e-09 0 1.01e-09 0.005 1.013e-09 0 1.207e-09 0 1.21e-09 0.005 1.213e-09 0 1.407e-09 0 1.41e-09 0.005 1.413e-09 0 1.607e-09 0 1.61e-09 0.005 1.613e-09 0 1.807e-09 0 1.81e-09 0.005 1.813e-09 0 2.007e-09 0 2.01e-09 0.005 2.013e-09 0 2.207e-09 0 2.21e-09 0.005 2.213e-09 0 2.407e-09 0 2.41e-09 0.005 2.413e-09 0 2.607e-09 0 2.61e-09 0.005 2.613e-09 0 2.807e-09 0 2.81e-09 0.005 2.813e-09 0 3.007e-09 0 3.01e-09 0.005 3.013e-09 0 3.207e-09 0 3.21e-09 0.005 3.213e-09 0 3.407e-09 0 3.41e-09 0.005 3.413e-09 0 3.607e-09 0 3.61e-09 0.005 3.613e-09 0 3.807e-09 0 3.81e-09 0.005 3.813e-09 0 4.007e-09 0 4.01e-09 0.005 4.013e-09 0 4.207e-09 0 4.21e-09 0.005 4.213e-09 0 4.407e-09 0 4.41e-09 0.005 4.413e-09 0 4.607e-09 0 4.61e-09 0.005 4.613e-09 0 4.807e-09 0 4.81e-09 0.005 4.813e-09 0 5.007e-09 0 5.01e-09 0.005 5.013e-09 0 5.207e-09 0 5.21e-09 0.005 5.213e-09 0 5.407e-09 0 5.41e-09 0.005 5.413e-09 0 5.607e-09 0 5.61e-09 0.005 5.613e-09 0 5.807e-09 0 5.81e-09 0.005 5.813e-09 0 6.007e-09 0 6.01e-09 0.005 6.013e-09 0 6.207e-09 0 6.21e-09 0.005 6.213e-09 0 6.407e-09 0 6.41e-09 0.005 6.413e-09 0 6.607e-09 0 6.61e-09 0.005 6.613e-09 0 6.807e-09 0 6.81e-09 0.005 6.813e-09 0 7.007e-09 0 7.01e-09 0.005 7.013e-09 0 7.207e-09 0 7.21e-09 0.005 7.213e-09 0 7.407e-09 0 7.41e-09 0.005 7.413e-09 0 7.607e-09 0 7.61e-09 0.005 7.613e-09 0)
IT1|T 0 CLK1  PWL(0 0 1.7e-11 0 2e-11 0.005 2.3e-11 0 2.17e-10 0 2.2e-10 0.005 2.23e-10 0 4.17e-10 0 4.2e-10 0.005 4.23e-10 0 6.17e-10 0 6.2e-10 0.005 6.23e-10 0 8.17e-10 0 8.2e-10 0.005 8.23e-10 0 1.017e-09 0 1.02e-09 0.005 1.023e-09 0 1.217e-09 0 1.22e-09 0.005 1.223e-09 0 1.417e-09 0 1.42e-09 0.005 1.423e-09 0 1.617e-09 0 1.62e-09 0.005 1.623e-09 0 1.817e-09 0 1.82e-09 0.005 1.823e-09 0 2.017e-09 0 2.02e-09 0.005 2.023e-09 0 2.217e-09 0 2.22e-09 0.005 2.223e-09 0 2.417e-09 0 2.42e-09 0.005 2.423e-09 0 2.617e-09 0 2.62e-09 0.005 2.623e-09 0 2.817e-09 0 2.82e-09 0.005 2.823e-09 0 3.017e-09 0 3.02e-09 0.005 3.023e-09 0 3.217e-09 0 3.22e-09 0.005 3.223e-09 0 3.417e-09 0 3.42e-09 0.005 3.423e-09 0 3.617e-09 0 3.62e-09 0.005 3.623e-09 0 3.817e-09 0 3.82e-09 0.005 3.823e-09 0 4.017e-09 0 4.02e-09 0.005 4.023e-09 0 4.217e-09 0 4.22e-09 0.005 4.223e-09 0 4.417e-09 0 4.42e-09 0.005 4.423e-09 0 4.617e-09 0 4.62e-09 0.005 4.623e-09 0 4.817e-09 0 4.82e-09 0.005 4.823e-09 0 5.017e-09 0 5.02e-09 0.005 5.023e-09 0 5.217e-09 0 5.22e-09 0.005 5.223e-09 0 5.417e-09 0 5.42e-09 0.005 5.423e-09 0 5.617e-09 0 5.62e-09 0.005 5.623e-09 0 5.817e-09 0 5.82e-09 0.005 5.823e-09 0 6.017e-09 0 6.02e-09 0.005 6.023e-09 0 6.217e-09 0 6.22e-09 0.005 6.223e-09 0 6.417e-09 0 6.42e-09 0.005 6.423e-09 0 6.617e-09 0 6.62e-09 0.005 6.623e-09 0 6.817e-09 0 6.82e-09 0.005 6.823e-09 0 7.017e-09 0 7.02e-09 0.005 7.023e-09 0 7.217e-09 0 7.22e-09 0.005 7.223e-09 0 7.417e-09 0 7.42e-09 0.005 7.423e-09 0 7.617e-09 0 7.62e-09 0.005 7.623e-09 0)
IT0|T 0 CLK0  PWL(0 0 2.7e-11 0 3e-11 0.005 3.3e-11 0 2.27e-10 0 2.3e-10 0.005 2.33e-10 0 4.27e-10 0 4.3e-10 0.005 4.33e-10 0 6.27e-10 0 6.3e-10 0.005 6.33e-10 0 8.27e-10 0 8.3e-10 0.005 8.33e-10 0 1.027e-09 0 1.03e-09 0.005 1.033e-09 0 1.227e-09 0 1.23e-09 0.005 1.233e-09 0 1.427e-09 0 1.43e-09 0.005 1.433e-09 0 1.627e-09 0 1.63e-09 0.005 1.633e-09 0 1.827e-09 0 1.83e-09 0.005 1.833e-09 0 2.027e-09 0 2.03e-09 0.005 2.033e-09 0 2.227e-09 0 2.23e-09 0.005 2.233e-09 0 2.427e-09 0 2.43e-09 0.005 2.433e-09 0 2.627e-09 0 2.63e-09 0.005 2.633e-09 0 2.827e-09 0 2.83e-09 0.005 2.833e-09 0 3.027e-09 0 3.03e-09 0.005 3.033e-09 0 3.227e-09 0 3.23e-09 0.005 3.233e-09 0 3.427e-09 0 3.43e-09 0.005 3.433e-09 0 3.627e-09 0 3.63e-09 0.005 3.633e-09 0 3.827e-09 0 3.83e-09 0.005 3.833e-09 0 4.027e-09 0 4.03e-09 0.005 4.033e-09 0 4.227e-09 0 4.23e-09 0.005 4.233e-09 0 4.427e-09 0 4.43e-09 0.005 4.433e-09 0 4.627e-09 0 4.63e-09 0.005 4.633e-09 0 4.827e-09 0 4.83e-09 0.005 4.833e-09 0 5.027e-09 0 5.03e-09 0.005 5.033e-09 0 5.227e-09 0 5.23e-09 0.005 5.233e-09 0 5.427e-09 0 5.43e-09 0.005 5.433e-09 0 5.627e-09 0 5.63e-09 0.005 5.633e-09 0 5.827e-09 0 5.83e-09 0.005 5.833e-09 0 6.027e-09 0 6.03e-09 0.005 6.033e-09 0 6.227e-09 0 6.23e-09 0.005 6.233e-09 0 6.427e-09 0 6.43e-09 0.005 6.433e-09 0 6.627e-09 0 6.63e-09 0.005 6.633e-09 0 6.827e-09 0 6.83e-09 0.005 6.833e-09 0 7.027e-09 0 7.03e-09 0.005 7.033e-09 0 7.227e-09 0 7.23e-09 0.005 7.233e-09 0 7.427e-09 0 7.43e-09 0.005 7.433e-09 0 7.627e-09 0 7.63e-09 0.005 7.633e-09 0)
IDATA_A0|A 0 A0I  PWL(0 0 2.47e-10 0 2.5e-10 0.0005 2.53e-10 0 6.47e-10 0 6.5e-10 0.0005 6.53e-10 0 1.047e-09 0 1.05e-09 0.0005 1.053e-09 0 1.447e-09 0 1.45e-09 0.0005 1.453e-09 0 1.847e-09 0 1.85e-09 0.0005 1.853e-09 0 2.247e-09 0 2.25e-09 0.0005 2.253e-09 0 2.647e-09 0 2.65e-09 0.0005 2.653e-09 0 3.047e-09 0 3.05e-09 0.0005 3.053e-09 0 3.447e-09 0 3.45e-09 0.0005 3.453e-09 0 3.847e-09 0 3.85e-09 0.0005 3.853e-09 0 4.247e-09 0 4.25e-09 0.0005 4.253e-09 0 4.647e-09 0 4.65e-09 0.0005 4.653e-09 0 5.047e-09 0 5.05e-09 0.0005 5.053e-09 0 5.447e-09 0 5.45e-09 0.0005 5.453e-09 0 5.847e-09 0 5.85e-09 0.0005 5.853e-09 0 6.247e-09 0 6.25e-09 0.0005 6.253e-09 0 6.647e-09 0 6.65e-09 0.0005 6.653e-09 0 7.047e-09 0 7.05e-09 0.0005 7.053e-09 0 7.447e-09 0 7.45e-09 0.0005 7.453e-09 0)
IDATA_B0|B 0 B0I  PWL(0 0 4.87e-10 0 4.9e-10 0.0005 4.93e-10 0 6.87e-10 0 6.9e-10 0.0005 6.93e-10 0 1.287e-09 0 1.29e-09 0.0005 1.293e-09 0 1.487e-09 0 1.49e-09 0.0005 1.493e-09 0 2.087e-09 0 2.09e-09 0.0005 2.093e-09 0 2.287e-09 0 2.29e-09 0.0005 2.293e-09 0 2.887e-09 0 2.89e-09 0.0005 2.893e-09 0 3.087e-09 0 3.09e-09 0.0005 3.093e-09 0 3.687e-09 0 3.69e-09 0.0005 3.693e-09 0 3.887e-09 0 3.89e-09 0.0005 3.893e-09 0 4.487e-09 0 4.49e-09 0.0005 4.493e-09 0 4.687e-09 0 4.69e-09 0.0005 4.693e-09 0 5.287e-09 0 5.29e-09 0.0005 5.293e-09 0 5.487e-09 0 5.49e-09 0.0005 5.493e-09 0 6.087e-09 0 6.09e-09 0.0005 6.093e-09 0 6.287e-09 0 6.29e-09 0.0005 6.293e-09 0 6.887e-09 0 6.89e-09 0.0005 6.893e-09 0 7.087e-09 0 7.09e-09 0.0005 7.093e-09 0 7.687e-09 0 7.69e-09 0.0005 7.693e-09 0)
IDATA_A1|C 0 A1I  PWL(0 0 9.27e-10 0 9.3e-10 0.0005 9.33e-10 0 1.127e-09 0 1.13e-09 0.0005 1.133e-09 0 1.327e-09 0 1.33e-09 0.0005 1.333e-09 0 1.527e-09 0 1.53e-09 0.0005 1.533e-09 0 2.527e-09 0 2.53e-09 0.0005 2.533e-09 0 2.727e-09 0 2.73e-09 0.0005 2.733e-09 0 2.927e-09 0 2.93e-09 0.0005 2.933e-09 0 3.127e-09 0 3.13e-09 0.0005 3.133e-09 0 4.127e-09 0 4.13e-09 0.0005 4.133e-09 0 4.327e-09 0 4.33e-09 0.0005 4.333e-09 0 4.527e-09 0 4.53e-09 0.0005 4.533e-09 0 4.727e-09 0 4.73e-09 0.0005 4.733e-09 0 5.727e-09 0 5.73e-09 0.0005 5.733e-09 0 5.927e-09 0 5.93e-09 0.0005 5.933e-09 0 6.127e-09 0 6.13e-09 0.0005 6.133e-09 0 6.327e-09 0 6.33e-09 0.0005 6.333e-09 0 7.327e-09 0 7.33e-09 0.0005 7.333e-09 0 7.527e-09 0 7.53e-09 0.0005 7.533e-09 0 7.727e-09 0 7.73e-09 0.0005 7.733e-09 0)
IDATA_B1|D 0 B1I  PWL(0 0 1.767e-09 0 1.77e-09 0.0005 1.773e-09 0 1.967e-09 0 1.97e-09 0.0005 1.973e-09 0 2.167e-09 0 2.17e-09 0.0005 2.173e-09 0 2.367e-09 0 2.37e-09 0.0005 2.373e-09 0 2.567e-09 0 2.57e-09 0.0005 2.573e-09 0 2.767e-09 0 2.77e-09 0.0005 2.773e-09 0 2.967e-09 0 2.97e-09 0.0005 2.973e-09 0 3.167e-09 0 3.17e-09 0.0005 3.173e-09 0 4.967e-09 0 4.97e-09 0.0005 4.973e-09 0 5.167e-09 0 5.17e-09 0.0005 5.173e-09 0 5.367e-09 0 5.37e-09 0.0005 5.373e-09 0 5.567e-09 0 5.57e-09 0.0005 5.573e-09 0 5.767e-09 0 5.77e-09 0.0005 5.773e-09 0 5.967e-09 0 5.97e-09 0.0005 5.973e-09 0 6.167e-09 0 6.17e-09 0.0005 6.173e-09 0 6.367e-09 0 6.37e-09 0.0005 6.373e-09 0)
L_SPL_P0_0|1 P0_0 _SPL_P0_0|D1  2e-12
L_SPL_P0_0|2 _SPL_P0_0|D1 _SPL_P0_0|D2  4.135667696e-12
L_SPL_P0_0|3 _SPL_P0_0|D2 _SPL_P0_0|JCT  1.4770241771428573e-12
L_SPL_P0_0|4 _SPL_P0_0|JCT _SPL_P0_0|QA1  1.4770241771428573e-12
L_SPL_P0_0|5 _SPL_P0_0|QA1 P0_0_B  2e-12
L_SPL_P0_0|6 _SPL_P0_0|JCT _SPL_P0_0|QB1  1.4770241771428573e-12
L_SPL_P0_0|7 _SPL_P0_0|QB1 P0_0_W  2e-12
L_SPL_G0_0|1 G0_0 _SPL_G0_0|D1  2e-12
L_SPL_G0_0|2 _SPL_G0_0|D1 _SPL_G0_0|D2  4.135667696e-12
L_SPL_G0_0|3 _SPL_G0_0|D2 _SPL_G0_0|JCT  1.4770241771428573e-12
L_SPL_G0_0|4 _SPL_G0_0|JCT _SPL_G0_0|QA1  1.4770241771428573e-12
L_SPL_G0_0|5 _SPL_G0_0|QA1 G0_0_B  2e-12
L_SPL_G0_0|6 _SPL_G0_0|JCT _SPL_G0_0|QB1  1.4770241771428573e-12
L_SPL_G0_0|7 _SPL_G0_0|QB1 G0_0_W  2e-12
L_SPL_P1_0|1 P1_0 _SPL_P1_0|D1  2e-12
L_SPL_P1_0|2 _SPL_P1_0|D1 _SPL_P1_0|D2  4.135667696e-12
L_SPL_P1_0|3 _SPL_P1_0|D2 _SPL_P1_0|JCT  1.4770241771428573e-12
L_SPL_P1_0|4 _SPL_P1_0|JCT _SPL_P1_0|QA1  1.4770241771428573e-12
L_SPL_P1_0|5 _SPL_P1_0|QA1 P1_0_B  2e-12
L_SPL_P1_0|6 _SPL_P1_0|JCT _SPL_P1_0|QB1  1.4770241771428573e-12
L_SPL_P1_0|7 _SPL_P1_0|QB1 P1_0_W  2e-12
L_DFF_P0_01|1 P0_0_W _DFF_P0_01|1  2.067833848e-12
L_DFF_P0_01|2 _DFF_P0_01|1 _DFF_P0_01|2  4.135667696e-12
L_DFF_P0_01|3 _DFF_P0_01|3 _DFF_P0_01|4  8.271335392e-12
L_DFF_P0_01|4 _DFF_P0_01|5 _DFF_P0_01|T1  4.135667696e-12
L_DFF_P0_01|T CLK1 _DFF_P0_01|T1  2.067833848e-12
L_DFF_P0_01|5 _DFF_P0_01|4 _DFF_P0_01|6  4.135667696e-12
L_DFF_P0_01|6 _DFF_P0_01|6 P0_1  2.067833848e-12
L_DFF_G0_01|1 G0_0_W _DFF_G0_01|1  2.067833848e-12
L_DFF_G0_01|2 _DFF_G0_01|1 _DFF_G0_01|2  4.135667696e-12
L_DFF_G0_01|3 _DFF_G0_01|3 _DFF_G0_01|4  8.271335392e-12
L_DFF_G0_01|4 _DFF_G0_01|5 _DFF_G0_01|T1  4.135667696e-12
L_DFF_G0_01|T CLK1 _DFF_G0_01|T1  2.067833848e-12
L_DFF_G0_01|5 _DFF_G0_01|4 _DFF_G0_01|6  4.135667696e-12
L_DFF_G0_01|6 _DFF_G0_01|6 G0_1  2.067833848e-12
L_DFF_P1_01|1 P1_0_W _DFF_P1_01|1  2.067833848e-12
L_DFF_P1_01|2 _DFF_P1_01|1 _DFF_P1_01|2  4.135667696e-12
L_DFF_P1_01|3 _DFF_P1_01|3 _DFF_P1_01|4  8.271335392e-12
L_DFF_P1_01|4 _DFF_P1_01|5 _DFF_P1_01|T1  4.135667696e-12
L_DFF_P1_01|T CLK1 _DFF_P1_01|T1  2.067833848e-12
L_DFF_P1_01|5 _DFF_P1_01|4 _DFF_P1_01|6  4.135667696e-12
L_DFF_P1_01|6 _DFF_P1_01|6 P1_1  2.067833848e-12
L_DFF_S0|1 P0_1 _DFF_S0|1  2.067833848e-12
L_DFF_S0|2 _DFF_S0|1 _DFF_S0|2  4.135667696e-12
L_DFF_S0|3 _DFF_S0|3 _DFF_S0|4  8.271335392e-12
L_DFF_S0|4 _DFF_S0|5 _DFF_S0|T1  4.135667696e-12
L_DFF_S0|T CLK2 _DFF_S0|T1  2.067833848e-12
L_DFF_S0|5 _DFF_S0|4 _DFF_S0|6  4.135667696e-12
L_DFF_S0|6 _DFF_S0|6 S0  2.067833848e-12
L_XOR_S1|A1 G0_1 _XOR_S1|A1  2.067833848e-12
L_XOR_S1|A2 _XOR_S1|A1 _XOR_S1|A2  4.135667696e-12
L_XOR_S1|A3 _XOR_S1|A3 _XOR_S1|AB  8.271335392e-12
L_XOR_S1|B1 P1_1 _XOR_S1|B1  2.067833848e-12
L_XOR_S1|B2 _XOR_S1|B1 _XOR_S1|B2  4.135667696e-12
L_XOR_S1|B3 _XOR_S1|B3 _XOR_S1|AB  8.271335392e-12
L_XOR_S1|T1 CLK2 _XOR_S1|T1  2.067833848e-12
L_XOR_S1|T2 _XOR_S1|T1 _XOR_S1|T2  4.135667696e-12
L_XOR_S1|Q2 _XOR_S1|ABTQ _XOR_S1|Q1  4.135667696e-12
L_XOR_S1|Q1 _XOR_S1|Q1 S1  2.067833848e-12
L_DFF_S2|1 G1_1 _DFF_S2|1  2.067833848e-12
L_DFF_S2|2 _DFF_S2|1 _DFF_S2|2  4.135667696e-12
L_DFF_S2|3 _DFF_S2|3 _DFF_S2|4  8.271335392e-12
L_DFF_S2|4 _DFF_S2|5 _DFF_S2|T1  4.135667696e-12
L_DFF_S2|T CLK2 _DFF_S2|T1  2.067833848e-12
L_DFF_S2|5 _DFF_S2|4 _DFF_S2|6  4.135667696e-12
L_DFF_S2|6 _DFF_S2|6 S2  2.067833848e-12
L_INIT_0|_SPL_A|1 A0I _INIT_0|_SPL_A|D1  2e-12
L_INIT_0|_SPL_A|2 _INIT_0|_SPL_A|D1 _INIT_0|_SPL_A|D2  4.135667696e-12
L_INIT_0|_SPL_A|3 _INIT_0|_SPL_A|D2 _INIT_0|_SPL_A|JCT  1.4770241771428573e-12
L_INIT_0|_SPL_A|4 _INIT_0|_SPL_A|JCT _INIT_0|_SPL_A|QA1  1.4770241771428573e-12
L_INIT_0|_SPL_A|5 _INIT_0|_SPL_A|QA1 _INIT_0|A1  2e-12
L_INIT_0|_SPL_A|6 _INIT_0|_SPL_A|JCT _INIT_0|_SPL_A|QB1  1.4770241771428573e-12
L_INIT_0|_SPL_A|7 _INIT_0|_SPL_A|QB1 _INIT_0|A2  2e-12
L_INIT_0|_SPL_B|1 B0I _INIT_0|_SPL_B|D1  2e-12
L_INIT_0|_SPL_B|2 _INIT_0|_SPL_B|D1 _INIT_0|_SPL_B|D2  4.135667696e-12
L_INIT_0|_SPL_B|3 _INIT_0|_SPL_B|D2 _INIT_0|_SPL_B|JCT  1.4770241771428573e-12
L_INIT_0|_SPL_B|4 _INIT_0|_SPL_B|JCT _INIT_0|_SPL_B|QA1  1.4770241771428573e-12
L_INIT_0|_SPL_B|5 _INIT_0|_SPL_B|QA1 _INIT_0|B1  2e-12
L_INIT_0|_SPL_B|6 _INIT_0|_SPL_B|JCT _INIT_0|_SPL_B|QB1  1.4770241771428573e-12
L_INIT_0|_SPL_B|7 _INIT_0|_SPL_B|QB1 _INIT_0|B2  2e-12
L_INIT_0|_DFF_A|1 _INIT_0|A1 _INIT_0|_DFF_A|1  2.067833848e-12
L_INIT_0|_DFF_A|2 _INIT_0|_DFF_A|1 _INIT_0|_DFF_A|2  4.135667696e-12
L_INIT_0|_DFF_A|3 _INIT_0|_DFF_A|3 _INIT_0|_DFF_A|4  8.271335392e-12
L_INIT_0|_DFF_A|4 _INIT_0|_DFF_A|5 _INIT_0|_DFF_A|T1  4.135667696e-12
L_INIT_0|_DFF_A|T CLK0 _INIT_0|_DFF_A|T1  2.067833848e-12
L_INIT_0|_DFF_A|5 _INIT_0|_DFF_A|4 _INIT_0|_DFF_A|6  4.135667696e-12
L_INIT_0|_DFF_A|6 _INIT_0|_DFF_A|6 _INIT_0|A1_SYNC  2.067833848e-12
L_INIT_0|_DFF_B|1 _INIT_0|B1 _INIT_0|_DFF_B|1  2.067833848e-12
L_INIT_0|_DFF_B|2 _INIT_0|_DFF_B|1 _INIT_0|_DFF_B|2  4.135667696e-12
L_INIT_0|_DFF_B|3 _INIT_0|_DFF_B|3 _INIT_0|_DFF_B|4  8.271335392e-12
L_INIT_0|_DFF_B|4 _INIT_0|_DFF_B|5 _INIT_0|_DFF_B|T1  4.135667696e-12
L_INIT_0|_DFF_B|T CLK0 _INIT_0|_DFF_B|T1  2.067833848e-12
L_INIT_0|_DFF_B|5 _INIT_0|_DFF_B|4 _INIT_0|_DFF_B|6  4.135667696e-12
L_INIT_0|_DFF_B|6 _INIT_0|_DFF_B|6 _INIT_0|B1_SYNC  2.067833848e-12
L_INIT_0|_XOR|A1 _INIT_0|A2 _INIT_0|_XOR|A1  2.067833848e-12
L_INIT_0|_XOR|A2 _INIT_0|_XOR|A1 _INIT_0|_XOR|A2  4.135667696e-12
L_INIT_0|_XOR|A3 _INIT_0|_XOR|A3 _INIT_0|_XOR|AB  8.271335392e-12
L_INIT_0|_XOR|B1 _INIT_0|B2 _INIT_0|_XOR|B1  2.067833848e-12
L_INIT_0|_XOR|B2 _INIT_0|_XOR|B1 _INIT_0|_XOR|B2  4.135667696e-12
L_INIT_0|_XOR|B3 _INIT_0|_XOR|B3 _INIT_0|_XOR|AB  8.271335392e-12
L_INIT_0|_XOR|T1 CLK0 _INIT_0|_XOR|T1  2.067833848e-12
L_INIT_0|_XOR|T2 _INIT_0|_XOR|T1 _INIT_0|_XOR|T2  4.135667696e-12
L_INIT_0|_XOR|Q2 _INIT_0|_XOR|ABTQ _INIT_0|_XOR|Q1  4.135667696e-12
L_INIT_0|_XOR|Q1 _INIT_0|_XOR|Q1 P0_0  2.067833848e-12
L_INIT_0|_AND|A1 _INIT_0|A1_SYNC _INIT_0|_AND|A1  2.067833848e-12
L_INIT_0|_AND|A2 _INIT_0|_AND|A1 _INIT_0|_AND|A2  4.135667696e-12
L_INIT_0|_AND|A3 _INIT_0|_AND|A3 _INIT_0|_AND|Q3  1.2e-12
L_INIT_0|_AND|B1 _INIT_0|B1_SYNC _INIT_0|_AND|B1  2.067833848e-12
L_INIT_0|_AND|B2 _INIT_0|_AND|B1 _INIT_0|_AND|B2  4.135667696e-12
L_INIT_0|_AND|B3 _INIT_0|_AND|B3 _INIT_0|_AND|Q3  1.2e-12
L_INIT_0|_AND|Q3 _INIT_0|_AND|Q3 _INIT_0|_AND|Q2  4.135667696e-12
L_INIT_0|_AND|Q2 _INIT_0|_AND|Q2 _INIT_0|_AND|Q1  4.135667696e-12
L_INIT_0|_AND|Q1 _INIT_0|_AND|Q1 G0_0  2.067833848e-12
L_INIT_1|_SPL_A|1 A1I _INIT_1|_SPL_A|D1  2e-12
L_INIT_1|_SPL_A|2 _INIT_1|_SPL_A|D1 _INIT_1|_SPL_A|D2  4.135667696e-12
L_INIT_1|_SPL_A|3 _INIT_1|_SPL_A|D2 _INIT_1|_SPL_A|JCT  1.4770241771428573e-12
L_INIT_1|_SPL_A|4 _INIT_1|_SPL_A|JCT _INIT_1|_SPL_A|QA1  1.4770241771428573e-12
L_INIT_1|_SPL_A|5 _INIT_1|_SPL_A|QA1 _INIT_1|A1  2e-12
L_INIT_1|_SPL_A|6 _INIT_1|_SPL_A|JCT _INIT_1|_SPL_A|QB1  1.4770241771428573e-12
L_INIT_1|_SPL_A|7 _INIT_1|_SPL_A|QB1 _INIT_1|A2  2e-12
L_INIT_1|_SPL_B|1 B1I _INIT_1|_SPL_B|D1  2e-12
L_INIT_1|_SPL_B|2 _INIT_1|_SPL_B|D1 _INIT_1|_SPL_B|D2  4.135667696e-12
L_INIT_1|_SPL_B|3 _INIT_1|_SPL_B|D2 _INIT_1|_SPL_B|JCT  1.4770241771428573e-12
L_INIT_1|_SPL_B|4 _INIT_1|_SPL_B|JCT _INIT_1|_SPL_B|QA1  1.4770241771428573e-12
L_INIT_1|_SPL_B|5 _INIT_1|_SPL_B|QA1 _INIT_1|B1  2e-12
L_INIT_1|_SPL_B|6 _INIT_1|_SPL_B|JCT _INIT_1|_SPL_B|QB1  1.4770241771428573e-12
L_INIT_1|_SPL_B|7 _INIT_1|_SPL_B|QB1 _INIT_1|B2  2e-12
L_INIT_1|_DFF_A|1 _INIT_1|A1 _INIT_1|_DFF_A|1  2.067833848e-12
L_INIT_1|_DFF_A|2 _INIT_1|_DFF_A|1 _INIT_1|_DFF_A|2  4.135667696e-12
L_INIT_1|_DFF_A|3 _INIT_1|_DFF_A|3 _INIT_1|_DFF_A|4  8.271335392e-12
L_INIT_1|_DFF_A|4 _INIT_1|_DFF_A|5 _INIT_1|_DFF_A|T1  4.135667696e-12
L_INIT_1|_DFF_A|T CLK0 _INIT_1|_DFF_A|T1  2.067833848e-12
L_INIT_1|_DFF_A|5 _INIT_1|_DFF_A|4 _INIT_1|_DFF_A|6  4.135667696e-12
L_INIT_1|_DFF_A|6 _INIT_1|_DFF_A|6 _INIT_1|A1_SYNC  2.067833848e-12
L_INIT_1|_DFF_B|1 _INIT_1|B1 _INIT_1|_DFF_B|1  2.067833848e-12
L_INIT_1|_DFF_B|2 _INIT_1|_DFF_B|1 _INIT_1|_DFF_B|2  4.135667696e-12
L_INIT_1|_DFF_B|3 _INIT_1|_DFF_B|3 _INIT_1|_DFF_B|4  8.271335392e-12
L_INIT_1|_DFF_B|4 _INIT_1|_DFF_B|5 _INIT_1|_DFF_B|T1  4.135667696e-12
L_INIT_1|_DFF_B|T CLK0 _INIT_1|_DFF_B|T1  2.067833848e-12
L_INIT_1|_DFF_B|5 _INIT_1|_DFF_B|4 _INIT_1|_DFF_B|6  4.135667696e-12
L_INIT_1|_DFF_B|6 _INIT_1|_DFF_B|6 _INIT_1|B1_SYNC  2.067833848e-12
L_INIT_1|_XOR|A1 _INIT_1|A2 _INIT_1|_XOR|A1  2.067833848e-12
L_INIT_1|_XOR|A2 _INIT_1|_XOR|A1 _INIT_1|_XOR|A2  4.135667696e-12
L_INIT_1|_XOR|A3 _INIT_1|_XOR|A3 _INIT_1|_XOR|AB  8.271335392e-12
L_INIT_1|_XOR|B1 _INIT_1|B2 _INIT_1|_XOR|B1  2.067833848e-12
L_INIT_1|_XOR|B2 _INIT_1|_XOR|B1 _INIT_1|_XOR|B2  4.135667696e-12
L_INIT_1|_XOR|B3 _INIT_1|_XOR|B3 _INIT_1|_XOR|AB  8.271335392e-12
L_INIT_1|_XOR|T1 CLK0 _INIT_1|_XOR|T1  2.067833848e-12
L_INIT_1|_XOR|T2 _INIT_1|_XOR|T1 _INIT_1|_XOR|T2  4.135667696e-12
L_INIT_1|_XOR|Q2 _INIT_1|_XOR|ABTQ _INIT_1|_XOR|Q1  4.135667696e-12
L_INIT_1|_XOR|Q1 _INIT_1|_XOR|Q1 P1_0  2.067833848e-12
L_INIT_1|_AND|A1 _INIT_1|A1_SYNC _INIT_1|_AND|A1  2.067833848e-12
L_INIT_1|_AND|A2 _INIT_1|_AND|A1 _INIT_1|_AND|A2  4.135667696e-12
L_INIT_1|_AND|A3 _INIT_1|_AND|A3 _INIT_1|_AND|Q3  1.2e-12
L_INIT_1|_AND|B1 _INIT_1|B1_SYNC _INIT_1|_AND|B1  2.067833848e-12
L_INIT_1|_AND|B2 _INIT_1|_AND|B1 _INIT_1|_AND|B2  4.135667696e-12
L_INIT_1|_AND|B3 _INIT_1|_AND|B3 _INIT_1|_AND|Q3  1.2e-12
L_INIT_1|_AND|Q3 _INIT_1|_AND|Q3 _INIT_1|_AND|Q2  4.135667696e-12
L_INIT_1|_AND|Q2 _INIT_1|_AND|Q2 _INIT_1|_AND|Q1  4.135667696e-12
L_INIT_1|_AND|Q1 _INIT_1|_AND|Q1 G1_0  2.067833848e-12
L_SPL_P0_0|I_D1|B _SPL_P0_0|D1 _SPL_P0_0|I_D1|MID  2e-12
I_SPL_P0_0|I_D1|B 0 _SPL_P0_0|I_D1|MID  0.000175
L_SPL_P0_0|I_D2|B _SPL_P0_0|D2 _SPL_P0_0|I_D2|MID  2e-12
I_SPL_P0_0|I_D2|B 0 _SPL_P0_0|I_D2|MID  0.000245
L_SPL_P0_0|I_Q1|B _SPL_P0_0|QA1 _SPL_P0_0|I_Q1|MID  2e-12
I_SPL_P0_0|I_Q1|B 0 _SPL_P0_0|I_Q1|MID  0.000175
L_SPL_P0_0|I_Q2|B _SPL_P0_0|QB1 _SPL_P0_0|I_Q2|MID  2e-12
I_SPL_P0_0|I_Q2|B 0 _SPL_P0_0|I_Q2|MID  0.000175
B_SPL_P0_0|1|1 _SPL_P0_0|D1 _SPL_P0_0|1|MID_SERIES JJMIT AREA=2.5
L_SPL_P0_0|1|P _SPL_P0_0|1|MID_SERIES 0  2e-13
R_SPL_P0_0|1|B _SPL_P0_0|D1 _SPL_P0_0|1|MID_SHUNT  2.7439617672
L_SPL_P0_0|1|RB _SPL_P0_0|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_P0_0|2|1 _SPL_P0_0|D2 _SPL_P0_0|2|MID_SERIES JJMIT AREA=2.5
L_SPL_P0_0|2|P _SPL_P0_0|2|MID_SERIES 0  2e-13
R_SPL_P0_0|2|B _SPL_P0_0|D2 _SPL_P0_0|2|MID_SHUNT  2.7439617672
L_SPL_P0_0|2|RB _SPL_P0_0|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_P0_0|A|1 _SPL_P0_0|QA1 _SPL_P0_0|A|MID_SERIES JJMIT AREA=2.5
L_SPL_P0_0|A|P _SPL_P0_0|A|MID_SERIES 0  2e-13
R_SPL_P0_0|A|B _SPL_P0_0|QA1 _SPL_P0_0|A|MID_SHUNT  2.7439617672
L_SPL_P0_0|A|RB _SPL_P0_0|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_P0_0|B|1 _SPL_P0_0|QB1 _SPL_P0_0|B|MID_SERIES JJMIT AREA=2.5
L_SPL_P0_0|B|P _SPL_P0_0|B|MID_SERIES 0  2e-13
R_SPL_P0_0|B|B _SPL_P0_0|QB1 _SPL_P0_0|B|MID_SHUNT  2.7439617672
L_SPL_P0_0|B|RB _SPL_P0_0|B|MID_SHUNT 0  1.550338398468e-12
L_SPL_G0_0|I_D1|B _SPL_G0_0|D1 _SPL_G0_0|I_D1|MID  2e-12
I_SPL_G0_0|I_D1|B 0 _SPL_G0_0|I_D1|MID  0.000175
L_SPL_G0_0|I_D2|B _SPL_G0_0|D2 _SPL_G0_0|I_D2|MID  2e-12
I_SPL_G0_0|I_D2|B 0 _SPL_G0_0|I_D2|MID  0.000245
L_SPL_G0_0|I_Q1|B _SPL_G0_0|QA1 _SPL_G0_0|I_Q1|MID  2e-12
I_SPL_G0_0|I_Q1|B 0 _SPL_G0_0|I_Q1|MID  0.000175
L_SPL_G0_0|I_Q2|B _SPL_G0_0|QB1 _SPL_G0_0|I_Q2|MID  2e-12
I_SPL_G0_0|I_Q2|B 0 _SPL_G0_0|I_Q2|MID  0.000175
B_SPL_G0_0|1|1 _SPL_G0_0|D1 _SPL_G0_0|1|MID_SERIES JJMIT AREA=2.5
L_SPL_G0_0|1|P _SPL_G0_0|1|MID_SERIES 0  2e-13
R_SPL_G0_0|1|B _SPL_G0_0|D1 _SPL_G0_0|1|MID_SHUNT  2.7439617672
L_SPL_G0_0|1|RB _SPL_G0_0|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_G0_0|2|1 _SPL_G0_0|D2 _SPL_G0_0|2|MID_SERIES JJMIT AREA=2.5
L_SPL_G0_0|2|P _SPL_G0_0|2|MID_SERIES 0  2e-13
R_SPL_G0_0|2|B _SPL_G0_0|D2 _SPL_G0_0|2|MID_SHUNT  2.7439617672
L_SPL_G0_0|2|RB _SPL_G0_0|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_G0_0|A|1 _SPL_G0_0|QA1 _SPL_G0_0|A|MID_SERIES JJMIT AREA=2.5
L_SPL_G0_0|A|P _SPL_G0_0|A|MID_SERIES 0  2e-13
R_SPL_G0_0|A|B _SPL_G0_0|QA1 _SPL_G0_0|A|MID_SHUNT  2.7439617672
L_SPL_G0_0|A|RB _SPL_G0_0|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_G0_0|B|1 _SPL_G0_0|QB1 _SPL_G0_0|B|MID_SERIES JJMIT AREA=2.5
L_SPL_G0_0|B|P _SPL_G0_0|B|MID_SERIES 0  2e-13
R_SPL_G0_0|B|B _SPL_G0_0|QB1 _SPL_G0_0|B|MID_SHUNT  2.7439617672
L_SPL_G0_0|B|RB _SPL_G0_0|B|MID_SHUNT 0  1.550338398468e-12
L_SPL_P1_0|I_D1|B _SPL_P1_0|D1 _SPL_P1_0|I_D1|MID  2e-12
I_SPL_P1_0|I_D1|B 0 _SPL_P1_0|I_D1|MID  0.000175
L_SPL_P1_0|I_D2|B _SPL_P1_0|D2 _SPL_P1_0|I_D2|MID  2e-12
I_SPL_P1_0|I_D2|B 0 _SPL_P1_0|I_D2|MID  0.000245
L_SPL_P1_0|I_Q1|B _SPL_P1_0|QA1 _SPL_P1_0|I_Q1|MID  2e-12
I_SPL_P1_0|I_Q1|B 0 _SPL_P1_0|I_Q1|MID  0.000175
L_SPL_P1_0|I_Q2|B _SPL_P1_0|QB1 _SPL_P1_0|I_Q2|MID  2e-12
I_SPL_P1_0|I_Q2|B 0 _SPL_P1_0|I_Q2|MID  0.000175
B_SPL_P1_0|1|1 _SPL_P1_0|D1 _SPL_P1_0|1|MID_SERIES JJMIT AREA=2.5
L_SPL_P1_0|1|P _SPL_P1_0|1|MID_SERIES 0  2e-13
R_SPL_P1_0|1|B _SPL_P1_0|D1 _SPL_P1_0|1|MID_SHUNT  2.7439617672
L_SPL_P1_0|1|RB _SPL_P1_0|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_P1_0|2|1 _SPL_P1_0|D2 _SPL_P1_0|2|MID_SERIES JJMIT AREA=2.5
L_SPL_P1_0|2|P _SPL_P1_0|2|MID_SERIES 0  2e-13
R_SPL_P1_0|2|B _SPL_P1_0|D2 _SPL_P1_0|2|MID_SHUNT  2.7439617672
L_SPL_P1_0|2|RB _SPL_P1_0|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_P1_0|A|1 _SPL_P1_0|QA1 _SPL_P1_0|A|MID_SERIES JJMIT AREA=2.5
L_SPL_P1_0|A|P _SPL_P1_0|A|MID_SERIES 0  2e-13
R_SPL_P1_0|A|B _SPL_P1_0|QA1 _SPL_P1_0|A|MID_SHUNT  2.7439617672
L_SPL_P1_0|A|RB _SPL_P1_0|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_P1_0|B|1 _SPL_P1_0|QB1 _SPL_P1_0|B|MID_SERIES JJMIT AREA=2.5
L_SPL_P1_0|B|P _SPL_P1_0|B|MID_SERIES 0  2e-13
R_SPL_P1_0|B|B _SPL_P1_0|QB1 _SPL_P1_0|B|MID_SHUNT  2.7439617672
L_SPL_P1_0|B|RB _SPL_P1_0|B|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_SPL_G1|1 G1_0 _PG_01|_SPL_G1|D1  2e-12
L_PG_01|_SPL_G1|2 _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|D2  4.135667696e-12
L_PG_01|_SPL_G1|3 _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|JCT  1.4770241771428573e-12
L_PG_01|_SPL_G1|4 _PG_01|_SPL_G1|JCT _PG_01|_SPL_G1|QA1  1.4770241771428573e-12
L_PG_01|_SPL_G1|5 _PG_01|_SPL_G1|QA1 _PG_01|G1_COPY_1  2e-12
L_PG_01|_SPL_G1|6 _PG_01|_SPL_G1|JCT _PG_01|_SPL_G1|QB1  1.4770241771428573e-12
L_PG_01|_SPL_G1|7 _PG_01|_SPL_G1|QB1 _PG_01|G1_COPY_2  2e-12
L_PG_01|_SPL_P1|1 P1_0_B _PG_01|_SPL_P1|D1  2e-12
L_PG_01|_SPL_P1|2 _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|D2  4.135667696e-12
L_PG_01|_SPL_P1|3 _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|JCT  1.4770241771428573e-12
L_PG_01|_SPL_P1|4 _PG_01|_SPL_P1|JCT _PG_01|_SPL_P1|QA1  1.4770241771428573e-12
L_PG_01|_SPL_P1|5 _PG_01|_SPL_P1|QA1 _PG_01|P1_COPY_1  2e-12
L_PG_01|_SPL_P1|6 _PG_01|_SPL_P1|JCT _PG_01|_SPL_P1|QB1  1.4770241771428573e-12
L_PG_01|_SPL_P1|7 _PG_01|_SPL_P1|QB1 _PG_01|P1_COPY_2  2e-12
L_PG_01|_PG|A1 _PG_01|P1_COPY_1 _PG_01|_PG|A1  2.067833848e-12
L_PG_01|_PG|A2 _PG_01|_PG|A1 _PG_01|_PG|A2  4.135667696e-12
L_PG_01|_PG|A3 _PG_01|_PG|A3 _PG_01|_PG|Q3  1.2e-12
L_PG_01|_PG|B1 _PG_01|G1_COPY_1 _PG_01|_PG|B1  2.067833848e-12
L_PG_01|_PG|B2 _PG_01|_PG|B1 _PG_01|_PG|B2  4.135667696e-12
L_PG_01|_PG|B3 _PG_01|_PG|B3 _PG_01|_PG|Q3  1.2e-12
L_PG_01|_PG|Q3 _PG_01|_PG|Q3 _PG_01|_PG|Q2  4.135667696e-12
L_PG_01|_PG|Q2 _PG_01|_PG|Q2 _PG_01|_PG|Q1  4.135667696e-12
L_PG_01|_PG|Q1 _PG_01|_PG|Q1 _PG_01|PG  2.067833848e-12
L_PG_01|_GG|A1 G0_0_B _PG_01|_GG|A1  2.067833848e-12
L_PG_01|_GG|A2 _PG_01|_GG|A1 _PG_01|_GG|A2  4.135667696e-12
L_PG_01|_GG|A3 _PG_01|_GG|A3 _PG_01|_GG|Q3  1.2e-12
L_PG_01|_GG|B1 _PG_01|G1_COPY_2 _PG_01|_GG|B1  2.067833848e-12
L_PG_01|_GG|B2 _PG_01|_GG|B1 _PG_01|_GG|B2  4.135667696e-12
L_PG_01|_GG|B3 _PG_01|_GG|B3 _PG_01|_GG|Q3  1.2e-12
L_PG_01|_GG|Q3 _PG_01|_GG|Q3 _PG_01|_GG|Q2  4.135667696e-12
L_PG_01|_GG|Q2 _PG_01|_GG|Q2 _PG_01|_GG|Q1  4.135667696e-12
L_PG_01|_GG|Q1 _PG_01|_GG|Q1 _PG_01|GG  2.067833848e-12
L_PG_01|_DFF_P0|1 P0_0_B _PG_01|_DFF_P0|1  2.067833848e-12
L_PG_01|_DFF_P0|2 _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|2  4.135667696e-12
L_PG_01|_DFF_P0|3 _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|4  8.271335392e-12
L_PG_01|_DFF_P0|4 _PG_01|_DFF_P0|5 _PG_01|_DFF_P0|T1  4.135667696e-12
L_PG_01|_DFF_P0|T CLK1 _PG_01|_DFF_P0|T1  2.067833848e-12
L_PG_01|_DFF_P0|5 _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|6  4.135667696e-12
L_PG_01|_DFF_P0|6 _PG_01|_DFF_P0|6 _PG_01|P0_SYNC  2.067833848e-12
L_PG_01|_DFF_P1|1 _PG_01|P1_COPY_2 _PG_01|_DFF_P1|1  2.067833848e-12
L_PG_01|_DFF_P1|2 _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|2  4.135667696e-12
L_PG_01|_DFF_P1|3 _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|4  8.271335392e-12
L_PG_01|_DFF_P1|4 _PG_01|_DFF_P1|5 _PG_01|_DFF_P1|T1  4.135667696e-12
L_PG_01|_DFF_P1|T CLK1 _PG_01|_DFF_P1|T1  2.067833848e-12
L_PG_01|_DFF_P1|5 _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|6  4.135667696e-12
L_PG_01|_DFF_P1|6 _PG_01|_DFF_P1|6 _PG_01|P1_SYNC  2.067833848e-12
L_PG_01|_DFF_PG|1 _PG_01|PG _PG_01|_DFF_PG|1  2.067833848e-12
L_PG_01|_DFF_PG|2 _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|2  4.135667696e-12
L_PG_01|_DFF_PG|3 _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|4  8.271335392e-12
L_PG_01|_DFF_PG|4 _PG_01|_DFF_PG|5 _PG_01|_DFF_PG|T1  4.135667696e-12
L_PG_01|_DFF_PG|T CLK1 _PG_01|_DFF_PG|T1  2.067833848e-12
L_PG_01|_DFF_PG|5 _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|6  4.135667696e-12
L_PG_01|_DFF_PG|6 _PG_01|_DFF_PG|6 _PG_01|PG_SYNC  2.067833848e-12
L_PG_01|_DFF_GG|1 _PG_01|GG _PG_01|_DFF_GG|1  2.067833848e-12
L_PG_01|_DFF_GG|2 _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|2  4.135667696e-12
L_PG_01|_DFF_GG|3 _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|4  8.271335392e-12
L_PG_01|_DFF_GG|4 _PG_01|_DFF_GG|5 _PG_01|_DFF_GG|T1  4.135667696e-12
L_PG_01|_DFF_GG|T CLK1 _PG_01|_DFF_GG|T1  2.067833848e-12
L_PG_01|_DFF_GG|5 _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|6  4.135667696e-12
L_PG_01|_DFF_GG|6 _PG_01|_DFF_GG|6 _PG_01|GG_SYNC  2.067833848e-12
L_PG_01|_AND_G|A1 _PG_01|PG_SYNC _PG_01|_AND_G|A1  2.067833848e-12
L_PG_01|_AND_G|A2 _PG_01|_AND_G|A1 _PG_01|_AND_G|A2  4.135667696e-12
L_PG_01|_AND_G|A3 _PG_01|_AND_G|A3 _PG_01|_AND_G|Q3  1.2e-12
L_PG_01|_AND_G|B1 _PG_01|GG_SYNC _PG_01|_AND_G|B1  2.067833848e-12
L_PG_01|_AND_G|B2 _PG_01|_AND_G|B1 _PG_01|_AND_G|B2  4.135667696e-12
L_PG_01|_AND_G|B3 _PG_01|_AND_G|B3 _PG_01|_AND_G|Q3  1.2e-12
L_PG_01|_AND_G|Q3 _PG_01|_AND_G|Q3 _PG_01|_AND_G|Q2  4.135667696e-12
L_PG_01|_AND_G|Q2 _PG_01|_AND_G|Q2 _PG_01|_AND_G|Q1  4.135667696e-12
L_PG_01|_AND_G|Q1 _PG_01|_AND_G|Q1 G1_1  2.067833848e-12
L_PG_01|_AND_P|A1 _PG_01|P0_SYNC _PG_01|_AND_P|A1  2.067833848e-12
L_PG_01|_AND_P|A2 _PG_01|_AND_P|A1 _PG_01|_AND_P|A2  4.135667696e-12
L_PG_01|_AND_P|A3 _PG_01|_AND_P|A3 _PG_01|_AND_P|Q3  1.2e-12
L_PG_01|_AND_P|B1 _PG_01|P1_SYNC _PG_01|_AND_P|B1  2.067833848e-12
L_PG_01|_AND_P|B2 _PG_01|_AND_P|B1 _PG_01|_AND_P|B2  4.135667696e-12
L_PG_01|_AND_P|B3 _PG_01|_AND_P|B3 _PG_01|_AND_P|Q3  1.2e-12
L_PG_01|_AND_P|Q3 _PG_01|_AND_P|Q3 _PG_01|_AND_P|Q2  4.135667696e-12
L_PG_01|_AND_P|Q2 _PG_01|_AND_P|Q2 _PG_01|_AND_P|Q1  4.135667696e-12
L_PG_01|_AND_P|Q1 _PG_01|_AND_P|Q1 P1_1  2.067833848e-12
B_DFF_P0_01|1|1 _DFF_P0_01|1 _DFF_P0_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_P0_01|1|P _DFF_P0_01|1|MID_SERIES 0  2e-13
R_DFF_P0_01|1|B _DFF_P0_01|1 _DFF_P0_01|1|MID_SHUNT  2.7439617672
L_DFF_P0_01|1|RB _DFF_P0_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_P0_01|23|1 _DFF_P0_01|2 _DFF_P0_01|3 JJMIT AREA=1.7857142857142858
R_DFF_P0_01|23|B _DFF_P0_01|2 _DFF_P0_01|23|MID_SHUNT  3.84154647408
L_DFF_P0_01|23|RB _DFF_P0_01|23|MID_SHUNT _DFF_P0_01|3  2.1704737578552e-12
B_DFF_P0_01|3|1 _DFF_P0_01|3 _DFF_P0_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_P0_01|3|P _DFF_P0_01|3|MID_SERIES 0  2e-13
R_DFF_P0_01|3|B _DFF_P0_01|3 _DFF_P0_01|3|MID_SHUNT  2.7439617672
L_DFF_P0_01|3|RB _DFF_P0_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_P0_01|4|1 _DFF_P0_01|4 _DFF_P0_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_P0_01|4|P _DFF_P0_01|4|MID_SERIES 0  2e-13
R_DFF_P0_01|4|B _DFF_P0_01|4 _DFF_P0_01|4|MID_SHUNT  2.7439617672
L_DFF_P0_01|4|RB _DFF_P0_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_P0_01|45|1 _DFF_P0_01|4 _DFF_P0_01|5 JJMIT AREA=1.7857142857142858
R_DFF_P0_01|45|B _DFF_P0_01|4 _DFF_P0_01|45|MID_SHUNT  3.84154647408
L_DFF_P0_01|45|RB _DFF_P0_01|45|MID_SHUNT _DFF_P0_01|5  2.1704737578552e-12
B_DFF_P0_01|T|1 _DFF_P0_01|T1 _DFF_P0_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_P0_01|T|P _DFF_P0_01|T|MID_SERIES 0  2e-13
R_DFF_P0_01|T|B _DFF_P0_01|T1 _DFF_P0_01|T|MID_SHUNT  2.7439617672
L_DFF_P0_01|T|RB _DFF_P0_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_P0_01|6|1 _DFF_P0_01|6 _DFF_P0_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_P0_01|6|P _DFF_P0_01|6|MID_SERIES 0  2e-13
R_DFF_P0_01|6|B _DFF_P0_01|6 _DFF_P0_01|6|MID_SHUNT  2.7439617672
L_DFF_P0_01|6|RB _DFF_P0_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_P0_01|I_1|B _DFF_P0_01|1 _DFF_P0_01|I_1|MID  2e-12
I_DFF_P0_01|I_1|B 0 _DFF_P0_01|I_1|MID  0.000175
L_DFF_P0_01|I_3|B _DFF_P0_01|3 _DFF_P0_01|I_3|MID  2e-12
I_DFF_P0_01|I_3|B 0 _DFF_P0_01|I_3|MID  0.00025
L_DFF_P0_01|I_T|B _DFF_P0_01|T1 _DFF_P0_01|I_T|MID  2e-12
I_DFF_P0_01|I_T|B 0 _DFF_P0_01|I_T|MID  0.000175
L_DFF_P0_01|I_6|B _DFF_P0_01|6 _DFF_P0_01|I_6|MID  2e-12
I_DFF_P0_01|I_6|B 0 _DFF_P0_01|I_6|MID  0.000175
B_DFF_G0_01|1|1 _DFF_G0_01|1 _DFF_G0_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_G0_01|1|P _DFF_G0_01|1|MID_SERIES 0  2e-13
R_DFF_G0_01|1|B _DFF_G0_01|1 _DFF_G0_01|1|MID_SHUNT  2.7439617672
L_DFF_G0_01|1|RB _DFF_G0_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_G0_01|23|1 _DFF_G0_01|2 _DFF_G0_01|3 JJMIT AREA=1.7857142857142858
R_DFF_G0_01|23|B _DFF_G0_01|2 _DFF_G0_01|23|MID_SHUNT  3.84154647408
L_DFF_G0_01|23|RB _DFF_G0_01|23|MID_SHUNT _DFF_G0_01|3  2.1704737578552e-12
B_DFF_G0_01|3|1 _DFF_G0_01|3 _DFF_G0_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_G0_01|3|P _DFF_G0_01|3|MID_SERIES 0  2e-13
R_DFF_G0_01|3|B _DFF_G0_01|3 _DFF_G0_01|3|MID_SHUNT  2.7439617672
L_DFF_G0_01|3|RB _DFF_G0_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_G0_01|4|1 _DFF_G0_01|4 _DFF_G0_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_G0_01|4|P _DFF_G0_01|4|MID_SERIES 0  2e-13
R_DFF_G0_01|4|B _DFF_G0_01|4 _DFF_G0_01|4|MID_SHUNT  2.7439617672
L_DFF_G0_01|4|RB _DFF_G0_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_G0_01|45|1 _DFF_G0_01|4 _DFF_G0_01|5 JJMIT AREA=1.7857142857142858
R_DFF_G0_01|45|B _DFF_G0_01|4 _DFF_G0_01|45|MID_SHUNT  3.84154647408
L_DFF_G0_01|45|RB _DFF_G0_01|45|MID_SHUNT _DFF_G0_01|5  2.1704737578552e-12
B_DFF_G0_01|T|1 _DFF_G0_01|T1 _DFF_G0_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_G0_01|T|P _DFF_G0_01|T|MID_SERIES 0  2e-13
R_DFF_G0_01|T|B _DFF_G0_01|T1 _DFF_G0_01|T|MID_SHUNT  2.7439617672
L_DFF_G0_01|T|RB _DFF_G0_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_G0_01|6|1 _DFF_G0_01|6 _DFF_G0_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_G0_01|6|P _DFF_G0_01|6|MID_SERIES 0  2e-13
R_DFF_G0_01|6|B _DFF_G0_01|6 _DFF_G0_01|6|MID_SHUNT  2.7439617672
L_DFF_G0_01|6|RB _DFF_G0_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_G0_01|I_1|B _DFF_G0_01|1 _DFF_G0_01|I_1|MID  2e-12
I_DFF_G0_01|I_1|B 0 _DFF_G0_01|I_1|MID  0.000175
L_DFF_G0_01|I_3|B _DFF_G0_01|3 _DFF_G0_01|I_3|MID  2e-12
I_DFF_G0_01|I_3|B 0 _DFF_G0_01|I_3|MID  0.00025
L_DFF_G0_01|I_T|B _DFF_G0_01|T1 _DFF_G0_01|I_T|MID  2e-12
I_DFF_G0_01|I_T|B 0 _DFF_G0_01|I_T|MID  0.000175
L_DFF_G0_01|I_6|B _DFF_G0_01|6 _DFF_G0_01|I_6|MID  2e-12
I_DFF_G0_01|I_6|B 0 _DFF_G0_01|I_6|MID  0.000175
B_DFF_P1_01|1|1 _DFF_P1_01|1 _DFF_P1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_P1_01|1|P _DFF_P1_01|1|MID_SERIES 0  2e-13
R_DFF_P1_01|1|B _DFF_P1_01|1 _DFF_P1_01|1|MID_SHUNT  2.7439617672
L_DFF_P1_01|1|RB _DFF_P1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_P1_01|23|1 _DFF_P1_01|2 _DFF_P1_01|3 JJMIT AREA=1.7857142857142858
R_DFF_P1_01|23|B _DFF_P1_01|2 _DFF_P1_01|23|MID_SHUNT  3.84154647408
L_DFF_P1_01|23|RB _DFF_P1_01|23|MID_SHUNT _DFF_P1_01|3  2.1704737578552e-12
B_DFF_P1_01|3|1 _DFF_P1_01|3 _DFF_P1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_P1_01|3|P _DFF_P1_01|3|MID_SERIES 0  2e-13
R_DFF_P1_01|3|B _DFF_P1_01|3 _DFF_P1_01|3|MID_SHUNT  2.7439617672
L_DFF_P1_01|3|RB _DFF_P1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_P1_01|4|1 _DFF_P1_01|4 _DFF_P1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_P1_01|4|P _DFF_P1_01|4|MID_SERIES 0  2e-13
R_DFF_P1_01|4|B _DFF_P1_01|4 _DFF_P1_01|4|MID_SHUNT  2.7439617672
L_DFF_P1_01|4|RB _DFF_P1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_P1_01|45|1 _DFF_P1_01|4 _DFF_P1_01|5 JJMIT AREA=1.7857142857142858
R_DFF_P1_01|45|B _DFF_P1_01|4 _DFF_P1_01|45|MID_SHUNT  3.84154647408
L_DFF_P1_01|45|RB _DFF_P1_01|45|MID_SHUNT _DFF_P1_01|5  2.1704737578552e-12
B_DFF_P1_01|T|1 _DFF_P1_01|T1 _DFF_P1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_P1_01|T|P _DFF_P1_01|T|MID_SERIES 0  2e-13
R_DFF_P1_01|T|B _DFF_P1_01|T1 _DFF_P1_01|T|MID_SHUNT  2.7439617672
L_DFF_P1_01|T|RB _DFF_P1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_P1_01|6|1 _DFF_P1_01|6 _DFF_P1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_P1_01|6|P _DFF_P1_01|6|MID_SERIES 0  2e-13
R_DFF_P1_01|6|B _DFF_P1_01|6 _DFF_P1_01|6|MID_SHUNT  2.7439617672
L_DFF_P1_01|6|RB _DFF_P1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_P1_01|I_1|B _DFF_P1_01|1 _DFF_P1_01|I_1|MID  2e-12
I_DFF_P1_01|I_1|B 0 _DFF_P1_01|I_1|MID  0.000175
L_DFF_P1_01|I_3|B _DFF_P1_01|3 _DFF_P1_01|I_3|MID  2e-12
I_DFF_P1_01|I_3|B 0 _DFF_P1_01|I_3|MID  0.00025
L_DFF_P1_01|I_T|B _DFF_P1_01|T1 _DFF_P1_01|I_T|MID  2e-12
I_DFF_P1_01|I_T|B 0 _DFF_P1_01|I_T|MID  0.000175
L_DFF_P1_01|I_6|B _DFF_P1_01|6 _DFF_P1_01|I_6|MID  2e-12
I_DFF_P1_01|I_6|B 0 _DFF_P1_01|I_6|MID  0.000175
B_DFF_S0|1|1 _DFF_S0|1 _DFF_S0|1|MID_SERIES JJMIT AREA=2.5
L_DFF_S0|1|P _DFF_S0|1|MID_SERIES 0  2e-13
R_DFF_S0|1|B _DFF_S0|1 _DFF_S0|1|MID_SHUNT  2.7439617672
L_DFF_S0|1|RB _DFF_S0|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_S0|23|1 _DFF_S0|2 _DFF_S0|3 JJMIT AREA=1.7857142857142858
R_DFF_S0|23|B _DFF_S0|2 _DFF_S0|23|MID_SHUNT  3.84154647408
L_DFF_S0|23|RB _DFF_S0|23|MID_SHUNT _DFF_S0|3  2.1704737578552e-12
B_DFF_S0|3|1 _DFF_S0|3 _DFF_S0|3|MID_SERIES JJMIT AREA=2.5
L_DFF_S0|3|P _DFF_S0|3|MID_SERIES 0  2e-13
R_DFF_S0|3|B _DFF_S0|3 _DFF_S0|3|MID_SHUNT  2.7439617672
L_DFF_S0|3|RB _DFF_S0|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_S0|4|1 _DFF_S0|4 _DFF_S0|4|MID_SERIES JJMIT AREA=2.5
L_DFF_S0|4|P _DFF_S0|4|MID_SERIES 0  2e-13
R_DFF_S0|4|B _DFF_S0|4 _DFF_S0|4|MID_SHUNT  2.7439617672
L_DFF_S0|4|RB _DFF_S0|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_S0|45|1 _DFF_S0|4 _DFF_S0|5 JJMIT AREA=1.7857142857142858
R_DFF_S0|45|B _DFF_S0|4 _DFF_S0|45|MID_SHUNT  3.84154647408
L_DFF_S0|45|RB _DFF_S0|45|MID_SHUNT _DFF_S0|5  2.1704737578552e-12
B_DFF_S0|T|1 _DFF_S0|T1 _DFF_S0|T|MID_SERIES JJMIT AREA=2.5
L_DFF_S0|T|P _DFF_S0|T|MID_SERIES 0  2e-13
R_DFF_S0|T|B _DFF_S0|T1 _DFF_S0|T|MID_SHUNT  2.7439617672
L_DFF_S0|T|RB _DFF_S0|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_S0|6|1 _DFF_S0|6 _DFF_S0|6|MID_SERIES JJMIT AREA=2.5
L_DFF_S0|6|P _DFF_S0|6|MID_SERIES 0  2e-13
R_DFF_S0|6|B _DFF_S0|6 _DFF_S0|6|MID_SHUNT  2.7439617672
L_DFF_S0|6|RB _DFF_S0|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_S0|I_1|B _DFF_S0|1 _DFF_S0|I_1|MID  2e-12
I_DFF_S0|I_1|B 0 _DFF_S0|I_1|MID  0.000175
L_DFF_S0|I_3|B _DFF_S0|3 _DFF_S0|I_3|MID  2e-12
I_DFF_S0|I_3|B 0 _DFF_S0|I_3|MID  0.00025
L_DFF_S0|I_T|B _DFF_S0|T1 _DFF_S0|I_T|MID  2e-12
I_DFF_S0|I_T|B 0 _DFF_S0|I_T|MID  0.000175
L_DFF_S0|I_6|B _DFF_S0|6 _DFF_S0|I_6|MID  2e-12
I_DFF_S0|I_6|B 0 _DFF_S0|I_6|MID  0.000175
L_XOR_S1|I_A1|B _XOR_S1|A1 _XOR_S1|I_A1|MID  2e-12
I_XOR_S1|I_A1|B 0 _XOR_S1|I_A1|MID  0.000175
L_XOR_S1|I_A3|B _XOR_S1|A3 _XOR_S1|I_A3|MID  2e-12
I_XOR_S1|I_A3|B 0 _XOR_S1|I_A3|MID  0.000175
L_XOR_S1|I_B1|B _XOR_S1|B1 _XOR_S1|I_B1|MID  2e-12
I_XOR_S1|I_B1|B 0 _XOR_S1|I_B1|MID  0.000175
L_XOR_S1|I_B3|B _XOR_S1|B3 _XOR_S1|I_B3|MID  2e-12
I_XOR_S1|I_B3|B 0 _XOR_S1|I_B3|MID  0.000175
L_XOR_S1|I_T1|B _XOR_S1|T1 _XOR_S1|I_T1|MID  2e-12
I_XOR_S1|I_T1|B 0 _XOR_S1|I_T1|MID  0.000175
L_XOR_S1|I_Q1|B _XOR_S1|Q1 _XOR_S1|I_Q1|MID  2e-12
I_XOR_S1|I_Q1|B 0 _XOR_S1|I_Q1|MID  0.000175
B_XOR_S1|A1|1 _XOR_S1|A1 _XOR_S1|A1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|A1|P _XOR_S1|A1|MID_SERIES 0  5e-13
R_XOR_S1|A1|B _XOR_S1|A1 _XOR_S1|A1|MID_SHUNT  2.7439617672
L_XOR_S1|A1|RB _XOR_S1|A1|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|A2|1 _XOR_S1|A2 _XOR_S1|A2|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|A2|P _XOR_S1|A2|MID_SERIES 0  5e-13
R_XOR_S1|A2|B _XOR_S1|A2 _XOR_S1|A2|MID_SHUNT  2.7439617672
L_XOR_S1|A2|RB _XOR_S1|A2|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|A3|1 _XOR_S1|A2 _XOR_S1|A3|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|A3|P _XOR_S1|A3|MID_SERIES _XOR_S1|A3  1.2e-12
R_XOR_S1|A3|B _XOR_S1|A2 _XOR_S1|A3|MID_SHUNT  2.7439617672
L_XOR_S1|A3|RB _XOR_S1|A3|MID_SHUNT _XOR_S1|A3  2.050338398468e-12
B_XOR_S1|B1|1 _XOR_S1|B1 _XOR_S1|B1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|B1|P _XOR_S1|B1|MID_SERIES 0  5e-13
R_XOR_S1|B1|B _XOR_S1|B1 _XOR_S1|B1|MID_SHUNT  2.7439617672
L_XOR_S1|B1|RB _XOR_S1|B1|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|B2|1 _XOR_S1|B2 _XOR_S1|B2|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|B2|P _XOR_S1|B2|MID_SERIES 0  5e-13
R_XOR_S1|B2|B _XOR_S1|B2 _XOR_S1|B2|MID_SHUNT  2.7439617672
L_XOR_S1|B2|RB _XOR_S1|B2|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|B3|1 _XOR_S1|B2 _XOR_S1|B3|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|B3|P _XOR_S1|B3|MID_SERIES _XOR_S1|B3  1.2e-12
R_XOR_S1|B3|B _XOR_S1|B2 _XOR_S1|B3|MID_SHUNT  2.7439617672
L_XOR_S1|B3|RB _XOR_S1|B3|MID_SHUNT _XOR_S1|B3  2.050338398468e-12
B_XOR_S1|T1|1 _XOR_S1|T1 _XOR_S1|T1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|T1|P _XOR_S1|T1|MID_SERIES 0  5e-13
R_XOR_S1|T1|B _XOR_S1|T1 _XOR_S1|T1|MID_SHUNT  2.7439617672
L_XOR_S1|T1|RB _XOR_S1|T1|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|T2|1 _XOR_S1|T2 _XOR_S1|ABTQ JJMIT AREA=2.0
R_XOR_S1|T2|B _XOR_S1|T2 _XOR_S1|T2|MID_SHUNT  3.429952209
L_XOR_S1|T2|RB _XOR_S1|T2|MID_SHUNT _XOR_S1|ABTQ  2.437922998085e-12
B_XOR_S1|AB|1 _XOR_S1|AB _XOR_S1|AB|MID_SERIES JJMIT AREA=2.0
L_XOR_S1|AB|P _XOR_S1|AB|MID_SERIES _XOR_S1|ABTQ  1.2e-12
R_XOR_S1|AB|B _XOR_S1|AB _XOR_S1|AB|MID_SHUNT  3.429952209
L_XOR_S1|AB|RB _XOR_S1|AB|MID_SHUNT _XOR_S1|ABTQ  2.437922998085e-12
B_XOR_S1|ABTQ|1 _XOR_S1|ABTQ _XOR_S1|ABTQ|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|ABTQ|P _XOR_S1|ABTQ|MID_SERIES 0  5e-13
R_XOR_S1|ABTQ|B _XOR_S1|ABTQ _XOR_S1|ABTQ|MID_SHUNT  2.7439617672
L_XOR_S1|ABTQ|RB _XOR_S1|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|Q1|1 _XOR_S1|Q1 _XOR_S1|Q1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|Q1|P _XOR_S1|Q1|MID_SERIES 0  5e-13
R_XOR_S1|Q1|B _XOR_S1|Q1 _XOR_S1|Q1|MID_SHUNT  2.7439617672
L_XOR_S1|Q1|RB _XOR_S1|Q1|MID_SHUNT 0  2.050338398468e-12
B_DFF_S2|1|1 _DFF_S2|1 _DFF_S2|1|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|1|P _DFF_S2|1|MID_SERIES 0  2e-13
R_DFF_S2|1|B _DFF_S2|1 _DFF_S2|1|MID_SHUNT  2.7439617672
L_DFF_S2|1|RB _DFF_S2|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|23|1 _DFF_S2|2 _DFF_S2|3 JJMIT AREA=1.7857142857142858
R_DFF_S2|23|B _DFF_S2|2 _DFF_S2|23|MID_SHUNT  3.84154647408
L_DFF_S2|23|RB _DFF_S2|23|MID_SHUNT _DFF_S2|3  2.1704737578552e-12
B_DFF_S2|3|1 _DFF_S2|3 _DFF_S2|3|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|3|P _DFF_S2|3|MID_SERIES 0  2e-13
R_DFF_S2|3|B _DFF_S2|3 _DFF_S2|3|MID_SHUNT  2.7439617672
L_DFF_S2|3|RB _DFF_S2|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|4|1 _DFF_S2|4 _DFF_S2|4|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|4|P _DFF_S2|4|MID_SERIES 0  2e-13
R_DFF_S2|4|B _DFF_S2|4 _DFF_S2|4|MID_SHUNT  2.7439617672
L_DFF_S2|4|RB _DFF_S2|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|45|1 _DFF_S2|4 _DFF_S2|5 JJMIT AREA=1.7857142857142858
R_DFF_S2|45|B _DFF_S2|4 _DFF_S2|45|MID_SHUNT  3.84154647408
L_DFF_S2|45|RB _DFF_S2|45|MID_SHUNT _DFF_S2|5  2.1704737578552e-12
B_DFF_S2|T|1 _DFF_S2|T1 _DFF_S2|T|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|T|P _DFF_S2|T|MID_SERIES 0  2e-13
R_DFF_S2|T|B _DFF_S2|T1 _DFF_S2|T|MID_SHUNT  2.7439617672
L_DFF_S2|T|RB _DFF_S2|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|6|1 _DFF_S2|6 _DFF_S2|6|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|6|P _DFF_S2|6|MID_SERIES 0  2e-13
R_DFF_S2|6|B _DFF_S2|6 _DFF_S2|6|MID_SHUNT  2.7439617672
L_DFF_S2|6|RB _DFF_S2|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_S2|I_1|B _DFF_S2|1 _DFF_S2|I_1|MID  2e-12
I_DFF_S2|I_1|B 0 _DFF_S2|I_1|MID  0.000175
L_DFF_S2|I_3|B _DFF_S2|3 _DFF_S2|I_3|MID  2e-12
I_DFF_S2|I_3|B 0 _DFF_S2|I_3|MID  0.00025
L_DFF_S2|I_T|B _DFF_S2|T1 _DFF_S2|I_T|MID  2e-12
I_DFF_S2|I_T|B 0 _DFF_S2|I_T|MID  0.000175
L_DFF_S2|I_6|B _DFF_S2|6 _DFF_S2|I_6|MID  2e-12
I_DFF_S2|I_6|B 0 _DFF_S2|I_6|MID  0.000175
L_INIT_0|_SPL_A|I_D1|B _INIT_0|_SPL_A|D1 _INIT_0|_SPL_A|I_D1|MID  2e-12
I_INIT_0|_SPL_A|I_D1|B 0 _INIT_0|_SPL_A|I_D1|MID  0.000175
L_INIT_0|_SPL_A|I_D2|B _INIT_0|_SPL_A|D2 _INIT_0|_SPL_A|I_D2|MID  2e-12
I_INIT_0|_SPL_A|I_D2|B 0 _INIT_0|_SPL_A|I_D2|MID  0.000245
L_INIT_0|_SPL_A|I_Q1|B _INIT_0|_SPL_A|QA1 _INIT_0|_SPL_A|I_Q1|MID  2e-12
I_INIT_0|_SPL_A|I_Q1|B 0 _INIT_0|_SPL_A|I_Q1|MID  0.000175
L_INIT_0|_SPL_A|I_Q2|B _INIT_0|_SPL_A|QB1 _INIT_0|_SPL_A|I_Q2|MID  2e-12
I_INIT_0|_SPL_A|I_Q2|B 0 _INIT_0|_SPL_A|I_Q2|MID  0.000175
B_INIT_0|_SPL_A|1|1 _INIT_0|_SPL_A|D1 _INIT_0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_A|1|P _INIT_0|_SPL_A|1|MID_SERIES 0  2e-13
R_INIT_0|_SPL_A|1|B _INIT_0|_SPL_A|D1 _INIT_0|_SPL_A|1|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_A|1|RB _INIT_0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_SPL_A|2|1 _INIT_0|_SPL_A|D2 _INIT_0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_A|2|P _INIT_0|_SPL_A|2|MID_SERIES 0  2e-13
R_INIT_0|_SPL_A|2|B _INIT_0|_SPL_A|D2 _INIT_0|_SPL_A|2|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_A|2|RB _INIT_0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_SPL_A|A|1 _INIT_0|_SPL_A|QA1 _INIT_0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_A|A|P _INIT_0|_SPL_A|A|MID_SERIES 0  2e-13
R_INIT_0|_SPL_A|A|B _INIT_0|_SPL_A|QA1 _INIT_0|_SPL_A|A|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_A|A|RB _INIT_0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_SPL_A|B|1 _INIT_0|_SPL_A|QB1 _INIT_0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_A|B|P _INIT_0|_SPL_A|B|MID_SERIES 0  2e-13
R_INIT_0|_SPL_A|B|B _INIT_0|_SPL_A|QB1 _INIT_0|_SPL_A|B|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_A|B|RB _INIT_0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
L_INIT_0|_SPL_B|I_D1|B _INIT_0|_SPL_B|D1 _INIT_0|_SPL_B|I_D1|MID  2e-12
I_INIT_0|_SPL_B|I_D1|B 0 _INIT_0|_SPL_B|I_D1|MID  0.000175
L_INIT_0|_SPL_B|I_D2|B _INIT_0|_SPL_B|D2 _INIT_0|_SPL_B|I_D2|MID  2e-12
I_INIT_0|_SPL_B|I_D2|B 0 _INIT_0|_SPL_B|I_D2|MID  0.000245
L_INIT_0|_SPL_B|I_Q1|B _INIT_0|_SPL_B|QA1 _INIT_0|_SPL_B|I_Q1|MID  2e-12
I_INIT_0|_SPL_B|I_Q1|B 0 _INIT_0|_SPL_B|I_Q1|MID  0.000175
L_INIT_0|_SPL_B|I_Q2|B _INIT_0|_SPL_B|QB1 _INIT_0|_SPL_B|I_Q2|MID  2e-12
I_INIT_0|_SPL_B|I_Q2|B 0 _INIT_0|_SPL_B|I_Q2|MID  0.000175
B_INIT_0|_SPL_B|1|1 _INIT_0|_SPL_B|D1 _INIT_0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_B|1|P _INIT_0|_SPL_B|1|MID_SERIES 0  2e-13
R_INIT_0|_SPL_B|1|B _INIT_0|_SPL_B|D1 _INIT_0|_SPL_B|1|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_B|1|RB _INIT_0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_SPL_B|2|1 _INIT_0|_SPL_B|D2 _INIT_0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_B|2|P _INIT_0|_SPL_B|2|MID_SERIES 0  2e-13
R_INIT_0|_SPL_B|2|B _INIT_0|_SPL_B|D2 _INIT_0|_SPL_B|2|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_B|2|RB _INIT_0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_SPL_B|A|1 _INIT_0|_SPL_B|QA1 _INIT_0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_B|A|P _INIT_0|_SPL_B|A|MID_SERIES 0  2e-13
R_INIT_0|_SPL_B|A|B _INIT_0|_SPL_B|QA1 _INIT_0|_SPL_B|A|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_B|A|RB _INIT_0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_SPL_B|B|1 _INIT_0|_SPL_B|QB1 _INIT_0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_SPL_B|B|P _INIT_0|_SPL_B|B|MID_SERIES 0  2e-13
R_INIT_0|_SPL_B|B|B _INIT_0|_SPL_B|QB1 _INIT_0|_SPL_B|B|MID_SHUNT  2.7439617672
L_INIT_0|_SPL_B|B|RB _INIT_0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_A|1|1 _INIT_0|_DFF_A|1 _INIT_0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_A|1|P _INIT_0|_DFF_A|1|MID_SERIES 0  2e-13
R_INIT_0|_DFF_A|1|B _INIT_0|_DFF_A|1 _INIT_0|_DFF_A|1|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_A|1|RB _INIT_0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_A|23|1 _INIT_0|_DFF_A|2 _INIT_0|_DFF_A|3 JJMIT AREA=1.7857142857142858
R_INIT_0|_DFF_A|23|B _INIT_0|_DFF_A|2 _INIT_0|_DFF_A|23|MID_SHUNT  3.84154647408
L_INIT_0|_DFF_A|23|RB _INIT_0|_DFF_A|23|MID_SHUNT _INIT_0|_DFF_A|3  2.1704737578552e-12
B_INIT_0|_DFF_A|3|1 _INIT_0|_DFF_A|3 _INIT_0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_A|3|P _INIT_0|_DFF_A|3|MID_SERIES 0  2e-13
R_INIT_0|_DFF_A|3|B _INIT_0|_DFF_A|3 _INIT_0|_DFF_A|3|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_A|3|RB _INIT_0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_A|4|1 _INIT_0|_DFF_A|4 _INIT_0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_A|4|P _INIT_0|_DFF_A|4|MID_SERIES 0  2e-13
R_INIT_0|_DFF_A|4|B _INIT_0|_DFF_A|4 _INIT_0|_DFF_A|4|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_A|4|RB _INIT_0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_A|45|1 _INIT_0|_DFF_A|4 _INIT_0|_DFF_A|5 JJMIT AREA=1.7857142857142858
R_INIT_0|_DFF_A|45|B _INIT_0|_DFF_A|4 _INIT_0|_DFF_A|45|MID_SHUNT  3.84154647408
L_INIT_0|_DFF_A|45|RB _INIT_0|_DFF_A|45|MID_SHUNT _INIT_0|_DFF_A|5  2.1704737578552e-12
B_INIT_0|_DFF_A|T|1 _INIT_0|_DFF_A|T1 _INIT_0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_A|T|P _INIT_0|_DFF_A|T|MID_SERIES 0  2e-13
R_INIT_0|_DFF_A|T|B _INIT_0|_DFF_A|T1 _INIT_0|_DFF_A|T|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_A|T|RB _INIT_0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_A|6|1 _INIT_0|_DFF_A|6 _INIT_0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_A|6|P _INIT_0|_DFF_A|6|MID_SERIES 0  2e-13
R_INIT_0|_DFF_A|6|B _INIT_0|_DFF_A|6 _INIT_0|_DFF_A|6|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_A|6|RB _INIT_0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
L_INIT_0|_DFF_A|I_1|B _INIT_0|_DFF_A|1 _INIT_0|_DFF_A|I_1|MID  2e-12
I_INIT_0|_DFF_A|I_1|B 0 _INIT_0|_DFF_A|I_1|MID  0.000175
L_INIT_0|_DFF_A|I_3|B _INIT_0|_DFF_A|3 _INIT_0|_DFF_A|I_3|MID  2e-12
I_INIT_0|_DFF_A|I_3|B 0 _INIT_0|_DFF_A|I_3|MID  0.00025
L_INIT_0|_DFF_A|I_T|B _INIT_0|_DFF_A|T1 _INIT_0|_DFF_A|I_T|MID  2e-12
I_INIT_0|_DFF_A|I_T|B 0 _INIT_0|_DFF_A|I_T|MID  0.000175
L_INIT_0|_DFF_A|I_6|B _INIT_0|_DFF_A|6 _INIT_0|_DFF_A|I_6|MID  2e-12
I_INIT_0|_DFF_A|I_6|B 0 _INIT_0|_DFF_A|I_6|MID  0.000175
B_INIT_0|_DFF_B|1|1 _INIT_0|_DFF_B|1 _INIT_0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_B|1|P _INIT_0|_DFF_B|1|MID_SERIES 0  2e-13
R_INIT_0|_DFF_B|1|B _INIT_0|_DFF_B|1 _INIT_0|_DFF_B|1|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_B|1|RB _INIT_0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_B|23|1 _INIT_0|_DFF_B|2 _INIT_0|_DFF_B|3 JJMIT AREA=1.7857142857142858
R_INIT_0|_DFF_B|23|B _INIT_0|_DFF_B|2 _INIT_0|_DFF_B|23|MID_SHUNT  3.84154647408
L_INIT_0|_DFF_B|23|RB _INIT_0|_DFF_B|23|MID_SHUNT _INIT_0|_DFF_B|3  2.1704737578552e-12
B_INIT_0|_DFF_B|3|1 _INIT_0|_DFF_B|3 _INIT_0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_B|3|P _INIT_0|_DFF_B|3|MID_SERIES 0  2e-13
R_INIT_0|_DFF_B|3|B _INIT_0|_DFF_B|3 _INIT_0|_DFF_B|3|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_B|3|RB _INIT_0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_B|4|1 _INIT_0|_DFF_B|4 _INIT_0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_B|4|P _INIT_0|_DFF_B|4|MID_SERIES 0  2e-13
R_INIT_0|_DFF_B|4|B _INIT_0|_DFF_B|4 _INIT_0|_DFF_B|4|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_B|4|RB _INIT_0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_B|45|1 _INIT_0|_DFF_B|4 _INIT_0|_DFF_B|5 JJMIT AREA=1.7857142857142858
R_INIT_0|_DFF_B|45|B _INIT_0|_DFF_B|4 _INIT_0|_DFF_B|45|MID_SHUNT  3.84154647408
L_INIT_0|_DFF_B|45|RB _INIT_0|_DFF_B|45|MID_SHUNT _INIT_0|_DFF_B|5  2.1704737578552e-12
B_INIT_0|_DFF_B|T|1 _INIT_0|_DFF_B|T1 _INIT_0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_B|T|P _INIT_0|_DFF_B|T|MID_SERIES 0  2e-13
R_INIT_0|_DFF_B|T|B _INIT_0|_DFF_B|T1 _INIT_0|_DFF_B|T|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_B|T|RB _INIT_0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_DFF_B|6|1 _INIT_0|_DFF_B|6 _INIT_0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_DFF_B|6|P _INIT_0|_DFF_B|6|MID_SERIES 0  2e-13
R_INIT_0|_DFF_B|6|B _INIT_0|_DFF_B|6 _INIT_0|_DFF_B|6|MID_SHUNT  2.7439617672
L_INIT_0|_DFF_B|6|RB _INIT_0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
L_INIT_0|_DFF_B|I_1|B _INIT_0|_DFF_B|1 _INIT_0|_DFF_B|I_1|MID  2e-12
I_INIT_0|_DFF_B|I_1|B 0 _INIT_0|_DFF_B|I_1|MID  0.000175
L_INIT_0|_DFF_B|I_3|B _INIT_0|_DFF_B|3 _INIT_0|_DFF_B|I_3|MID  2e-12
I_INIT_0|_DFF_B|I_3|B 0 _INIT_0|_DFF_B|I_3|MID  0.00025
L_INIT_0|_DFF_B|I_T|B _INIT_0|_DFF_B|T1 _INIT_0|_DFF_B|I_T|MID  2e-12
I_INIT_0|_DFF_B|I_T|B 0 _INIT_0|_DFF_B|I_T|MID  0.000175
L_INIT_0|_DFF_B|I_6|B _INIT_0|_DFF_B|6 _INIT_0|_DFF_B|I_6|MID  2e-12
I_INIT_0|_DFF_B|I_6|B 0 _INIT_0|_DFF_B|I_6|MID  0.000175
L_INIT_0|_XOR|I_A1|B _INIT_0|_XOR|A1 _INIT_0|_XOR|I_A1|MID  2e-12
I_INIT_0|_XOR|I_A1|B 0 _INIT_0|_XOR|I_A1|MID  0.000175
L_INIT_0|_XOR|I_A3|B _INIT_0|_XOR|A3 _INIT_0|_XOR|I_A3|MID  2e-12
I_INIT_0|_XOR|I_A3|B 0 _INIT_0|_XOR|I_A3|MID  0.000175
L_INIT_0|_XOR|I_B1|B _INIT_0|_XOR|B1 _INIT_0|_XOR|I_B1|MID  2e-12
I_INIT_0|_XOR|I_B1|B 0 _INIT_0|_XOR|I_B1|MID  0.000175
L_INIT_0|_XOR|I_B3|B _INIT_0|_XOR|B3 _INIT_0|_XOR|I_B3|MID  2e-12
I_INIT_0|_XOR|I_B3|B 0 _INIT_0|_XOR|I_B3|MID  0.000175
L_INIT_0|_XOR|I_T1|B _INIT_0|_XOR|T1 _INIT_0|_XOR|I_T1|MID  2e-12
I_INIT_0|_XOR|I_T1|B 0 _INIT_0|_XOR|I_T1|MID  0.000175
L_INIT_0|_XOR|I_Q1|B _INIT_0|_XOR|Q1 _INIT_0|_XOR|I_Q1|MID  2e-12
I_INIT_0|_XOR|I_Q1|B 0 _INIT_0|_XOR|I_Q1|MID  0.000175
B_INIT_0|_XOR|A1|1 _INIT_0|_XOR|A1 _INIT_0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|A1|P _INIT_0|_XOR|A1|MID_SERIES 0  5e-13
R_INIT_0|_XOR|A1|B _INIT_0|_XOR|A1 _INIT_0|_XOR|A1|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|A1|RB _INIT_0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
B_INIT_0|_XOR|A2|1 _INIT_0|_XOR|A2 _INIT_0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|A2|P _INIT_0|_XOR|A2|MID_SERIES 0  5e-13
R_INIT_0|_XOR|A2|B _INIT_0|_XOR|A2 _INIT_0|_XOR|A2|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|A2|RB _INIT_0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
B_INIT_0|_XOR|A3|1 _INIT_0|_XOR|A2 _INIT_0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|A3|P _INIT_0|_XOR|A3|MID_SERIES _INIT_0|_XOR|A3  1.2e-12
R_INIT_0|_XOR|A3|B _INIT_0|_XOR|A2 _INIT_0|_XOR|A3|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|A3|RB _INIT_0|_XOR|A3|MID_SHUNT _INIT_0|_XOR|A3  2.050338398468e-12
B_INIT_0|_XOR|B1|1 _INIT_0|_XOR|B1 _INIT_0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|B1|P _INIT_0|_XOR|B1|MID_SERIES 0  5e-13
R_INIT_0|_XOR|B1|B _INIT_0|_XOR|B1 _INIT_0|_XOR|B1|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|B1|RB _INIT_0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
B_INIT_0|_XOR|B2|1 _INIT_0|_XOR|B2 _INIT_0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|B2|P _INIT_0|_XOR|B2|MID_SERIES 0  5e-13
R_INIT_0|_XOR|B2|B _INIT_0|_XOR|B2 _INIT_0|_XOR|B2|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|B2|RB _INIT_0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
B_INIT_0|_XOR|B3|1 _INIT_0|_XOR|B2 _INIT_0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|B3|P _INIT_0|_XOR|B3|MID_SERIES _INIT_0|_XOR|B3  1.2e-12
R_INIT_0|_XOR|B3|B _INIT_0|_XOR|B2 _INIT_0|_XOR|B3|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|B3|RB _INIT_0|_XOR|B3|MID_SHUNT _INIT_0|_XOR|B3  2.050338398468e-12
B_INIT_0|_XOR|T1|1 _INIT_0|_XOR|T1 _INIT_0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|T1|P _INIT_0|_XOR|T1|MID_SERIES 0  5e-13
R_INIT_0|_XOR|T1|B _INIT_0|_XOR|T1 _INIT_0|_XOR|T1|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|T1|RB _INIT_0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
B_INIT_0|_XOR|T2|1 _INIT_0|_XOR|T2 _INIT_0|_XOR|ABTQ JJMIT AREA=2.0
R_INIT_0|_XOR|T2|B _INIT_0|_XOR|T2 _INIT_0|_XOR|T2|MID_SHUNT  3.429952209
L_INIT_0|_XOR|T2|RB _INIT_0|_XOR|T2|MID_SHUNT _INIT_0|_XOR|ABTQ  2.437922998085e-12
B_INIT_0|_XOR|AB|1 _INIT_0|_XOR|AB _INIT_0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
L_INIT_0|_XOR|AB|P _INIT_0|_XOR|AB|MID_SERIES _INIT_0|_XOR|ABTQ  1.2e-12
R_INIT_0|_XOR|AB|B _INIT_0|_XOR|AB _INIT_0|_XOR|AB|MID_SHUNT  3.429952209
L_INIT_0|_XOR|AB|RB _INIT_0|_XOR|AB|MID_SHUNT _INIT_0|_XOR|ABTQ  2.437922998085e-12
B_INIT_0|_XOR|ABTQ|1 _INIT_0|_XOR|ABTQ _INIT_0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|ABTQ|P _INIT_0|_XOR|ABTQ|MID_SERIES 0  5e-13
R_INIT_0|_XOR|ABTQ|B _INIT_0|_XOR|ABTQ _INIT_0|_XOR|ABTQ|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|ABTQ|RB _INIT_0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_INIT_0|_XOR|Q1|1 _INIT_0|_XOR|Q1 _INIT_0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_XOR|Q1|P _INIT_0|_XOR|Q1|MID_SERIES 0  5e-13
R_INIT_0|_XOR|Q1|B _INIT_0|_XOR|Q1 _INIT_0|_XOR|Q1|MID_SHUNT  2.7439617672
L_INIT_0|_XOR|Q1|RB _INIT_0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
L_INIT_0|_AND|I_A1|B _INIT_0|_AND|A1 _INIT_0|_AND|I_A1|MID  2e-12
I_INIT_0|_AND|I_A1|B 0 _INIT_0|_AND|I_A1|MID  0.000175
L_INIT_0|_AND|I_B1|B _INIT_0|_AND|B1 _INIT_0|_AND|I_B1|MID  2e-12
I_INIT_0|_AND|I_B1|B 0 _INIT_0|_AND|I_B1|MID  0.000175
L_INIT_0|_AND|I_Q3|B _INIT_0|_AND|Q3 _INIT_0|_AND|I_Q3|MID  2e-12
I_INIT_0|_AND|I_Q3|B 0 _INIT_0|_AND|I_Q3|MID  7.5e-05
L_INIT_0|_AND|I_Q2|B _INIT_0|_AND|Q2 _INIT_0|_AND|I_Q2|MID  2e-12
I_INIT_0|_AND|I_Q2|B 0 _INIT_0|_AND|I_Q2|MID  0.000175
L_INIT_0|_AND|I_Q1|B _INIT_0|_AND|Q1 _INIT_0|_AND|I_Q1|MID  2e-12
I_INIT_0|_AND|I_Q1|B 0 _INIT_0|_AND|I_Q1|MID  0.000175
B_INIT_0|_AND|A1|1 _INIT_0|_AND|A1 _INIT_0|_AND|A1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_AND|A1|P _INIT_0|_AND|A1|MID_SERIES 0  2e-13
R_INIT_0|_AND|A1|B _INIT_0|_AND|A1 _INIT_0|_AND|A1|MID_SHUNT  2.7439617672
L_INIT_0|_AND|A1|RB _INIT_0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_AND|A2|1 _INIT_0|_AND|A2 _INIT_0|_AND|A2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_AND|A2|P _INIT_0|_AND|A2|MID_SERIES 0  2e-13
R_INIT_0|_AND|A2|B _INIT_0|_AND|A2 _INIT_0|_AND|A2|MID_SHUNT  2.7439617672
L_INIT_0|_AND|A2|RB _INIT_0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_AND|A12|1 _INIT_0|_AND|A2 _INIT_0|_AND|A3 JJMIT AREA=1.7857142857142858
R_INIT_0|_AND|A12|B _INIT_0|_AND|A2 _INIT_0|_AND|A12|MID_SHUNT  3.84154647408
L_INIT_0|_AND|A12|RB _INIT_0|_AND|A12|MID_SHUNT _INIT_0|_AND|A3  2.1704737578552e-12
B_INIT_0|_AND|B1|1 _INIT_0|_AND|B1 _INIT_0|_AND|B1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_AND|B1|P _INIT_0|_AND|B1|MID_SERIES 0  2e-13
R_INIT_0|_AND|B1|B _INIT_0|_AND|B1 _INIT_0|_AND|B1|MID_SHUNT  2.7439617672
L_INIT_0|_AND|B1|RB _INIT_0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_AND|B2|1 _INIT_0|_AND|B2 _INIT_0|_AND|B2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_AND|B2|P _INIT_0|_AND|B2|MID_SERIES 0  2e-13
R_INIT_0|_AND|B2|B _INIT_0|_AND|B2 _INIT_0|_AND|B2|MID_SHUNT  2.7439617672
L_INIT_0|_AND|B2|RB _INIT_0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_AND|B12|1 _INIT_0|_AND|B2 _INIT_0|_AND|B3 JJMIT AREA=1.7857142857142858
R_INIT_0|_AND|B12|B _INIT_0|_AND|B2 _INIT_0|_AND|B12|MID_SHUNT  3.84154647408
L_INIT_0|_AND|B12|RB _INIT_0|_AND|B12|MID_SHUNT _INIT_0|_AND|B3  2.1704737578552e-12
B_INIT_0|_AND|Q2|1 _INIT_0|_AND|Q2 _INIT_0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_AND|Q2|P _INIT_0|_AND|Q2|MID_SERIES 0  2e-13
R_INIT_0|_AND|Q2|B _INIT_0|_AND|Q2 _INIT_0|_AND|Q2|MID_SHUNT  2.7439617672
L_INIT_0|_AND|Q2|RB _INIT_0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
B_INIT_0|_AND|Q1|1 _INIT_0|_AND|Q1 _INIT_0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
L_INIT_0|_AND|Q1|P _INIT_0|_AND|Q1|MID_SERIES 0  2e-13
R_INIT_0|_AND|Q1|B _INIT_0|_AND|Q1 _INIT_0|_AND|Q1|MID_SHUNT  2.7439617672
L_INIT_0|_AND|Q1|RB _INIT_0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
L_INIT_1|_SPL_A|I_D1|B _INIT_1|_SPL_A|D1 _INIT_1|_SPL_A|I_D1|MID  2e-12
I_INIT_1|_SPL_A|I_D1|B 0 _INIT_1|_SPL_A|I_D1|MID  0.000175
L_INIT_1|_SPL_A|I_D2|B _INIT_1|_SPL_A|D2 _INIT_1|_SPL_A|I_D2|MID  2e-12
I_INIT_1|_SPL_A|I_D2|B 0 _INIT_1|_SPL_A|I_D2|MID  0.000245
L_INIT_1|_SPL_A|I_Q1|B _INIT_1|_SPL_A|QA1 _INIT_1|_SPL_A|I_Q1|MID  2e-12
I_INIT_1|_SPL_A|I_Q1|B 0 _INIT_1|_SPL_A|I_Q1|MID  0.000175
L_INIT_1|_SPL_A|I_Q2|B _INIT_1|_SPL_A|QB1 _INIT_1|_SPL_A|I_Q2|MID  2e-12
I_INIT_1|_SPL_A|I_Q2|B 0 _INIT_1|_SPL_A|I_Q2|MID  0.000175
B_INIT_1|_SPL_A|1|1 _INIT_1|_SPL_A|D1 _INIT_1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_A|1|P _INIT_1|_SPL_A|1|MID_SERIES 0  2e-13
R_INIT_1|_SPL_A|1|B _INIT_1|_SPL_A|D1 _INIT_1|_SPL_A|1|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_A|1|RB _INIT_1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_SPL_A|2|1 _INIT_1|_SPL_A|D2 _INIT_1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_A|2|P _INIT_1|_SPL_A|2|MID_SERIES 0  2e-13
R_INIT_1|_SPL_A|2|B _INIT_1|_SPL_A|D2 _INIT_1|_SPL_A|2|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_A|2|RB _INIT_1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_SPL_A|A|1 _INIT_1|_SPL_A|QA1 _INIT_1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_A|A|P _INIT_1|_SPL_A|A|MID_SERIES 0  2e-13
R_INIT_1|_SPL_A|A|B _INIT_1|_SPL_A|QA1 _INIT_1|_SPL_A|A|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_A|A|RB _INIT_1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_SPL_A|B|1 _INIT_1|_SPL_A|QB1 _INIT_1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_A|B|P _INIT_1|_SPL_A|B|MID_SERIES 0  2e-13
R_INIT_1|_SPL_A|B|B _INIT_1|_SPL_A|QB1 _INIT_1|_SPL_A|B|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_A|B|RB _INIT_1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
L_INIT_1|_SPL_B|I_D1|B _INIT_1|_SPL_B|D1 _INIT_1|_SPL_B|I_D1|MID  2e-12
I_INIT_1|_SPL_B|I_D1|B 0 _INIT_1|_SPL_B|I_D1|MID  0.000175
L_INIT_1|_SPL_B|I_D2|B _INIT_1|_SPL_B|D2 _INIT_1|_SPL_B|I_D2|MID  2e-12
I_INIT_1|_SPL_B|I_D2|B 0 _INIT_1|_SPL_B|I_D2|MID  0.000245
L_INIT_1|_SPL_B|I_Q1|B _INIT_1|_SPL_B|QA1 _INIT_1|_SPL_B|I_Q1|MID  2e-12
I_INIT_1|_SPL_B|I_Q1|B 0 _INIT_1|_SPL_B|I_Q1|MID  0.000175
L_INIT_1|_SPL_B|I_Q2|B _INIT_1|_SPL_B|QB1 _INIT_1|_SPL_B|I_Q2|MID  2e-12
I_INIT_1|_SPL_B|I_Q2|B 0 _INIT_1|_SPL_B|I_Q2|MID  0.000175
B_INIT_1|_SPL_B|1|1 _INIT_1|_SPL_B|D1 _INIT_1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_B|1|P _INIT_1|_SPL_B|1|MID_SERIES 0  2e-13
R_INIT_1|_SPL_B|1|B _INIT_1|_SPL_B|D1 _INIT_1|_SPL_B|1|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_B|1|RB _INIT_1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_SPL_B|2|1 _INIT_1|_SPL_B|D2 _INIT_1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_B|2|P _INIT_1|_SPL_B|2|MID_SERIES 0  2e-13
R_INIT_1|_SPL_B|2|B _INIT_1|_SPL_B|D2 _INIT_1|_SPL_B|2|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_B|2|RB _INIT_1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_SPL_B|A|1 _INIT_1|_SPL_B|QA1 _INIT_1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_B|A|P _INIT_1|_SPL_B|A|MID_SERIES 0  2e-13
R_INIT_1|_SPL_B|A|B _INIT_1|_SPL_B|QA1 _INIT_1|_SPL_B|A|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_B|A|RB _INIT_1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_SPL_B|B|1 _INIT_1|_SPL_B|QB1 _INIT_1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_SPL_B|B|P _INIT_1|_SPL_B|B|MID_SERIES 0  2e-13
R_INIT_1|_SPL_B|B|B _INIT_1|_SPL_B|QB1 _INIT_1|_SPL_B|B|MID_SHUNT  2.7439617672
L_INIT_1|_SPL_B|B|RB _INIT_1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_A|1|1 _INIT_1|_DFF_A|1 _INIT_1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_A|1|P _INIT_1|_DFF_A|1|MID_SERIES 0  2e-13
R_INIT_1|_DFF_A|1|B _INIT_1|_DFF_A|1 _INIT_1|_DFF_A|1|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_A|1|RB _INIT_1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_A|23|1 _INIT_1|_DFF_A|2 _INIT_1|_DFF_A|3 JJMIT AREA=1.7857142857142858
R_INIT_1|_DFF_A|23|B _INIT_1|_DFF_A|2 _INIT_1|_DFF_A|23|MID_SHUNT  3.84154647408
L_INIT_1|_DFF_A|23|RB _INIT_1|_DFF_A|23|MID_SHUNT _INIT_1|_DFF_A|3  2.1704737578552e-12
B_INIT_1|_DFF_A|3|1 _INIT_1|_DFF_A|3 _INIT_1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_A|3|P _INIT_1|_DFF_A|3|MID_SERIES 0  2e-13
R_INIT_1|_DFF_A|3|B _INIT_1|_DFF_A|3 _INIT_1|_DFF_A|3|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_A|3|RB _INIT_1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_A|4|1 _INIT_1|_DFF_A|4 _INIT_1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_A|4|P _INIT_1|_DFF_A|4|MID_SERIES 0  2e-13
R_INIT_1|_DFF_A|4|B _INIT_1|_DFF_A|4 _INIT_1|_DFF_A|4|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_A|4|RB _INIT_1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_A|45|1 _INIT_1|_DFF_A|4 _INIT_1|_DFF_A|5 JJMIT AREA=1.7857142857142858
R_INIT_1|_DFF_A|45|B _INIT_1|_DFF_A|4 _INIT_1|_DFF_A|45|MID_SHUNT  3.84154647408
L_INIT_1|_DFF_A|45|RB _INIT_1|_DFF_A|45|MID_SHUNT _INIT_1|_DFF_A|5  2.1704737578552e-12
B_INIT_1|_DFF_A|T|1 _INIT_1|_DFF_A|T1 _INIT_1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_A|T|P _INIT_1|_DFF_A|T|MID_SERIES 0  2e-13
R_INIT_1|_DFF_A|T|B _INIT_1|_DFF_A|T1 _INIT_1|_DFF_A|T|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_A|T|RB _INIT_1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_A|6|1 _INIT_1|_DFF_A|6 _INIT_1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_A|6|P _INIT_1|_DFF_A|6|MID_SERIES 0  2e-13
R_INIT_1|_DFF_A|6|B _INIT_1|_DFF_A|6 _INIT_1|_DFF_A|6|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_A|6|RB _INIT_1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
L_INIT_1|_DFF_A|I_1|B _INIT_1|_DFF_A|1 _INIT_1|_DFF_A|I_1|MID  2e-12
I_INIT_1|_DFF_A|I_1|B 0 _INIT_1|_DFF_A|I_1|MID  0.000175
L_INIT_1|_DFF_A|I_3|B _INIT_1|_DFF_A|3 _INIT_1|_DFF_A|I_3|MID  2e-12
I_INIT_1|_DFF_A|I_3|B 0 _INIT_1|_DFF_A|I_3|MID  0.00025
L_INIT_1|_DFF_A|I_T|B _INIT_1|_DFF_A|T1 _INIT_1|_DFF_A|I_T|MID  2e-12
I_INIT_1|_DFF_A|I_T|B 0 _INIT_1|_DFF_A|I_T|MID  0.000175
L_INIT_1|_DFF_A|I_6|B _INIT_1|_DFF_A|6 _INIT_1|_DFF_A|I_6|MID  2e-12
I_INIT_1|_DFF_A|I_6|B 0 _INIT_1|_DFF_A|I_6|MID  0.000175
B_INIT_1|_DFF_B|1|1 _INIT_1|_DFF_B|1 _INIT_1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_B|1|P _INIT_1|_DFF_B|1|MID_SERIES 0  2e-13
R_INIT_1|_DFF_B|1|B _INIT_1|_DFF_B|1 _INIT_1|_DFF_B|1|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_B|1|RB _INIT_1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_B|23|1 _INIT_1|_DFF_B|2 _INIT_1|_DFF_B|3 JJMIT AREA=1.7857142857142858
R_INIT_1|_DFF_B|23|B _INIT_1|_DFF_B|2 _INIT_1|_DFF_B|23|MID_SHUNT  3.84154647408
L_INIT_1|_DFF_B|23|RB _INIT_1|_DFF_B|23|MID_SHUNT _INIT_1|_DFF_B|3  2.1704737578552e-12
B_INIT_1|_DFF_B|3|1 _INIT_1|_DFF_B|3 _INIT_1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_B|3|P _INIT_1|_DFF_B|3|MID_SERIES 0  2e-13
R_INIT_1|_DFF_B|3|B _INIT_1|_DFF_B|3 _INIT_1|_DFF_B|3|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_B|3|RB _INIT_1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_B|4|1 _INIT_1|_DFF_B|4 _INIT_1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_B|4|P _INIT_1|_DFF_B|4|MID_SERIES 0  2e-13
R_INIT_1|_DFF_B|4|B _INIT_1|_DFF_B|4 _INIT_1|_DFF_B|4|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_B|4|RB _INIT_1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_B|45|1 _INIT_1|_DFF_B|4 _INIT_1|_DFF_B|5 JJMIT AREA=1.7857142857142858
R_INIT_1|_DFF_B|45|B _INIT_1|_DFF_B|4 _INIT_1|_DFF_B|45|MID_SHUNT  3.84154647408
L_INIT_1|_DFF_B|45|RB _INIT_1|_DFF_B|45|MID_SHUNT _INIT_1|_DFF_B|5  2.1704737578552e-12
B_INIT_1|_DFF_B|T|1 _INIT_1|_DFF_B|T1 _INIT_1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_B|T|P _INIT_1|_DFF_B|T|MID_SERIES 0  2e-13
R_INIT_1|_DFF_B|T|B _INIT_1|_DFF_B|T1 _INIT_1|_DFF_B|T|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_B|T|RB _INIT_1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_DFF_B|6|1 _INIT_1|_DFF_B|6 _INIT_1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_DFF_B|6|P _INIT_1|_DFF_B|6|MID_SERIES 0  2e-13
R_INIT_1|_DFF_B|6|B _INIT_1|_DFF_B|6 _INIT_1|_DFF_B|6|MID_SHUNT  2.7439617672
L_INIT_1|_DFF_B|6|RB _INIT_1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
L_INIT_1|_DFF_B|I_1|B _INIT_1|_DFF_B|1 _INIT_1|_DFF_B|I_1|MID  2e-12
I_INIT_1|_DFF_B|I_1|B 0 _INIT_1|_DFF_B|I_1|MID  0.000175
L_INIT_1|_DFF_B|I_3|B _INIT_1|_DFF_B|3 _INIT_1|_DFF_B|I_3|MID  2e-12
I_INIT_1|_DFF_B|I_3|B 0 _INIT_1|_DFF_B|I_3|MID  0.00025
L_INIT_1|_DFF_B|I_T|B _INIT_1|_DFF_B|T1 _INIT_1|_DFF_B|I_T|MID  2e-12
I_INIT_1|_DFF_B|I_T|B 0 _INIT_1|_DFF_B|I_T|MID  0.000175
L_INIT_1|_DFF_B|I_6|B _INIT_1|_DFF_B|6 _INIT_1|_DFF_B|I_6|MID  2e-12
I_INIT_1|_DFF_B|I_6|B 0 _INIT_1|_DFF_B|I_6|MID  0.000175
L_INIT_1|_XOR|I_A1|B _INIT_1|_XOR|A1 _INIT_1|_XOR|I_A1|MID  2e-12
I_INIT_1|_XOR|I_A1|B 0 _INIT_1|_XOR|I_A1|MID  0.000175
L_INIT_1|_XOR|I_A3|B _INIT_1|_XOR|A3 _INIT_1|_XOR|I_A3|MID  2e-12
I_INIT_1|_XOR|I_A3|B 0 _INIT_1|_XOR|I_A3|MID  0.000175
L_INIT_1|_XOR|I_B1|B _INIT_1|_XOR|B1 _INIT_1|_XOR|I_B1|MID  2e-12
I_INIT_1|_XOR|I_B1|B 0 _INIT_1|_XOR|I_B1|MID  0.000175
L_INIT_1|_XOR|I_B3|B _INIT_1|_XOR|B3 _INIT_1|_XOR|I_B3|MID  2e-12
I_INIT_1|_XOR|I_B3|B 0 _INIT_1|_XOR|I_B3|MID  0.000175
L_INIT_1|_XOR|I_T1|B _INIT_1|_XOR|T1 _INIT_1|_XOR|I_T1|MID  2e-12
I_INIT_1|_XOR|I_T1|B 0 _INIT_1|_XOR|I_T1|MID  0.000175
L_INIT_1|_XOR|I_Q1|B _INIT_1|_XOR|Q1 _INIT_1|_XOR|I_Q1|MID  2e-12
I_INIT_1|_XOR|I_Q1|B 0 _INIT_1|_XOR|I_Q1|MID  0.000175
B_INIT_1|_XOR|A1|1 _INIT_1|_XOR|A1 _INIT_1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|A1|P _INIT_1|_XOR|A1|MID_SERIES 0  5e-13
R_INIT_1|_XOR|A1|B _INIT_1|_XOR|A1 _INIT_1|_XOR|A1|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|A1|RB _INIT_1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
B_INIT_1|_XOR|A2|1 _INIT_1|_XOR|A2 _INIT_1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|A2|P _INIT_1|_XOR|A2|MID_SERIES 0  5e-13
R_INIT_1|_XOR|A2|B _INIT_1|_XOR|A2 _INIT_1|_XOR|A2|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|A2|RB _INIT_1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
B_INIT_1|_XOR|A3|1 _INIT_1|_XOR|A2 _INIT_1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|A3|P _INIT_1|_XOR|A3|MID_SERIES _INIT_1|_XOR|A3  1.2e-12
R_INIT_1|_XOR|A3|B _INIT_1|_XOR|A2 _INIT_1|_XOR|A3|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|A3|RB _INIT_1|_XOR|A3|MID_SHUNT _INIT_1|_XOR|A3  2.050338398468e-12
B_INIT_1|_XOR|B1|1 _INIT_1|_XOR|B1 _INIT_1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|B1|P _INIT_1|_XOR|B1|MID_SERIES 0  5e-13
R_INIT_1|_XOR|B1|B _INIT_1|_XOR|B1 _INIT_1|_XOR|B1|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|B1|RB _INIT_1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
B_INIT_1|_XOR|B2|1 _INIT_1|_XOR|B2 _INIT_1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|B2|P _INIT_1|_XOR|B2|MID_SERIES 0  5e-13
R_INIT_1|_XOR|B2|B _INIT_1|_XOR|B2 _INIT_1|_XOR|B2|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|B2|RB _INIT_1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
B_INIT_1|_XOR|B3|1 _INIT_1|_XOR|B2 _INIT_1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|B3|P _INIT_1|_XOR|B3|MID_SERIES _INIT_1|_XOR|B3  1.2e-12
R_INIT_1|_XOR|B3|B _INIT_1|_XOR|B2 _INIT_1|_XOR|B3|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|B3|RB _INIT_1|_XOR|B3|MID_SHUNT _INIT_1|_XOR|B3  2.050338398468e-12
B_INIT_1|_XOR|T1|1 _INIT_1|_XOR|T1 _INIT_1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|T1|P _INIT_1|_XOR|T1|MID_SERIES 0  5e-13
R_INIT_1|_XOR|T1|B _INIT_1|_XOR|T1 _INIT_1|_XOR|T1|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|T1|RB _INIT_1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
B_INIT_1|_XOR|T2|1 _INIT_1|_XOR|T2 _INIT_1|_XOR|ABTQ JJMIT AREA=2.0
R_INIT_1|_XOR|T2|B _INIT_1|_XOR|T2 _INIT_1|_XOR|T2|MID_SHUNT  3.429952209
L_INIT_1|_XOR|T2|RB _INIT_1|_XOR|T2|MID_SHUNT _INIT_1|_XOR|ABTQ  2.437922998085e-12
B_INIT_1|_XOR|AB|1 _INIT_1|_XOR|AB _INIT_1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
L_INIT_1|_XOR|AB|P _INIT_1|_XOR|AB|MID_SERIES _INIT_1|_XOR|ABTQ  1.2e-12
R_INIT_1|_XOR|AB|B _INIT_1|_XOR|AB _INIT_1|_XOR|AB|MID_SHUNT  3.429952209
L_INIT_1|_XOR|AB|RB _INIT_1|_XOR|AB|MID_SHUNT _INIT_1|_XOR|ABTQ  2.437922998085e-12
B_INIT_1|_XOR|ABTQ|1 _INIT_1|_XOR|ABTQ _INIT_1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|ABTQ|P _INIT_1|_XOR|ABTQ|MID_SERIES 0  5e-13
R_INIT_1|_XOR|ABTQ|B _INIT_1|_XOR|ABTQ _INIT_1|_XOR|ABTQ|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|ABTQ|RB _INIT_1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_INIT_1|_XOR|Q1|1 _INIT_1|_XOR|Q1 _INIT_1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_XOR|Q1|P _INIT_1|_XOR|Q1|MID_SERIES 0  5e-13
R_INIT_1|_XOR|Q1|B _INIT_1|_XOR|Q1 _INIT_1|_XOR|Q1|MID_SHUNT  2.7439617672
L_INIT_1|_XOR|Q1|RB _INIT_1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
L_INIT_1|_AND|I_A1|B _INIT_1|_AND|A1 _INIT_1|_AND|I_A1|MID  2e-12
I_INIT_1|_AND|I_A1|B 0 _INIT_1|_AND|I_A1|MID  0.000175
L_INIT_1|_AND|I_B1|B _INIT_1|_AND|B1 _INIT_1|_AND|I_B1|MID  2e-12
I_INIT_1|_AND|I_B1|B 0 _INIT_1|_AND|I_B1|MID  0.000175
L_INIT_1|_AND|I_Q3|B _INIT_1|_AND|Q3 _INIT_1|_AND|I_Q3|MID  2e-12
I_INIT_1|_AND|I_Q3|B 0 _INIT_1|_AND|I_Q3|MID  7.5e-05
L_INIT_1|_AND|I_Q2|B _INIT_1|_AND|Q2 _INIT_1|_AND|I_Q2|MID  2e-12
I_INIT_1|_AND|I_Q2|B 0 _INIT_1|_AND|I_Q2|MID  0.000175
L_INIT_1|_AND|I_Q1|B _INIT_1|_AND|Q1 _INIT_1|_AND|I_Q1|MID  2e-12
I_INIT_1|_AND|I_Q1|B 0 _INIT_1|_AND|I_Q1|MID  0.000175
B_INIT_1|_AND|A1|1 _INIT_1|_AND|A1 _INIT_1|_AND|A1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_AND|A1|P _INIT_1|_AND|A1|MID_SERIES 0  2e-13
R_INIT_1|_AND|A1|B _INIT_1|_AND|A1 _INIT_1|_AND|A1|MID_SHUNT  2.7439617672
L_INIT_1|_AND|A1|RB _INIT_1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_AND|A2|1 _INIT_1|_AND|A2 _INIT_1|_AND|A2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_AND|A2|P _INIT_1|_AND|A2|MID_SERIES 0  2e-13
R_INIT_1|_AND|A2|B _INIT_1|_AND|A2 _INIT_1|_AND|A2|MID_SHUNT  2.7439617672
L_INIT_1|_AND|A2|RB _INIT_1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_AND|A12|1 _INIT_1|_AND|A2 _INIT_1|_AND|A3 JJMIT AREA=1.7857142857142858
R_INIT_1|_AND|A12|B _INIT_1|_AND|A2 _INIT_1|_AND|A12|MID_SHUNT  3.84154647408
L_INIT_1|_AND|A12|RB _INIT_1|_AND|A12|MID_SHUNT _INIT_1|_AND|A3  2.1704737578552e-12
B_INIT_1|_AND|B1|1 _INIT_1|_AND|B1 _INIT_1|_AND|B1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_AND|B1|P _INIT_1|_AND|B1|MID_SERIES 0  2e-13
R_INIT_1|_AND|B1|B _INIT_1|_AND|B1 _INIT_1|_AND|B1|MID_SHUNT  2.7439617672
L_INIT_1|_AND|B1|RB _INIT_1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_AND|B2|1 _INIT_1|_AND|B2 _INIT_1|_AND|B2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_AND|B2|P _INIT_1|_AND|B2|MID_SERIES 0  2e-13
R_INIT_1|_AND|B2|B _INIT_1|_AND|B2 _INIT_1|_AND|B2|MID_SHUNT  2.7439617672
L_INIT_1|_AND|B2|RB _INIT_1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_AND|B12|1 _INIT_1|_AND|B2 _INIT_1|_AND|B3 JJMIT AREA=1.7857142857142858
R_INIT_1|_AND|B12|B _INIT_1|_AND|B2 _INIT_1|_AND|B12|MID_SHUNT  3.84154647408
L_INIT_1|_AND|B12|RB _INIT_1|_AND|B12|MID_SHUNT _INIT_1|_AND|B3  2.1704737578552e-12
B_INIT_1|_AND|Q2|1 _INIT_1|_AND|Q2 _INIT_1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_AND|Q2|P _INIT_1|_AND|Q2|MID_SERIES 0  2e-13
R_INIT_1|_AND|Q2|B _INIT_1|_AND|Q2 _INIT_1|_AND|Q2|MID_SHUNT  2.7439617672
L_INIT_1|_AND|Q2|RB _INIT_1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
B_INIT_1|_AND|Q1|1 _INIT_1|_AND|Q1 _INIT_1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
L_INIT_1|_AND|Q1|P _INIT_1|_AND|Q1|MID_SERIES 0  2e-13
R_INIT_1|_AND|Q1|B _INIT_1|_AND|Q1 _INIT_1|_AND|Q1|MID_SHUNT  2.7439617672
L_INIT_1|_AND|Q1|RB _INIT_1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_SPL_G1|I_D1|B _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|I_D1|MID  2e-12
I_PG_01|_SPL_G1|I_D1|B 0 _PG_01|_SPL_G1|I_D1|MID  0.000175
L_PG_01|_SPL_G1|I_D2|B _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|I_D2|MID  2e-12
I_PG_01|_SPL_G1|I_D2|B 0 _PG_01|_SPL_G1|I_D2|MID  0.000245
L_PG_01|_SPL_G1|I_Q1|B _PG_01|_SPL_G1|QA1 _PG_01|_SPL_G1|I_Q1|MID  2e-12
I_PG_01|_SPL_G1|I_Q1|B 0 _PG_01|_SPL_G1|I_Q1|MID  0.000175
L_PG_01|_SPL_G1|I_Q2|B _PG_01|_SPL_G1|QB1 _PG_01|_SPL_G1|I_Q2|MID  2e-12
I_PG_01|_SPL_G1|I_Q2|B 0 _PG_01|_SPL_G1|I_Q2|MID  0.000175
B_PG_01|_SPL_G1|1|1 _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|1|P _PG_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|1|B _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|1|RB _PG_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_G1|2|1 _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|2|P _PG_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|2|B _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|2|RB _PG_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_G1|A|1 _PG_01|_SPL_G1|QA1 _PG_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|A|P _PG_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|A|B _PG_01|_SPL_G1|QA1 _PG_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|A|RB _PG_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_G1|B|1 _PG_01|_SPL_G1|QB1 _PG_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|B|P _PG_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|B|B _PG_01|_SPL_G1|QB1 _PG_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|B|RB _PG_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_SPL_P1|I_D1|B _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|I_D1|MID  2e-12
I_PG_01|_SPL_P1|I_D1|B 0 _PG_01|_SPL_P1|I_D1|MID  0.000175
L_PG_01|_SPL_P1|I_D2|B _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|I_D2|MID  2e-12
I_PG_01|_SPL_P1|I_D2|B 0 _PG_01|_SPL_P1|I_D2|MID  0.000245
L_PG_01|_SPL_P1|I_Q1|B _PG_01|_SPL_P1|QA1 _PG_01|_SPL_P1|I_Q1|MID  2e-12
I_PG_01|_SPL_P1|I_Q1|B 0 _PG_01|_SPL_P1|I_Q1|MID  0.000175
L_PG_01|_SPL_P1|I_Q2|B _PG_01|_SPL_P1|QB1 _PG_01|_SPL_P1|I_Q2|MID  2e-12
I_PG_01|_SPL_P1|I_Q2|B 0 _PG_01|_SPL_P1|I_Q2|MID  0.000175
B_PG_01|_SPL_P1|1|1 _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|1|P _PG_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|1|B _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|1|RB _PG_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_P1|2|1 _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|2|P _PG_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|2|B _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|2|RB _PG_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_P1|A|1 _PG_01|_SPL_P1|QA1 _PG_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|A|P _PG_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|A|B _PG_01|_SPL_P1|QA1 _PG_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|A|RB _PG_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_P1|B|1 _PG_01|_SPL_P1|QB1 _PG_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|B|P _PG_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|B|B _PG_01|_SPL_P1|QB1 _PG_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|B|RB _PG_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_PG|I_A1|B _PG_01|_PG|A1 _PG_01|_PG|I_A1|MID  2e-12
I_PG_01|_PG|I_A1|B 0 _PG_01|_PG|I_A1|MID  0.000175
L_PG_01|_PG|I_B1|B _PG_01|_PG|B1 _PG_01|_PG|I_B1|MID  2e-12
I_PG_01|_PG|I_B1|B 0 _PG_01|_PG|I_B1|MID  0.000175
L_PG_01|_PG|I_Q3|B _PG_01|_PG|Q3 _PG_01|_PG|I_Q3|MID  2e-12
I_PG_01|_PG|I_Q3|B 0 _PG_01|_PG|I_Q3|MID  0.00025
L_PG_01|_PG|I_Q2|B _PG_01|_PG|Q2 _PG_01|_PG|I_Q2|MID  2e-12
I_PG_01|_PG|I_Q2|B 0 _PG_01|_PG|I_Q2|MID  0.000175
L_PG_01|_PG|I_Q1|B _PG_01|_PG|Q1 _PG_01|_PG|I_Q1|MID  2e-12
I_PG_01|_PG|I_Q1|B 0 _PG_01|_PG|I_Q1|MID  0.000175
B_PG_01|_PG|A1|1 _PG_01|_PG|A1 _PG_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|A1|P _PG_01|_PG|A1|MID_SERIES 0  2e-13
R_PG_01|_PG|A1|B _PG_01|_PG|A1 _PG_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG_01|_PG|A1|RB _PG_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|A2|1 _PG_01|_PG|A2 _PG_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|A2|P _PG_01|_PG|A2|MID_SERIES 0  2e-13
R_PG_01|_PG|A2|B _PG_01|_PG|A2 _PG_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG_01|_PG|A2|RB _PG_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|A12|1 _PG_01|_PG|A2 _PG_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_PG|A12|B _PG_01|_PG|A2 _PG_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG_01|_PG|A12|RB _PG_01|_PG|A12|MID_SHUNT _PG_01|_PG|A3  2.1704737578552e-12
B_PG_01|_PG|B1|1 _PG_01|_PG|B1 _PG_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|B1|P _PG_01|_PG|B1|MID_SERIES 0  2e-13
R_PG_01|_PG|B1|B _PG_01|_PG|B1 _PG_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG_01|_PG|B1|RB _PG_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|B2|1 _PG_01|_PG|B2 _PG_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|B2|P _PG_01|_PG|B2|MID_SERIES 0  2e-13
R_PG_01|_PG|B2|B _PG_01|_PG|B2 _PG_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG_01|_PG|B2|RB _PG_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|B12|1 _PG_01|_PG|B2 _PG_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_PG|B12|B _PG_01|_PG|B2 _PG_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG_01|_PG|B12|RB _PG_01|_PG|B12|MID_SHUNT _PG_01|_PG|B3  2.1704737578552e-12
B_PG_01|_PG|Q2|1 _PG_01|_PG|Q2 _PG_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|Q2|P _PG_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG_01|_PG|Q2|B _PG_01|_PG|Q2 _PG_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG_01|_PG|Q2|RB _PG_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|Q1|1 _PG_01|_PG|Q1 _PG_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|Q1|P _PG_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG_01|_PG|Q1|B _PG_01|_PG|Q1 _PG_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG_01|_PG|Q1|RB _PG_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_GG|I_A1|B _PG_01|_GG|A1 _PG_01|_GG|I_A1|MID  2e-12
I_PG_01|_GG|I_A1|B 0 _PG_01|_GG|I_A1|MID  0.000175
L_PG_01|_GG|I_B1|B _PG_01|_GG|B1 _PG_01|_GG|I_B1|MID  2e-12
I_PG_01|_GG|I_B1|B 0 _PG_01|_GG|I_B1|MID  0.000175
L_PG_01|_GG|I_Q3|B _PG_01|_GG|Q3 _PG_01|_GG|I_Q3|MID  2e-12
I_PG_01|_GG|I_Q3|B 0 _PG_01|_GG|I_Q3|MID  0.00025
L_PG_01|_GG|I_Q2|B _PG_01|_GG|Q2 _PG_01|_GG|I_Q2|MID  2e-12
I_PG_01|_GG|I_Q2|B 0 _PG_01|_GG|I_Q2|MID  0.000175
L_PG_01|_GG|I_Q1|B _PG_01|_GG|Q1 _PG_01|_GG|I_Q1|MID  2e-12
I_PG_01|_GG|I_Q1|B 0 _PG_01|_GG|I_Q1|MID  0.000175
B_PG_01|_GG|A1|1 _PG_01|_GG|A1 _PG_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|A1|P _PG_01|_GG|A1|MID_SERIES 0  2e-13
R_PG_01|_GG|A1|B _PG_01|_GG|A1 _PG_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG_01|_GG|A1|RB _PG_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|A2|1 _PG_01|_GG|A2 _PG_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|A2|P _PG_01|_GG|A2|MID_SERIES 0  2e-13
R_PG_01|_GG|A2|B _PG_01|_GG|A2 _PG_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG_01|_GG|A2|RB _PG_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|A12|1 _PG_01|_GG|A2 _PG_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_GG|A12|B _PG_01|_GG|A2 _PG_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG_01|_GG|A12|RB _PG_01|_GG|A12|MID_SHUNT _PG_01|_GG|A3  2.1704737578552e-12
B_PG_01|_GG|B1|1 _PG_01|_GG|B1 _PG_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|B1|P _PG_01|_GG|B1|MID_SERIES 0  2e-13
R_PG_01|_GG|B1|B _PG_01|_GG|B1 _PG_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG_01|_GG|B1|RB _PG_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|B2|1 _PG_01|_GG|B2 _PG_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|B2|P _PG_01|_GG|B2|MID_SERIES 0  2e-13
R_PG_01|_GG|B2|B _PG_01|_GG|B2 _PG_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG_01|_GG|B2|RB _PG_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|B12|1 _PG_01|_GG|B2 _PG_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_GG|B12|B _PG_01|_GG|B2 _PG_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG_01|_GG|B12|RB _PG_01|_GG|B12|MID_SHUNT _PG_01|_GG|B3  2.1704737578552e-12
B_PG_01|_GG|Q2|1 _PG_01|_GG|Q2 _PG_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|Q2|P _PG_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG_01|_GG|Q2|B _PG_01|_GG|Q2 _PG_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG_01|_GG|Q2|RB _PG_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|Q1|1 _PG_01|_GG|Q1 _PG_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|Q1|P _PG_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG_01|_GG|Q1|B _PG_01|_GG|Q1 _PG_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG_01|_GG|Q1|RB _PG_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|1|1 _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|1|P _PG_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|1|B _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|1|RB _PG_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|23|1 _PG_01|_DFF_P0|2 _PG_01|_DFF_P0|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P0|23|B _PG_01|_DFF_P0|2 _PG_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P0|23|RB _PG_01|_DFF_P0|23|MID_SHUNT _PG_01|_DFF_P0|3  2.1704737578552e-12
B_PG_01|_DFF_P0|3|1 _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|3|P _PG_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|3|B _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|3|RB _PG_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|4|1 _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|4|P _PG_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|4|B _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|4|RB _PG_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|45|1 _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P0|45|B _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P0|45|RB _PG_01|_DFF_P0|45|MID_SHUNT _PG_01|_DFF_P0|5  2.1704737578552e-12
B_PG_01|_DFF_P0|T|1 _PG_01|_DFF_P0|T1 _PG_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|T|P _PG_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|T|B _PG_01|_DFF_P0|T1 _PG_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|T|RB _PG_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|6|1 _PG_01|_DFF_P0|6 _PG_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|6|P _PG_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|6|B _PG_01|_DFF_P0|6 _PG_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|6|RB _PG_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_P0|I_1|B _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|I_1|MID  2e-12
I_PG_01|_DFF_P0|I_1|B 0 _PG_01|_DFF_P0|I_1|MID  0.000175
L_PG_01|_DFF_P0|I_3|B _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|I_3|MID  2e-12
I_PG_01|_DFF_P0|I_3|B 0 _PG_01|_DFF_P0|I_3|MID  0.00025
L_PG_01|_DFF_P0|I_T|B _PG_01|_DFF_P0|T1 _PG_01|_DFF_P0|I_T|MID  2e-12
I_PG_01|_DFF_P0|I_T|B 0 _PG_01|_DFF_P0|I_T|MID  0.000175
L_PG_01|_DFF_P0|I_6|B _PG_01|_DFF_P0|6 _PG_01|_DFF_P0|I_6|MID  2e-12
I_PG_01|_DFF_P0|I_6|B 0 _PG_01|_DFF_P0|I_6|MID  0.000175
B_PG_01|_DFF_P1|1|1 _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|1|P _PG_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|1|B _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|1|RB _PG_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|23|1 _PG_01|_DFF_P1|2 _PG_01|_DFF_P1|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P1|23|B _PG_01|_DFF_P1|2 _PG_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P1|23|RB _PG_01|_DFF_P1|23|MID_SHUNT _PG_01|_DFF_P1|3  2.1704737578552e-12
B_PG_01|_DFF_P1|3|1 _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|3|P _PG_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|3|B _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|3|RB _PG_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|4|1 _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|4|P _PG_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|4|B _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|4|RB _PG_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|45|1 _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P1|45|B _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P1|45|RB _PG_01|_DFF_P1|45|MID_SHUNT _PG_01|_DFF_P1|5  2.1704737578552e-12
B_PG_01|_DFF_P1|T|1 _PG_01|_DFF_P1|T1 _PG_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|T|P _PG_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|T|B _PG_01|_DFF_P1|T1 _PG_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|T|RB _PG_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|6|1 _PG_01|_DFF_P1|6 _PG_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|6|P _PG_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|6|B _PG_01|_DFF_P1|6 _PG_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|6|RB _PG_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_P1|I_1|B _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|I_1|MID  2e-12
I_PG_01|_DFF_P1|I_1|B 0 _PG_01|_DFF_P1|I_1|MID  0.000175
L_PG_01|_DFF_P1|I_3|B _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|I_3|MID  2e-12
I_PG_01|_DFF_P1|I_3|B 0 _PG_01|_DFF_P1|I_3|MID  0.00025
L_PG_01|_DFF_P1|I_T|B _PG_01|_DFF_P1|T1 _PG_01|_DFF_P1|I_T|MID  2e-12
I_PG_01|_DFF_P1|I_T|B 0 _PG_01|_DFF_P1|I_T|MID  0.000175
L_PG_01|_DFF_P1|I_6|B _PG_01|_DFF_P1|6 _PG_01|_DFF_P1|I_6|MID  2e-12
I_PG_01|_DFF_P1|I_6|B 0 _PG_01|_DFF_P1|I_6|MID  0.000175
B_PG_01|_DFF_PG|1|1 _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|1|P _PG_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|1|B _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|1|RB _PG_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|23|1 _PG_01|_DFF_PG|2 _PG_01|_DFF_PG|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_PG|23|B _PG_01|_DFF_PG|2 _PG_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_PG|23|RB _PG_01|_DFF_PG|23|MID_SHUNT _PG_01|_DFF_PG|3  2.1704737578552e-12
B_PG_01|_DFF_PG|3|1 _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|3|P _PG_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|3|B _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|3|RB _PG_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|4|1 _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|4|P _PG_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|4|B _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|4|RB _PG_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|45|1 _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_PG|45|B _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_PG|45|RB _PG_01|_DFF_PG|45|MID_SHUNT _PG_01|_DFF_PG|5  2.1704737578552e-12
B_PG_01|_DFF_PG|T|1 _PG_01|_DFF_PG|T1 _PG_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|T|P _PG_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|T|B _PG_01|_DFF_PG|T1 _PG_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|T|RB _PG_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|6|1 _PG_01|_DFF_PG|6 _PG_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|6|P _PG_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|6|B _PG_01|_DFF_PG|6 _PG_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|6|RB _PG_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_PG|I_1|B _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|I_1|MID  2e-12
I_PG_01|_DFF_PG|I_1|B 0 _PG_01|_DFF_PG|I_1|MID  0.000175
L_PG_01|_DFF_PG|I_3|B _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|I_3|MID  2e-12
I_PG_01|_DFF_PG|I_3|B 0 _PG_01|_DFF_PG|I_3|MID  0.00025
L_PG_01|_DFF_PG|I_T|B _PG_01|_DFF_PG|T1 _PG_01|_DFF_PG|I_T|MID  2e-12
I_PG_01|_DFF_PG|I_T|B 0 _PG_01|_DFF_PG|I_T|MID  0.000175
L_PG_01|_DFF_PG|I_6|B _PG_01|_DFF_PG|6 _PG_01|_DFF_PG|I_6|MID  2e-12
I_PG_01|_DFF_PG|I_6|B 0 _PG_01|_DFF_PG|I_6|MID  0.000175
B_PG_01|_DFF_GG|1|1 _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|1|P _PG_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|1|B _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|1|RB _PG_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|23|1 _PG_01|_DFF_GG|2 _PG_01|_DFF_GG|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_GG|23|B _PG_01|_DFF_GG|2 _PG_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_GG|23|RB _PG_01|_DFF_GG|23|MID_SHUNT _PG_01|_DFF_GG|3  2.1704737578552e-12
B_PG_01|_DFF_GG|3|1 _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|3|P _PG_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|3|B _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|3|RB _PG_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|4|1 _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|4|P _PG_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|4|B _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|4|RB _PG_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|45|1 _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_GG|45|B _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_GG|45|RB _PG_01|_DFF_GG|45|MID_SHUNT _PG_01|_DFF_GG|5  2.1704737578552e-12
B_PG_01|_DFF_GG|T|1 _PG_01|_DFF_GG|T1 _PG_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|T|P _PG_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|T|B _PG_01|_DFF_GG|T1 _PG_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|T|RB _PG_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|6|1 _PG_01|_DFF_GG|6 _PG_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|6|P _PG_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|6|B _PG_01|_DFF_GG|6 _PG_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|6|RB _PG_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_GG|I_1|B _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|I_1|MID  2e-12
I_PG_01|_DFF_GG|I_1|B 0 _PG_01|_DFF_GG|I_1|MID  0.000175
L_PG_01|_DFF_GG|I_3|B _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|I_3|MID  2e-12
I_PG_01|_DFF_GG|I_3|B 0 _PG_01|_DFF_GG|I_3|MID  0.00025
L_PG_01|_DFF_GG|I_T|B _PG_01|_DFF_GG|T1 _PG_01|_DFF_GG|I_T|MID  2e-12
I_PG_01|_DFF_GG|I_T|B 0 _PG_01|_DFF_GG|I_T|MID  0.000175
L_PG_01|_DFF_GG|I_6|B _PG_01|_DFF_GG|6 _PG_01|_DFF_GG|I_6|MID  2e-12
I_PG_01|_DFF_GG|I_6|B 0 _PG_01|_DFF_GG|I_6|MID  0.000175
L_PG_01|_AND_G|I_A1|B _PG_01|_AND_G|A1 _PG_01|_AND_G|I_A1|MID  2e-12
I_PG_01|_AND_G|I_A1|B 0 _PG_01|_AND_G|I_A1|MID  0.000175
L_PG_01|_AND_G|I_B1|B _PG_01|_AND_G|B1 _PG_01|_AND_G|I_B1|MID  2e-12
I_PG_01|_AND_G|I_B1|B 0 _PG_01|_AND_G|I_B1|MID  0.000175
L_PG_01|_AND_G|I_Q3|B _PG_01|_AND_G|Q3 _PG_01|_AND_G|I_Q3|MID  2e-12
I_PG_01|_AND_G|I_Q3|B 0 _PG_01|_AND_G|I_Q3|MID  7.5e-05
L_PG_01|_AND_G|I_Q2|B _PG_01|_AND_G|Q2 _PG_01|_AND_G|I_Q2|MID  2e-12
I_PG_01|_AND_G|I_Q2|B 0 _PG_01|_AND_G|I_Q2|MID  0.000175
L_PG_01|_AND_G|I_Q1|B _PG_01|_AND_G|Q1 _PG_01|_AND_G|I_Q1|MID  2e-12
I_PG_01|_AND_G|I_Q1|B 0 _PG_01|_AND_G|I_Q1|MID  0.000175
B_PG_01|_AND_G|A1|1 _PG_01|_AND_G|A1 _PG_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|A1|P _PG_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG_01|_AND_G|A1|B _PG_01|_AND_G|A1 _PG_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|A1|RB _PG_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|A2|1 _PG_01|_AND_G|A2 _PG_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|A2|P _PG_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG_01|_AND_G|A2|B _PG_01|_AND_G|A2 _PG_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|A2|RB _PG_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|A12|1 _PG_01|_AND_G|A2 _PG_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_G|A12|B _PG_01|_AND_G|A2 _PG_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG_01|_AND_G|A12|RB _PG_01|_AND_G|A12|MID_SHUNT _PG_01|_AND_G|A3  2.1704737578552e-12
B_PG_01|_AND_G|B1|1 _PG_01|_AND_G|B1 _PG_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|B1|P _PG_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG_01|_AND_G|B1|B _PG_01|_AND_G|B1 _PG_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|B1|RB _PG_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|B2|1 _PG_01|_AND_G|B2 _PG_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|B2|P _PG_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG_01|_AND_G|B2|B _PG_01|_AND_G|B2 _PG_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|B2|RB _PG_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|B12|1 _PG_01|_AND_G|B2 _PG_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_G|B12|B _PG_01|_AND_G|B2 _PG_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG_01|_AND_G|B12|RB _PG_01|_AND_G|B12|MID_SHUNT _PG_01|_AND_G|B3  2.1704737578552e-12
B_PG_01|_AND_G|Q2|1 _PG_01|_AND_G|Q2 _PG_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|Q2|P _PG_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG_01|_AND_G|Q2|B _PG_01|_AND_G|Q2 _PG_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|Q2|RB _PG_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|Q1|1 _PG_01|_AND_G|Q1 _PG_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|Q1|P _PG_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG_01|_AND_G|Q1|B _PG_01|_AND_G|Q1 _PG_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|Q1|RB _PG_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_AND_P|I_A1|B _PG_01|_AND_P|A1 _PG_01|_AND_P|I_A1|MID  2e-12
I_PG_01|_AND_P|I_A1|B 0 _PG_01|_AND_P|I_A1|MID  0.000175
L_PG_01|_AND_P|I_B1|B _PG_01|_AND_P|B1 _PG_01|_AND_P|I_B1|MID  2e-12
I_PG_01|_AND_P|I_B1|B 0 _PG_01|_AND_P|I_B1|MID  0.000175
L_PG_01|_AND_P|I_Q3|B _PG_01|_AND_P|Q3 _PG_01|_AND_P|I_Q3|MID  2e-12
I_PG_01|_AND_P|I_Q3|B 0 _PG_01|_AND_P|I_Q3|MID  7.5e-05
L_PG_01|_AND_P|I_Q2|B _PG_01|_AND_P|Q2 _PG_01|_AND_P|I_Q2|MID  2e-12
I_PG_01|_AND_P|I_Q2|B 0 _PG_01|_AND_P|I_Q2|MID  0.000175
L_PG_01|_AND_P|I_Q1|B _PG_01|_AND_P|Q1 _PG_01|_AND_P|I_Q1|MID  2e-12
I_PG_01|_AND_P|I_Q1|B 0 _PG_01|_AND_P|I_Q1|MID  0.000175
B_PG_01|_AND_P|A1|1 _PG_01|_AND_P|A1 _PG_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|A1|P _PG_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG_01|_AND_P|A1|B _PG_01|_AND_P|A1 _PG_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|A1|RB _PG_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|A2|1 _PG_01|_AND_P|A2 _PG_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|A2|P _PG_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG_01|_AND_P|A2|B _PG_01|_AND_P|A2 _PG_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|A2|RB _PG_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|A12|1 _PG_01|_AND_P|A2 _PG_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_P|A12|B _PG_01|_AND_P|A2 _PG_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG_01|_AND_P|A12|RB _PG_01|_AND_P|A12|MID_SHUNT _PG_01|_AND_P|A3  2.1704737578552e-12
B_PG_01|_AND_P|B1|1 _PG_01|_AND_P|B1 _PG_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|B1|P _PG_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG_01|_AND_P|B1|B _PG_01|_AND_P|B1 _PG_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|B1|RB _PG_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|B2|1 _PG_01|_AND_P|B2 _PG_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|B2|P _PG_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG_01|_AND_P|B2|B _PG_01|_AND_P|B2 _PG_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|B2|RB _PG_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|B12|1 _PG_01|_AND_P|B2 _PG_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_P|B12|B _PG_01|_AND_P|B2 _PG_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG_01|_AND_P|B12|RB _PG_01|_AND_P|B12|MID_SHUNT _PG_01|_AND_P|B3  2.1704737578552e-12
B_PG_01|_AND_P|Q2|1 _PG_01|_AND_P|Q2 _PG_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|Q2|P _PG_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG_01|_AND_P|Q2|B _PG_01|_AND_P|Q2 _PG_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|Q2|RB _PG_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|Q1|1 _PG_01|_AND_P|Q1 _PG_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|Q1|P _PG_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG_01|_AND_P|Q1|B _PG_01|_AND_P|Q1 _PG_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|Q1|RB _PG_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI RS0
.print DEVI RS1
.print DEVI RS2
.print DEVI IT2|T
.print DEVI IT1|T
.print DEVI IT0|T
.print DEVI IDATA_A0|A
.print DEVI IDATA_B0|B
.print DEVI IDATA_A1|C
.print DEVI IDATA_B1|D
.print DEVI L_SPL_P0_0|1
.print DEVI L_SPL_P0_0|2
.print DEVI L_SPL_P0_0|3
.print DEVI L_SPL_P0_0|4
.print DEVI L_SPL_P0_0|5
.print DEVI L_SPL_P0_0|6
.print DEVI L_SPL_P0_0|7
.print DEVI L_SPL_G0_0|1
.print DEVI L_SPL_G0_0|2
.print DEVI L_SPL_G0_0|3
.print DEVI L_SPL_G0_0|4
.print DEVI L_SPL_G0_0|5
.print DEVI L_SPL_G0_0|6
.print DEVI L_SPL_G0_0|7
.print DEVI L_SPL_P1_0|1
.print DEVI L_SPL_P1_0|2
.print DEVI L_SPL_P1_0|3
.print DEVI L_SPL_P1_0|4
.print DEVI L_SPL_P1_0|5
.print DEVI L_SPL_P1_0|6
.print DEVI L_SPL_P1_0|7
.print DEVI L_DFF_P0_01|1
.print DEVI L_DFF_P0_01|2
.print DEVI L_DFF_P0_01|3
.print DEVI L_DFF_P0_01|4
.print DEVI L_DFF_P0_01|T
.print DEVI L_DFF_P0_01|5
.print DEVI L_DFF_P0_01|6
.print DEVI L_DFF_G0_01|1
.print DEVI L_DFF_G0_01|2
.print DEVI L_DFF_G0_01|3
.print DEVI L_DFF_G0_01|4
.print DEVI L_DFF_G0_01|T
.print DEVI L_DFF_G0_01|5
.print DEVI L_DFF_G0_01|6
.print DEVI L_DFF_P1_01|1
.print DEVI L_DFF_P1_01|2
.print DEVI L_DFF_P1_01|3
.print DEVI L_DFF_P1_01|4
.print DEVI L_DFF_P1_01|T
.print DEVI L_DFF_P1_01|5
.print DEVI L_DFF_P1_01|6
.print DEVI L_DFF_S0|1
.print DEVI L_DFF_S0|2
.print DEVI L_DFF_S0|3
.print DEVI L_DFF_S0|4
.print DEVI L_DFF_S0|T
.print DEVI L_DFF_S0|5
.print DEVI L_DFF_S0|6
.print DEVI L_XOR_S1|A1
.print DEVI L_XOR_S1|A2
.print DEVI L_XOR_S1|A3
.print DEVI L_XOR_S1|B1
.print DEVI L_XOR_S1|B2
.print DEVI L_XOR_S1|B3
.print DEVI L_XOR_S1|T1
.print DEVI L_XOR_S1|T2
.print DEVI L_XOR_S1|Q2
.print DEVI L_XOR_S1|Q1
.print DEVI L_DFF_S2|1
.print DEVI L_DFF_S2|2
.print DEVI L_DFF_S2|3
.print DEVI L_DFF_S2|4
.print DEVI L_DFF_S2|T
.print DEVI L_DFF_S2|5
.print DEVI L_DFF_S2|6
.print V _SPL_P1_0|QA1
.print V _DFF_S2|3
.print V _DFF_G0_01|4
.print V _DFF_P0_01|T1
.print V B1I
.print V _DFF_P1_01|2
.print V _DFF_S2|T1
.print V _DFF_P0_01|6
.print V _SPL_P0_0|QB1
.print V _INIT_0|A1_SYNC
.print V _PG_01|G1_COPY_1
.print V G0_1
.print V B0I
.print V _DFF_P1_01|6
.print V _INIT_1|A2
.print V _DFF_P1_01|5
.print V _DFF_S0|2
.print V CLK1
.print V _DFF_S0|5
.print V CLK2
.print V G0_0_W
.print V _XOR_S1|B1
.print V _SPL_P0_0|D1
.print V _PG_01|P1_COPY_1
.print V _DFF_P0_01|2
.print V _XOR_S1|A1
.print V _INIT_0|B1_SYNC
.print V _XOR_S1|AB
.print V _PG_01|P1_SYNC
.print V _PG_01|G1_COPY_2
.print V _SPL_G0_0|JCT
.print V _PG_01|PG_SYNC
.print V _INIT_1|A1
.print V _XOR_S1|T2
.print V _SPL_P0_0|QA1
.print V _DFF_S0|T1
.print V _XOR_S1|ABTQ
.print V P1_0
.print V G1_0
.print V _DFF_P1_01|T1
.print V S0
.print V _PG_01|GG_SYNC
.print V _DFF_G0_01|6
.print V _XOR_S1|B2
.print V _DFF_P0_01|4
.print V _DFF_S2|2
.print V _DFF_S2|6
.print V _PG_01|PG
.print V _XOR_S1|Q1
.print V P0_0
.print V _INIT_0|A1
.print V P0_0_W
.print V _DFF_P1_01|1
.print V _XOR_S1|A2
.print V P1_0_B
.print V _PG_01|P1_COPY_2
.print V A1I
.print V _XOR_S1|A3
.print V _XOR_S1|B3
.print V P0_0_B
.print V _DFF_P0_01|5
.print V _DFF_S2|1
.print V _SPL_P1_0|QB1
.print V _DFF_S0|6
.print V _DFF_G0_01|1
.print V _SPL_G0_0|D2
.print V _DFF_P1_01|3
.print V _DFF_P1_01|4
.print V _DFF_G0_01|3
.print V _PG_01|GG
.print V _SPL_P1_0|D1
.print V _XOR_S1|T1
.print V _INIT_1|B2
.print V _SPL_P0_0|D2
.print V _SPL_P1_0|D2
.print V P1_1
.print V _SPL_G0_0|QA1
.print V _DFF_S0|1
.print V _DFF_S2|4
.print V G0_0
.print V _SPL_G0_0|QB1
.print V _DFF_S2|5
.print V CLK0
.print V P1_0_W
.print V _INIT_0|A2
.print V _DFF_P0_01|1
.print V G1_1
.print V A0I
.print V S1
.print V _DFF_G0_01|T1
.print V _DFF_S0|4
.print V _SPL_G0_0|D1
.print V _INIT_1|B1_SYNC
.print V _INIT_0|B2
.print V _INIT_1|B1
.print V G0_0_B
.print V _SPL_P1_0|JCT
.print V _DFF_S0|3
.print V S2
.print V _PG_01|P0_SYNC
.print V _INIT_0|B1
.print V _DFF_G0_01|2
.print V _DFF_G0_01|5
.print V _INIT_1|A1_SYNC
.print V _SPL_P0_0|JCT
.print V _DFF_P0_01|3
.print V P0_1
