*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OS=1e-11
.PARAM TCLOCK=1e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.25E-12 21E-10
RS0 S0 0  1
RS1 S1 0  1
RIG1 IG1_1 0  1
RS2 S2 0  1
RP1 P1_1 0  1
RG1 G1_1 0  1
IDATA_A0|A 0 A0  PWL(0 0 1.17e-10 0 1.2e-10 0.0005 1.23e-10 0 3.17e-10 0 3.2e-10 0.0005 3.23e-10 0 5.17e-10 0 5.2e-10 0.0005 5.23e-10 0 7.17e-10 0 7.2e-10 0.0005 7.23e-10 0 9.17e-10 0 9.2e-10 0.0005 9.23e-10 0 1.117e-09 0 1.12e-09 0.0005 1.123e-09 0 1.317e-09 0 1.32e-09 0.0005 1.323e-09 0 1.517e-09 0 1.52e-09 0.0005 1.523e-09 0 1.717e-09 0 1.72e-09 0.0005 1.723e-09 0 1.917e-09 0 1.92e-09 0.0005 1.923e-09 0 2.117e-09 0 2.12e-09 0.0005 2.123e-09 0 2.317e-09 0 2.32e-09 0.0005 2.323e-09 0 2.517e-09 0 2.52e-09 0.0005 2.523e-09 0 2.717e-09 0 2.72e-09 0.0005 2.723e-09 0 2.917e-09 0 2.92e-09 0.0005 2.923e-09 0 3.117e-09 0 3.12e-09 0.0005 3.123e-09 0 3.317e-09 0 3.32e-09 0.0005 3.323e-09 0 3.517e-09 0 3.52e-09 0.0005 3.523e-09 0 3.717e-09 0 3.72e-09 0.0005 3.723e-09 0)
IDATA_B0|B 0 B0  PWL(0 0 2.37e-10 0 2.4e-10 0.0005 2.43e-10 0 3.37e-10 0 3.4e-10 0.0005 3.43e-10 0 6.37e-10 0 6.4e-10 0.0005 6.43e-10 0 7.37e-10 0 7.4e-10 0.0005 7.43e-10 0 1.037e-09 0 1.04e-09 0.0005 1.043e-09 0 1.137e-09 0 1.14e-09 0.0005 1.143e-09 0 1.437e-09 0 1.44e-09 0.0005 1.443e-09 0 1.537e-09 0 1.54e-09 0.0005 1.543e-09 0 1.837e-09 0 1.84e-09 0.0005 1.843e-09 0 1.937e-09 0 1.94e-09 0.0005 1.943e-09 0 2.237e-09 0 2.24e-09 0.0005 2.243e-09 0 2.337e-09 0 2.34e-09 0.0005 2.343e-09 0 2.637e-09 0 2.64e-09 0.0005 2.643e-09 0 2.737e-09 0 2.74e-09 0.0005 2.743e-09 0 3.037e-09 0 3.04e-09 0.0005 3.043e-09 0 3.137e-09 0 3.14e-09 0.0005 3.143e-09 0 3.437e-09 0 3.44e-09 0.0005 3.443e-09 0 3.537e-09 0 3.54e-09 0.0005 3.543e-09 0 3.837e-09 0 3.84e-09 0.0005 3.843e-09 0)
IDATA_A1|C 0 A1  PWL(0 0 4.57e-10 0 4.6e-10 0.0005 4.63e-10 0 5.57e-10 0 5.6e-10 0.0005 5.63e-10 0 6.57e-10 0 6.6e-10 0.0005 6.63e-10 0 7.57e-10 0 7.6e-10 0.0005 7.63e-10 0 1.257e-09 0 1.26e-09 0.0005 1.263e-09 0 1.357e-09 0 1.36e-09 0.0005 1.363e-09 0 1.457e-09 0 1.46e-09 0.0005 1.463e-09 0 1.557e-09 0 1.56e-09 0.0005 1.563e-09 0 2.057e-09 0 2.06e-09 0.0005 2.063e-09 0 2.157e-09 0 2.16e-09 0.0005 2.163e-09 0 2.257e-09 0 2.26e-09 0.0005 2.263e-09 0 2.357e-09 0 2.36e-09 0.0005 2.363e-09 0 2.857e-09 0 2.86e-09 0.0005 2.863e-09 0 2.957e-09 0 2.96e-09 0.0005 2.963e-09 0 3.057e-09 0 3.06e-09 0.0005 3.063e-09 0 3.157e-09 0 3.16e-09 0.0005 3.163e-09 0 3.657e-09 0 3.66e-09 0.0005 3.663e-09 0 3.757e-09 0 3.76e-09 0.0005 3.763e-09 0 3.857e-09 0 3.86e-09 0.0005 3.863e-09 0)
IDATA_B1|D 0 B1  PWL(0 0 8.77e-10 0 8.8e-10 0.0005 8.83e-10 0 9.77e-10 0 9.8e-10 0.0005 9.83e-10 0 1.077e-09 0 1.08e-09 0.0005 1.083e-09 0 1.177e-09 0 1.18e-09 0.0005 1.183e-09 0 1.277e-09 0 1.28e-09 0.0005 1.283e-09 0 1.377e-09 0 1.38e-09 0.0005 1.383e-09 0 1.477e-09 0 1.48e-09 0.0005 1.483e-09 0 1.577e-09 0 1.58e-09 0.0005 1.583e-09 0 2.477e-09 0 2.48e-09 0.0005 2.483e-09 0 2.577e-09 0 2.58e-09 0.0005 2.583e-09 0 2.677e-09 0 2.68e-09 0.0005 2.683e-09 0 2.777e-09 0 2.78e-09 0.0005 2.783e-09 0 2.877e-09 0 2.88e-09 0.0005 2.883e-09 0 2.977e-09 0 2.98e-09 0.0005 2.983e-09 0 3.077e-09 0 3.08e-09 0.0005 3.083e-09 0 3.177e-09 0 3.18e-09 0.0005 3.183e-09 0)
IT1|T 0 CLK1  PWL(0 0 7e-12 0 1e-11 0.0015 1.3e-11 0 1.07e-10 0 1.1e-10 0.0015 1.13e-10 0 2.07e-10 0 2.1e-10 0.0015 2.13e-10 0 3.07e-10 0 3.1e-10 0.0015 3.13e-10 0 4.07e-10 0 4.1e-10 0.0015 4.13e-10 0 5.07e-10 0 5.1e-10 0.0015 5.13e-10 0 6.07e-10 0 6.1e-10 0.0015 6.13e-10 0 7.07e-10 0 7.1e-10 0.0015 7.13e-10 0 8.07e-10 0 8.1e-10 0.0015 8.13e-10 0 9.07e-10 0 9.1e-10 0.0015 9.13e-10 0 1.007e-09 0 1.01e-09 0.0015 1.013e-09 0 1.107e-09 0 1.11e-09 0.0015 1.113e-09 0 1.207e-09 0 1.21e-09 0.0015 1.213e-09 0 1.307e-09 0 1.31e-09 0.0015 1.313e-09 0 1.407e-09 0 1.41e-09 0.0015 1.413e-09 0 1.507e-09 0 1.51e-09 0.0015 1.513e-09 0 1.607e-09 0 1.61e-09 0.0015 1.613e-09 0 1.707e-09 0 1.71e-09 0.0015 1.713e-09 0 1.807e-09 0 1.81e-09 0.0015 1.813e-09 0 1.907e-09 0 1.91e-09 0.0015 1.913e-09 0 2.007e-09 0 2.01e-09 0.0015 2.013e-09 0 2.107e-09 0 2.11e-09 0.0015 2.113e-09 0 2.207e-09 0 2.21e-09 0.0015 2.213e-09 0 2.307e-09 0 2.31e-09 0.0015 2.313e-09 0 2.407e-09 0 2.41e-09 0.0015 2.413e-09 0 2.507e-09 0 2.51e-09 0.0015 2.513e-09 0 2.607e-09 0 2.61e-09 0.0015 2.613e-09 0 2.707e-09 0 2.71e-09 0.0015 2.713e-09 0 2.807e-09 0 2.81e-09 0.0015 2.813e-09 0 2.907e-09 0 2.91e-09 0.0015 2.913e-09 0 3.007e-09 0 3.01e-09 0.0015 3.013e-09 0 3.107e-09 0 3.11e-09 0.0015 3.113e-09 0 3.207e-09 0 3.21e-09 0.0015 3.213e-09 0 3.307e-09 0 3.31e-09 0.0015 3.313e-09 0 3.407e-09 0 3.41e-09 0.0015 3.413e-09 0 3.507e-09 0 3.51e-09 0.0015 3.513e-09 0 3.607e-09 0 3.61e-09 0.0015 3.613e-09 0 3.707e-09 0 3.71e-09 0.0015 3.713e-09 0 3.807e-09 0 3.81e-09 0.0015 3.813e-09 0)
IT2|T 0 CLK2  PWL(0 0 7e-12 0 1e-11 0.0015 1.3e-11 0 1.07e-10 0 1.1e-10 0.0015 1.13e-10 0 2.07e-10 0 2.1e-10 0.0015 2.13e-10 0 3.07e-10 0 3.1e-10 0.0015 3.13e-10 0 4.07e-10 0 4.1e-10 0.0015 4.13e-10 0 5.07e-10 0 5.1e-10 0.0015 5.13e-10 0 6.07e-10 0 6.1e-10 0.0015 6.13e-10 0 7.07e-10 0 7.1e-10 0.0015 7.13e-10 0 8.07e-10 0 8.1e-10 0.0015 8.13e-10 0 9.07e-10 0 9.1e-10 0.0015 9.13e-10 0 1.007e-09 0 1.01e-09 0.0015 1.013e-09 0 1.107e-09 0 1.11e-09 0.0015 1.113e-09 0 1.207e-09 0 1.21e-09 0.0015 1.213e-09 0 1.307e-09 0 1.31e-09 0.0015 1.313e-09 0 1.407e-09 0 1.41e-09 0.0015 1.413e-09 0 1.507e-09 0 1.51e-09 0.0015 1.513e-09 0 1.607e-09 0 1.61e-09 0.0015 1.613e-09 0 1.707e-09 0 1.71e-09 0.0015 1.713e-09 0 1.807e-09 0 1.81e-09 0.0015 1.813e-09 0 1.907e-09 0 1.91e-09 0.0015 1.913e-09 0 2.007e-09 0 2.01e-09 0.0015 2.013e-09 0 2.107e-09 0 2.11e-09 0.0015 2.113e-09 0 2.207e-09 0 2.21e-09 0.0015 2.213e-09 0 2.307e-09 0 2.31e-09 0.0015 2.313e-09 0 2.407e-09 0 2.41e-09 0.0015 2.413e-09 0 2.507e-09 0 2.51e-09 0.0015 2.513e-09 0 2.607e-09 0 2.61e-09 0.0015 2.613e-09 0 2.707e-09 0 2.71e-09 0.0015 2.713e-09 0 2.807e-09 0 2.81e-09 0.0015 2.813e-09 0 2.907e-09 0 2.91e-09 0.0015 2.913e-09 0 3.007e-09 0 3.01e-09 0.0015 3.013e-09 0 3.107e-09 0 3.11e-09 0.0015 3.113e-09 0 3.207e-09 0 3.21e-09 0.0015 3.213e-09 0 3.307e-09 0 3.31e-09 0.0015 3.313e-09 0 3.407e-09 0 3.41e-09 0.0015 3.413e-09 0 3.507e-09 0 3.51e-09 0.0015 3.513e-09 0 3.607e-09 0 3.61e-09 0.0015 3.613e-09 0 3.707e-09 0 3.71e-09 0.0015 3.713e-09 0 3.807e-09 0 3.81e-09 0.0015 3.813e-09 0)
L_SPL_P0|1 IP0_0 _SPL_P0|D1  2e-12
L_SPL_P0|2 _SPL_P0|D1 _SPL_P0|D2  4.135667696e-12
L_SPL_P0|3 _SPL_P0|D2 _SPL_P0|JCT  1.4770241771428573e-12
L_SPL_P0|4 _SPL_P0|JCT _SPL_P0|QA1  1.4770241771428573e-12
L_SPL_P0|5 _SPL_P0|QA1 IP0_0_B  2e-12
L_SPL_P0|6 _SPL_P0|JCT _SPL_P0|QB1  1.4770241771428573e-12
L_SPL_P0|7 _SPL_P0|QB1 IP0_0_W  2e-12
L_SPL_G0|1 IG0_0 _SPL_G0|D1  2e-12
L_SPL_G0|2 _SPL_G0|D1 _SPL_G0|D2  4.135667696e-12
L_SPL_G0|3 _SPL_G0|D2 _SPL_G0|JCT  1.4770241771428573e-12
L_SPL_G0|4 _SPL_G0|JCT _SPL_G0|QA1  1.4770241771428573e-12
L_SPL_G0|5 _SPL_G0|QA1 IG0_0_B  2e-12
L_SPL_G0|6 _SPL_G0|JCT _SPL_G0|QB1  1.4770241771428573e-12
L_SPL_G0|7 _SPL_G0|QB1 IG0_0_W  2e-12
L_SPL_P1|1 IP1_0 _SPL_P1|D1  2e-12
L_SPL_P1|2 _SPL_P1|D1 _SPL_P1|D2  4.135667696e-12
L_SPL_P1|3 _SPL_P1|D2 _SPL_P1|JCT  1.4770241771428573e-12
L_SPL_P1|4 _SPL_P1|JCT _SPL_P1|QA1  1.4770241771428573e-12
L_SPL_P1|5 _SPL_P1|QA1 IP1_0_B  2e-12
L_SPL_P1|6 _SPL_P1|JCT _SPL_P1|QB1  1.4770241771428573e-12
L_SPL_P1|7 _SPL_P1|QB1 IP1_0_W  2e-12
L_SPL_G1|1 IG1_0 _SPL_G1|D1  2e-12
L_SPL_G1|2 _SPL_G1|D1 _SPL_G1|D2  4.135667696e-12
L_SPL_G1|3 _SPL_G1|D2 _SPL_G1|JCT  1.4770241771428573e-12
L_SPL_G1|4 _SPL_G1|JCT _SPL_G1|QA1  1.4770241771428573e-12
L_SPL_G1|5 _SPL_G1|QA1 IG1_0_B  2e-12
L_SPL_G1|6 _SPL_G1|JCT _SPL_G1|QB1  1.4770241771428573e-12
L_SPL_G1|7 _SPL_G1|QB1 IG1_0_W  2e-12
IT3|T 0 CLK3  PWL(0 0 -3e-12 0 0 0.002 3e-12 0 9.7e-11 0 1e-10 0.002 1.03e-10 0 1.97e-10 0 2e-10 0.002 2.03e-10 0 2.97e-10 0 3e-10 0.002 3.03e-10 0 3.97e-10 0 4e-10 0.002 4.03e-10 0 4.97e-10 0 5e-10 0.002 5.03e-10 0 5.97e-10 0 6e-10 0.002 6.03e-10 0 6.97e-10 0 7e-10 0.002 7.03e-10 0 7.97e-10 0 8e-10 0.002 8.03e-10 0 8.97e-10 0 9e-10 0.002 9.03e-10 0 9.97e-10 0 1e-09 0.002 1.003e-09 0 1.097e-09 0 1.1e-09 0.002 1.103e-09 0 1.197e-09 0 1.2e-09 0.002 1.203e-09 0 1.297e-09 0 1.3e-09 0.002 1.303e-09 0 1.397e-09 0 1.4e-09 0.002 1.403e-09 0 1.497e-09 0 1.5e-09 0.002 1.503e-09 0 1.597e-09 0 1.6e-09 0.002 1.603e-09 0 1.697e-09 0 1.7e-09 0.002 1.703e-09 0 1.797e-09 0 1.8e-09 0.002 1.803e-09 0 1.897e-09 0 1.9e-09 0.002 1.903e-09 0 1.997e-09 0 2e-09 0.002 2.003e-09 0 2.097e-09 0 2.1e-09 0.002 2.103e-09 0 2.197e-09 0 2.2e-09 0.002 2.203e-09 0 2.297e-09 0 2.3e-09 0.002 2.303e-09 0 2.397e-09 0 2.4e-09 0.002 2.403e-09 0 2.497e-09 0 2.5e-09 0.002 2.503e-09 0 2.597e-09 0 2.6e-09 0.002 2.603e-09 0 2.697e-09 0 2.7e-09 0.002 2.703e-09 0 2.797e-09 0 2.8e-09 0.002 2.803e-09 0 2.897e-09 0 2.9e-09 0.002 2.903e-09 0 2.997e-09 0 3e-09 0.002 3.003e-09 0 3.097e-09 0 3.1e-09 0.002 3.103e-09 0 3.197e-09 0 3.2e-09 0.002 3.203e-09 0 3.297e-09 0 3.3e-09 0.002 3.303e-09 0 3.397e-09 0 3.4e-09 0.002 3.403e-09 0 3.497e-09 0 3.5e-09 0.002 3.503e-09 0 3.597e-09 0 3.6e-09 0.002 3.603e-09 0 3.697e-09 0 3.7e-09 0.002 3.703e-09 0 3.797e-09 0 3.8e-09 0.002 3.803e-09 0)
IT4|T 0 CLK4  PWL(0 0 -3e-12 0 0 0.0005 3e-12 0 9.7e-11 0 1e-10 0.0005 1.03e-10 0 1.97e-10 0 2e-10 0.0005 2.03e-10 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 3.97e-10 0 4e-10 0.0005 4.03e-10 0 4.97e-10 0 5e-10 0.0005 5.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 6.97e-10 0 7e-10 0.0005 7.03e-10 0 7.97e-10 0 8e-10 0.0005 8.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 9.97e-10 0 1e-09 0.0005 1.003e-09 0 1.097e-09 0 1.1e-09 0.0005 1.103e-09 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.297e-09 0 1.3e-09 0.0005 1.303e-09 0 1.397e-09 0 1.4e-09 0.0005 1.403e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.597e-09 0 1.6e-09 0.0005 1.603e-09 0 1.697e-09 0 1.7e-09 0.0005 1.703e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 1.897e-09 0 1.9e-09 0.0005 1.903e-09 0 1.997e-09 0 2e-09 0.0005 2.003e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.197e-09 0 2.2e-09 0.0005 2.203e-09 0 2.297e-09 0 2.3e-09 0.0005 2.303e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.497e-09 0 2.5e-09 0.0005 2.503e-09 0 2.597e-09 0 2.6e-09 0.0005 2.603e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.797e-09 0 2.8e-09 0.0005 2.803e-09 0 2.897e-09 0 2.9e-09 0.0005 2.903e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.097e-09 0 3.1e-09 0.0005 3.103e-09 0 3.197e-09 0 3.2e-09 0.0005 3.203e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.397e-09 0 3.4e-09 0.0005 3.403e-09 0 3.497e-09 0 3.5e-09 0.0005 3.503e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.697e-09 0 3.7e-09 0.0005 3.703e-09 0 3.797e-09 0 3.8e-09 0.0005 3.803e-09 0)
L_DFF_IP0_01|1 IP0_0_W _DFF_IP0_01|1  2.067833848e-12
L_DFF_IP0_01|2 _DFF_IP0_01|1 _DFF_IP0_01|2  4.135667696e-12
L_DFF_IP0_01|3 _DFF_IP0_01|3 _DFF_IP0_01|4  8.271335392e-12
L_DFF_IP0_01|4 _DFF_IP0_01|5 _DFF_IP0_01|T1  4.135667696e-12
L_DFF_IP0_01|T CLK4 _DFF_IP0_01|T1  2.067833848e-12
L_DFF_IP0_01|5 _DFF_IP0_01|4 _DFF_IP0_01|6  4.135667696e-12
L_DFF_IP0_01|6 _DFF_IP0_01|6 IP0_1  2.067833848e-12
IT5|T 0 CLK5  PWL(0 0 -1.3e-11 0 -1e-11 0.0005 -7e-12 0 8.7e-11 0 9e-11 0.0005 9.3e-11 0 1.87e-10 0 1.9e-10 0.0005 1.93e-10 0 2.87e-10 0 2.9e-10 0.0005 2.93e-10 0 3.87e-10 0 3.9e-10 0.0005 3.93e-10 0 4.87e-10 0 4.9e-10 0.0005 4.93e-10 0 5.87e-10 0 5.9e-10 0.0005 5.93e-10 0 6.87e-10 0 6.9e-10 0.0005 6.93e-10 0 7.87e-10 0 7.9e-10 0.0005 7.93e-10 0 8.87e-10 0 8.9e-10 0.0005 8.93e-10 0 9.87e-10 0 9.9e-10 0.0005 9.93e-10 0 1.087e-09 0 1.09e-09 0.0005 1.093e-09 0 1.187e-09 0 1.19e-09 0.0005 1.193e-09 0 1.287e-09 0 1.29e-09 0.0005 1.293e-09 0 1.387e-09 0 1.39e-09 0.0005 1.393e-09 0 1.487e-09 0 1.49e-09 0.0005 1.493e-09 0 1.587e-09 0 1.59e-09 0.0005 1.593e-09 0 1.687e-09 0 1.69e-09 0.0005 1.693e-09 0 1.787e-09 0 1.79e-09 0.0005 1.793e-09 0 1.887e-09 0 1.89e-09 0.0005 1.893e-09 0 1.987e-09 0 1.99e-09 0.0005 1.993e-09 0 2.087e-09 0 2.09e-09 0.0005 2.093e-09 0 2.187e-09 0 2.19e-09 0.0005 2.193e-09 0 2.287e-09 0 2.29e-09 0.0005 2.293e-09 0 2.387e-09 0 2.39e-09 0.0005 2.393e-09 0 2.487e-09 0 2.49e-09 0.0005 2.493e-09 0 2.587e-09 0 2.59e-09 0.0005 2.593e-09 0 2.687e-09 0 2.69e-09 0.0005 2.693e-09 0 2.787e-09 0 2.79e-09 0.0005 2.793e-09 0 2.887e-09 0 2.89e-09 0.0005 2.893e-09 0 2.987e-09 0 2.99e-09 0.0005 2.993e-09 0 3.087e-09 0 3.09e-09 0.0005 3.093e-09 0 3.187e-09 0 3.19e-09 0.0005 3.193e-09 0 3.287e-09 0 3.29e-09 0.0005 3.293e-09 0 3.387e-09 0 3.39e-09 0.0005 3.393e-09 0 3.487e-09 0 3.49e-09 0.0005 3.493e-09 0 3.587e-09 0 3.59e-09 0.0005 3.593e-09 0 3.687e-09 0 3.69e-09 0.0005 3.693e-09 0 3.787e-09 0 3.79e-09 0.0005 3.793e-09 0)
L_DFF_IP0_12|1 IP0_1 _DFF_IP0_12|1  2.067833848e-12
L_DFF_IP0_12|2 _DFF_IP0_12|1 _DFF_IP0_12|2  4.135667696e-12
L_DFF_IP0_12|3 _DFF_IP0_12|3 _DFF_IP0_12|4  8.271335392e-12
L_DFF_IP0_12|4 _DFF_IP0_12|5 _DFF_IP0_12|T1  4.135667696e-12
L_DFF_IP0_12|T CLK5 _DFF_IP0_12|T1  2.067833848e-12
L_DFF_IP0_12|5 _DFF_IP0_12|4 _DFF_IP0_12|6  4.135667696e-12
L_DFF_IP0_12|6 _DFF_IP0_12|6 S0  2.067833848e-12
IT6|T 0 CLK6  PWL(0 0 -3e-12 0 0 0.0005 3e-12 0 9.7e-11 0 1e-10 0.0005 1.03e-10 0 1.97e-10 0 2e-10 0.0005 2.03e-10 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 3.97e-10 0 4e-10 0.0005 4.03e-10 0 4.97e-10 0 5e-10 0.0005 5.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 6.97e-10 0 7e-10 0.0005 7.03e-10 0 7.97e-10 0 8e-10 0.0005 8.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 9.97e-10 0 1e-09 0.0005 1.003e-09 0 1.097e-09 0 1.1e-09 0.0005 1.103e-09 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.297e-09 0 1.3e-09 0.0005 1.303e-09 0 1.397e-09 0 1.4e-09 0.0005 1.403e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.597e-09 0 1.6e-09 0.0005 1.603e-09 0 1.697e-09 0 1.7e-09 0.0005 1.703e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 1.897e-09 0 1.9e-09 0.0005 1.903e-09 0 1.997e-09 0 2e-09 0.0005 2.003e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.197e-09 0 2.2e-09 0.0005 2.203e-09 0 2.297e-09 0 2.3e-09 0.0005 2.303e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.497e-09 0 2.5e-09 0.0005 2.503e-09 0 2.597e-09 0 2.6e-09 0.0005 2.603e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.797e-09 0 2.8e-09 0.0005 2.803e-09 0 2.897e-09 0 2.9e-09 0.0005 2.903e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.097e-09 0 3.1e-09 0.0005 3.103e-09 0 3.197e-09 0 3.2e-09 0.0005 3.203e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.397e-09 0 3.4e-09 0.0005 3.403e-09 0 3.497e-09 0 3.5e-09 0.0005 3.503e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.697e-09 0 3.7e-09 0.0005 3.703e-09 0 3.797e-09 0 3.8e-09 0.0005 3.803e-09 0)
L_DFF_IG0_01|1 IG0_0_W _DFF_IG0_01|1  2.067833848e-12
L_DFF_IG0_01|2 _DFF_IG0_01|1 _DFF_IG0_01|2  4.135667696e-12
L_DFF_IG0_01|3 _DFF_IG0_01|3 _DFF_IG0_01|4  8.271335392e-12
L_DFF_IG0_01|4 _DFF_IG0_01|5 _DFF_IG0_01|T1  4.135667696e-12
L_DFF_IG0_01|T CLK6 _DFF_IG0_01|T1  2.067833848e-12
L_DFF_IG0_01|5 _DFF_IG0_01|4 _DFF_IG0_01|6  4.135667696e-12
L_DFF_IG0_01|6 _DFF_IG0_01|6 IG0_1  2.067833848e-12
IT7|T 0 CLK7  PWL(0 0 -3e-12 0 0 0.0005 3e-12 0 9.7e-11 0 1e-10 0.0005 1.03e-10 0 1.97e-10 0 2e-10 0.0005 2.03e-10 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 3.97e-10 0 4e-10 0.0005 4.03e-10 0 4.97e-10 0 5e-10 0.0005 5.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 6.97e-10 0 7e-10 0.0005 7.03e-10 0 7.97e-10 0 8e-10 0.0005 8.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 9.97e-10 0 1e-09 0.0005 1.003e-09 0 1.097e-09 0 1.1e-09 0.0005 1.103e-09 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.297e-09 0 1.3e-09 0.0005 1.303e-09 0 1.397e-09 0 1.4e-09 0.0005 1.403e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.597e-09 0 1.6e-09 0.0005 1.603e-09 0 1.697e-09 0 1.7e-09 0.0005 1.703e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 1.897e-09 0 1.9e-09 0.0005 1.903e-09 0 1.997e-09 0 2e-09 0.0005 2.003e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.197e-09 0 2.2e-09 0.0005 2.203e-09 0 2.297e-09 0 2.3e-09 0.0005 2.303e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.497e-09 0 2.5e-09 0.0005 2.503e-09 0 2.597e-09 0 2.6e-09 0.0005 2.603e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.797e-09 0 2.8e-09 0.0005 2.803e-09 0 2.897e-09 0 2.9e-09 0.0005 2.903e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.097e-09 0 3.1e-09 0.0005 3.103e-09 0 3.197e-09 0 3.2e-09 0.0005 3.203e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.397e-09 0 3.4e-09 0.0005 3.403e-09 0 3.497e-09 0 3.5e-09 0.0005 3.503e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.697e-09 0 3.7e-09 0.0005 3.703e-09 0 3.797e-09 0 3.8e-09 0.0005 3.803e-09 0)
L_DFF_IP1_01|1 IP1_0_W _DFF_IP1_01|1  2.067833848e-12
L_DFF_IP1_01|2 _DFF_IP1_01|1 _DFF_IP1_01|2  4.135667696e-12
L_DFF_IP1_01|3 _DFF_IP1_01|3 _DFF_IP1_01|4  8.271335392e-12
L_DFF_IP1_01|4 _DFF_IP1_01|5 _DFF_IP1_01|T1  4.135667696e-12
L_DFF_IP1_01|T CLK7 _DFF_IP1_01|T1  2.067833848e-12
L_DFF_IP1_01|5 _DFF_IP1_01|4 _DFF_IP1_01|6  4.135667696e-12
L_DFF_IP1_01|6 _DFF_IP1_01|6 IP1_1  2.067833848e-12
IT8|T 0 CLK8  PWL(0 0 -1.3e-11 0 -1e-11 0.0005 -7e-12 0 8.7e-11 0 9e-11 0.0005 9.3e-11 0 1.87e-10 0 1.9e-10 0.0005 1.93e-10 0 2.87e-10 0 2.9e-10 0.0005 2.93e-10 0 3.87e-10 0 3.9e-10 0.0005 3.93e-10 0 4.87e-10 0 4.9e-10 0.0005 4.93e-10 0 5.87e-10 0 5.9e-10 0.0005 5.93e-10 0 6.87e-10 0 6.9e-10 0.0005 6.93e-10 0 7.87e-10 0 7.9e-10 0.0005 7.93e-10 0 8.87e-10 0 8.9e-10 0.0005 8.93e-10 0 9.87e-10 0 9.9e-10 0.0005 9.93e-10 0 1.087e-09 0 1.09e-09 0.0005 1.093e-09 0 1.187e-09 0 1.19e-09 0.0005 1.193e-09 0 1.287e-09 0 1.29e-09 0.0005 1.293e-09 0 1.387e-09 0 1.39e-09 0.0005 1.393e-09 0 1.487e-09 0 1.49e-09 0.0005 1.493e-09 0 1.587e-09 0 1.59e-09 0.0005 1.593e-09 0 1.687e-09 0 1.69e-09 0.0005 1.693e-09 0 1.787e-09 0 1.79e-09 0.0005 1.793e-09 0 1.887e-09 0 1.89e-09 0.0005 1.893e-09 0 1.987e-09 0 1.99e-09 0.0005 1.993e-09 0 2.087e-09 0 2.09e-09 0.0005 2.093e-09 0 2.187e-09 0 2.19e-09 0.0005 2.193e-09 0 2.287e-09 0 2.29e-09 0.0005 2.293e-09 0 2.387e-09 0 2.39e-09 0.0005 2.393e-09 0 2.487e-09 0 2.49e-09 0.0005 2.493e-09 0 2.587e-09 0 2.59e-09 0.0005 2.593e-09 0 2.687e-09 0 2.69e-09 0.0005 2.693e-09 0 2.787e-09 0 2.79e-09 0.0005 2.793e-09 0 2.887e-09 0 2.89e-09 0.0005 2.893e-09 0 2.987e-09 0 2.99e-09 0.0005 2.993e-09 0 3.087e-09 0 3.09e-09 0.0005 3.093e-09 0 3.187e-09 0 3.19e-09 0.0005 3.193e-09 0 3.287e-09 0 3.29e-09 0.0005 3.293e-09 0 3.387e-09 0 3.39e-09 0.0005 3.393e-09 0 3.487e-09 0 3.49e-09 0.0005 3.493e-09 0 3.587e-09 0 3.59e-09 0.0005 3.593e-09 0 3.687e-09 0 3.69e-09 0.0005 3.693e-09 0 3.787e-09 0 3.79e-09 0.0005 3.793e-09 0)
L_XOR_S1|A1 IG0_1 _XOR_S1|A1  2.067833848e-12
L_XOR_S1|A2 _XOR_S1|A1 _XOR_S1|A2  4.135667696e-12
L_XOR_S1|A3 _XOR_S1|A3 _XOR_S1|AB  8.271335392e-12
L_XOR_S1|B1 IP1_1 _XOR_S1|B1  2.067833848e-12
L_XOR_S1|B2 _XOR_S1|B1 _XOR_S1|B2  4.135667696e-12
L_XOR_S1|B3 _XOR_S1|B3 _XOR_S1|AB  8.271335392e-12
L_XOR_S1|T1 CLK8 _XOR_S1|T1  2.067833848e-12
L_XOR_S1|T2 _XOR_S1|T1 _XOR_S1|T2  4.135667696e-12
L_XOR_S1|Q2 _XOR_S1|ABTQ _XOR_S1|Q1  4.135667696e-12
L_XOR_S1|Q1 _XOR_S1|Q1 S1  2.067833848e-12
IT9|T 0 CLK9  PWL(0 0 -3e-12 0 0 0.0005 3e-12 0 9.7e-11 0 1e-10 0.0005 1.03e-10 0 1.97e-10 0 2e-10 0.0005 2.03e-10 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 3.97e-10 0 4e-10 0.0005 4.03e-10 0 4.97e-10 0 5e-10 0.0005 5.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 6.97e-10 0 7e-10 0.0005 7.03e-10 0 7.97e-10 0 8e-10 0.0005 8.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 9.97e-10 0 1e-09 0.0005 1.003e-09 0 1.097e-09 0 1.1e-09 0.0005 1.103e-09 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.297e-09 0 1.3e-09 0.0005 1.303e-09 0 1.397e-09 0 1.4e-09 0.0005 1.403e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.597e-09 0 1.6e-09 0.0005 1.603e-09 0 1.697e-09 0 1.7e-09 0.0005 1.703e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 1.897e-09 0 1.9e-09 0.0005 1.903e-09 0 1.997e-09 0 2e-09 0.0005 2.003e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.197e-09 0 2.2e-09 0.0005 2.203e-09 0 2.297e-09 0 2.3e-09 0.0005 2.303e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.497e-09 0 2.5e-09 0.0005 2.503e-09 0 2.597e-09 0 2.6e-09 0.0005 2.603e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.797e-09 0 2.8e-09 0.0005 2.803e-09 0 2.897e-09 0 2.9e-09 0.0005 2.903e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.097e-09 0 3.1e-09 0.0005 3.103e-09 0 3.197e-09 0 3.2e-09 0.0005 3.203e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.397e-09 0 3.4e-09 0.0005 3.403e-09 0 3.497e-09 0 3.5e-09 0.0005 3.503e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.697e-09 0 3.7e-09 0.0005 3.703e-09 0 3.797e-09 0 3.8e-09 0.0005 3.803e-09 0)
L_DFF_IG1_01|1 IG1_0_W _DFF_IG1_01|1  2.067833848e-12
L_DFF_IG1_01|2 _DFF_IG1_01|1 _DFF_IG1_01|2  4.135667696e-12
L_DFF_IG1_01|3 _DFF_IG1_01|3 _DFF_IG1_01|4  8.271335392e-12
L_DFF_IG1_01|4 _DFF_IG1_01|5 _DFF_IG1_01|T1  4.135667696e-12
L_DFF_IG1_01|T CLK9 _DFF_IG1_01|T1  2.067833848e-12
L_DFF_IG1_01|5 _DFF_IG1_01|4 _DFF_IG1_01|6  4.135667696e-12
L_DFF_IG1_01|6 _DFF_IG1_01|6 IG1_1  2.067833848e-12
IT10|T 0 CLK10  PWL(0 0 -1.3e-11 0 -1e-11 0.0005 -7e-12 0 8.7e-11 0 9e-11 0.0005 9.3e-11 0 1.87e-10 0 1.9e-10 0.0005 1.93e-10 0 2.87e-10 0 2.9e-10 0.0005 2.93e-10 0 3.87e-10 0 3.9e-10 0.0005 3.93e-10 0 4.87e-10 0 4.9e-10 0.0005 4.93e-10 0 5.87e-10 0 5.9e-10 0.0005 5.93e-10 0 6.87e-10 0 6.9e-10 0.0005 6.93e-10 0 7.87e-10 0 7.9e-10 0.0005 7.93e-10 0 8.87e-10 0 8.9e-10 0.0005 8.93e-10 0 9.87e-10 0 9.9e-10 0.0005 9.93e-10 0 1.087e-09 0 1.09e-09 0.0005 1.093e-09 0 1.187e-09 0 1.19e-09 0.0005 1.193e-09 0 1.287e-09 0 1.29e-09 0.0005 1.293e-09 0 1.387e-09 0 1.39e-09 0.0005 1.393e-09 0 1.487e-09 0 1.49e-09 0.0005 1.493e-09 0 1.587e-09 0 1.59e-09 0.0005 1.593e-09 0 1.687e-09 0 1.69e-09 0.0005 1.693e-09 0 1.787e-09 0 1.79e-09 0.0005 1.793e-09 0 1.887e-09 0 1.89e-09 0.0005 1.893e-09 0 1.987e-09 0 1.99e-09 0.0005 1.993e-09 0 2.087e-09 0 2.09e-09 0.0005 2.093e-09 0 2.187e-09 0 2.19e-09 0.0005 2.193e-09 0 2.287e-09 0 2.29e-09 0.0005 2.293e-09 0 2.387e-09 0 2.39e-09 0.0005 2.393e-09 0 2.487e-09 0 2.49e-09 0.0005 2.493e-09 0 2.587e-09 0 2.59e-09 0.0005 2.593e-09 0 2.687e-09 0 2.69e-09 0.0005 2.693e-09 0 2.787e-09 0 2.79e-09 0.0005 2.793e-09 0 2.887e-09 0 2.89e-09 0.0005 2.893e-09 0 2.987e-09 0 2.99e-09 0.0005 2.993e-09 0 3.087e-09 0 3.09e-09 0.0005 3.093e-09 0 3.187e-09 0 3.19e-09 0.0005 3.193e-09 0 3.287e-09 0 3.29e-09 0.0005 3.293e-09 0 3.387e-09 0 3.39e-09 0.0005 3.393e-09 0 3.487e-09 0 3.49e-09 0.0005 3.493e-09 0 3.587e-09 0 3.59e-09 0.0005 3.593e-09 0 3.687e-09 0 3.69e-09 0.0005 3.693e-09 0 3.787e-09 0 3.79e-09 0.0005 3.793e-09 0)
L_DFF_S2|1 G1_1 _DFF_S2|1  2.067833848e-12
L_DFF_S2|2 _DFF_S2|1 _DFF_S2|2  4.135667696e-12
L_DFF_S2|3 _DFF_S2|3 _DFF_S2|4  8.271335392e-12
L_DFF_S2|4 _DFF_S2|5 _DFF_S2|T1  4.135667696e-12
L_DFF_S2|T CLK10 _DFF_S2|T1  2.067833848e-12
L_DFF_S2|5 _DFF_S2|4 _DFF_S2|6  4.135667696e-12
L_DFF_S2|6 _DFF_S2|6 S2  2.067833848e-12
L_INITIAL_0|_SPL_A|1 A0 _INITIAL_0|_SPL_A|D1  2e-12
L_INITIAL_0|_SPL_A|2 _INITIAL_0|_SPL_A|D1 _INITIAL_0|_SPL_A|D2  4.135667696e-12
L_INITIAL_0|_SPL_A|3 _INITIAL_0|_SPL_A|D2 _INITIAL_0|_SPL_A|JCT  1.4770241771428573e-12
L_INITIAL_0|_SPL_A|4 _INITIAL_0|_SPL_A|JCT _INITIAL_0|_SPL_A|QA1  1.4770241771428573e-12
L_INITIAL_0|_SPL_A|5 _INITIAL_0|_SPL_A|QA1 _INITIAL_0|A1  2e-12
L_INITIAL_0|_SPL_A|6 _INITIAL_0|_SPL_A|JCT _INITIAL_0|_SPL_A|QB1  1.4770241771428573e-12
L_INITIAL_0|_SPL_A|7 _INITIAL_0|_SPL_A|QB1 _INITIAL_0|A2  2e-12
L_INITIAL_0|_SPL_B|1 B0 _INITIAL_0|_SPL_B|D1  2e-12
L_INITIAL_0|_SPL_B|2 _INITIAL_0|_SPL_B|D1 _INITIAL_0|_SPL_B|D2  4.135667696e-12
L_INITIAL_0|_SPL_B|3 _INITIAL_0|_SPL_B|D2 _INITIAL_0|_SPL_B|JCT  1.4770241771428573e-12
L_INITIAL_0|_SPL_B|4 _INITIAL_0|_SPL_B|JCT _INITIAL_0|_SPL_B|QA1  1.4770241771428573e-12
L_INITIAL_0|_SPL_B|5 _INITIAL_0|_SPL_B|QA1 _INITIAL_0|B1  2e-12
L_INITIAL_0|_SPL_B|6 _INITIAL_0|_SPL_B|JCT _INITIAL_0|_SPL_B|QB1  1.4770241771428573e-12
L_INITIAL_0|_SPL_B|7 _INITIAL_0|_SPL_B|QB1 _INITIAL_0|B2  2e-12
L_INITIAL_0|_DFF_A|1 _INITIAL_0|A1 _INITIAL_0|_DFF_A|1  2.067833848e-12
L_INITIAL_0|_DFF_A|2 _INITIAL_0|_DFF_A|1 _INITIAL_0|_DFF_A|2  4.135667696e-12
L_INITIAL_0|_DFF_A|3 _INITIAL_0|_DFF_A|3 _INITIAL_0|_DFF_A|4  8.271335392e-12
L_INITIAL_0|_DFF_A|4 _INITIAL_0|_DFF_A|5 _INITIAL_0|_DFF_A|T1  4.135667696e-12
L_INITIAL_0|_DFF_A|T CLK1 _INITIAL_0|_DFF_A|T1  2.067833848e-12
L_INITIAL_0|_DFF_A|5 _INITIAL_0|_DFF_A|4 _INITIAL_0|_DFF_A|6  4.135667696e-12
L_INITIAL_0|_DFF_A|6 _INITIAL_0|_DFF_A|6 _INITIAL_0|A1_SYNC  2.067833848e-12
L_INITIAL_0|_DFF_B|1 _INITIAL_0|B1 _INITIAL_0|_DFF_B|1  2.067833848e-12
L_INITIAL_0|_DFF_B|2 _INITIAL_0|_DFF_B|1 _INITIAL_0|_DFF_B|2  4.135667696e-12
L_INITIAL_0|_DFF_B|3 _INITIAL_0|_DFF_B|3 _INITIAL_0|_DFF_B|4  8.271335392e-12
L_INITIAL_0|_DFF_B|4 _INITIAL_0|_DFF_B|5 _INITIAL_0|_DFF_B|T1  4.135667696e-12
L_INITIAL_0|_DFF_B|T CLK1 _INITIAL_0|_DFF_B|T1  2.067833848e-12
L_INITIAL_0|_DFF_B|5 _INITIAL_0|_DFF_B|4 _INITIAL_0|_DFF_B|6  4.135667696e-12
L_INITIAL_0|_DFF_B|6 _INITIAL_0|_DFF_B|6 _INITIAL_0|B1_SYNC  2.067833848e-12
L_INITIAL_0|_XOR|A1 _INITIAL_0|A2 _INITIAL_0|_XOR|A1  2.067833848e-12
L_INITIAL_0|_XOR|A2 _INITIAL_0|_XOR|A1 _INITIAL_0|_XOR|A2  4.135667696e-12
L_INITIAL_0|_XOR|A3 _INITIAL_0|_XOR|A3 _INITIAL_0|_XOR|AB  8.271335392e-12
L_INITIAL_0|_XOR|B1 _INITIAL_0|B2 _INITIAL_0|_XOR|B1  2.067833848e-12
L_INITIAL_0|_XOR|B2 _INITIAL_0|_XOR|B1 _INITIAL_0|_XOR|B2  4.135667696e-12
L_INITIAL_0|_XOR|B3 _INITIAL_0|_XOR|B3 _INITIAL_0|_XOR|AB  8.271335392e-12
L_INITIAL_0|_XOR|T1 CLK1 _INITIAL_0|_XOR|T1  2.067833848e-12
L_INITIAL_0|_XOR|T2 _INITIAL_0|_XOR|T1 _INITIAL_0|_XOR|T2  4.135667696e-12
L_INITIAL_0|_XOR|Q2 _INITIAL_0|_XOR|ABTQ _INITIAL_0|_XOR|Q1  4.135667696e-12
L_INITIAL_0|_XOR|Q1 _INITIAL_0|_XOR|Q1 IP0_0  2.067833848e-12
L_INITIAL_0|_AND|A1 _INITIAL_0|A1_SYNC _INITIAL_0|_AND|A1  2.067833848e-12
L_INITIAL_0|_AND|A2 _INITIAL_0|_AND|A1 _INITIAL_0|_AND|A2  4.135667696e-12
L_INITIAL_0|_AND|A3 _INITIAL_0|_AND|A3 _INITIAL_0|_AND|Q3  1.2e-12
L_INITIAL_0|_AND|B1 _INITIAL_0|B1_SYNC _INITIAL_0|_AND|B1  2.067833848e-12
L_INITIAL_0|_AND|B2 _INITIAL_0|_AND|B1 _INITIAL_0|_AND|B2  4.135667696e-12
L_INITIAL_0|_AND|B3 _INITIAL_0|_AND|B3 _INITIAL_0|_AND|Q3  1.2e-12
L_INITIAL_0|_AND|Q3 _INITIAL_0|_AND|Q3 _INITIAL_0|_AND|Q2  4.135667696e-12
L_INITIAL_0|_AND|Q2 _INITIAL_0|_AND|Q2 _INITIAL_0|_AND|Q1  4.135667696e-12
L_INITIAL_0|_AND|Q1 _INITIAL_0|_AND|Q1 IG0_0  2.067833848e-12
L_INITIAL_1|_SPL_A|1 A1 _INITIAL_1|_SPL_A|D1  2e-12
L_INITIAL_1|_SPL_A|2 _INITIAL_1|_SPL_A|D1 _INITIAL_1|_SPL_A|D2  4.135667696e-12
L_INITIAL_1|_SPL_A|3 _INITIAL_1|_SPL_A|D2 _INITIAL_1|_SPL_A|JCT  1.4770241771428573e-12
L_INITIAL_1|_SPL_A|4 _INITIAL_1|_SPL_A|JCT _INITIAL_1|_SPL_A|QA1  1.4770241771428573e-12
L_INITIAL_1|_SPL_A|5 _INITIAL_1|_SPL_A|QA1 _INITIAL_1|A1  2e-12
L_INITIAL_1|_SPL_A|6 _INITIAL_1|_SPL_A|JCT _INITIAL_1|_SPL_A|QB1  1.4770241771428573e-12
L_INITIAL_1|_SPL_A|7 _INITIAL_1|_SPL_A|QB1 _INITIAL_1|A2  2e-12
L_INITIAL_1|_SPL_B|1 B1 _INITIAL_1|_SPL_B|D1  2e-12
L_INITIAL_1|_SPL_B|2 _INITIAL_1|_SPL_B|D1 _INITIAL_1|_SPL_B|D2  4.135667696e-12
L_INITIAL_1|_SPL_B|3 _INITIAL_1|_SPL_B|D2 _INITIAL_1|_SPL_B|JCT  1.4770241771428573e-12
L_INITIAL_1|_SPL_B|4 _INITIAL_1|_SPL_B|JCT _INITIAL_1|_SPL_B|QA1  1.4770241771428573e-12
L_INITIAL_1|_SPL_B|5 _INITIAL_1|_SPL_B|QA1 _INITIAL_1|B1  2e-12
L_INITIAL_1|_SPL_B|6 _INITIAL_1|_SPL_B|JCT _INITIAL_1|_SPL_B|QB1  1.4770241771428573e-12
L_INITIAL_1|_SPL_B|7 _INITIAL_1|_SPL_B|QB1 _INITIAL_1|B2  2e-12
L_INITIAL_1|_DFF_A|1 _INITIAL_1|A1 _INITIAL_1|_DFF_A|1  2.067833848e-12
L_INITIAL_1|_DFF_A|2 _INITIAL_1|_DFF_A|1 _INITIAL_1|_DFF_A|2  4.135667696e-12
L_INITIAL_1|_DFF_A|3 _INITIAL_1|_DFF_A|3 _INITIAL_1|_DFF_A|4  8.271335392e-12
L_INITIAL_1|_DFF_A|4 _INITIAL_1|_DFF_A|5 _INITIAL_1|_DFF_A|T1  4.135667696e-12
L_INITIAL_1|_DFF_A|T CLK2 _INITIAL_1|_DFF_A|T1  2.067833848e-12
L_INITIAL_1|_DFF_A|5 _INITIAL_1|_DFF_A|4 _INITIAL_1|_DFF_A|6  4.135667696e-12
L_INITIAL_1|_DFF_A|6 _INITIAL_1|_DFF_A|6 _INITIAL_1|A1_SYNC  2.067833848e-12
L_INITIAL_1|_DFF_B|1 _INITIAL_1|B1 _INITIAL_1|_DFF_B|1  2.067833848e-12
L_INITIAL_1|_DFF_B|2 _INITIAL_1|_DFF_B|1 _INITIAL_1|_DFF_B|2  4.135667696e-12
L_INITIAL_1|_DFF_B|3 _INITIAL_1|_DFF_B|3 _INITIAL_1|_DFF_B|4  8.271335392e-12
L_INITIAL_1|_DFF_B|4 _INITIAL_1|_DFF_B|5 _INITIAL_1|_DFF_B|T1  4.135667696e-12
L_INITIAL_1|_DFF_B|T CLK2 _INITIAL_1|_DFF_B|T1  2.067833848e-12
L_INITIAL_1|_DFF_B|5 _INITIAL_1|_DFF_B|4 _INITIAL_1|_DFF_B|6  4.135667696e-12
L_INITIAL_1|_DFF_B|6 _INITIAL_1|_DFF_B|6 _INITIAL_1|B1_SYNC  2.067833848e-12
L_INITIAL_1|_XOR|A1 _INITIAL_1|A2 _INITIAL_1|_XOR|A1  2.067833848e-12
L_INITIAL_1|_XOR|A2 _INITIAL_1|_XOR|A1 _INITIAL_1|_XOR|A2  4.135667696e-12
L_INITIAL_1|_XOR|A3 _INITIAL_1|_XOR|A3 _INITIAL_1|_XOR|AB  8.271335392e-12
L_INITIAL_1|_XOR|B1 _INITIAL_1|B2 _INITIAL_1|_XOR|B1  2.067833848e-12
L_INITIAL_1|_XOR|B2 _INITIAL_1|_XOR|B1 _INITIAL_1|_XOR|B2  4.135667696e-12
L_INITIAL_1|_XOR|B3 _INITIAL_1|_XOR|B3 _INITIAL_1|_XOR|AB  8.271335392e-12
L_INITIAL_1|_XOR|T1 CLK2 _INITIAL_1|_XOR|T1  2.067833848e-12
L_INITIAL_1|_XOR|T2 _INITIAL_1|_XOR|T1 _INITIAL_1|_XOR|T2  4.135667696e-12
L_INITIAL_1|_XOR|Q2 _INITIAL_1|_XOR|ABTQ _INITIAL_1|_XOR|Q1  4.135667696e-12
L_INITIAL_1|_XOR|Q1 _INITIAL_1|_XOR|Q1 IP1_0  2.067833848e-12
L_INITIAL_1|_AND|A1 _INITIAL_1|A1_SYNC _INITIAL_1|_AND|A1  2.067833848e-12
L_INITIAL_1|_AND|A2 _INITIAL_1|_AND|A1 _INITIAL_1|_AND|A2  4.135667696e-12
L_INITIAL_1|_AND|A3 _INITIAL_1|_AND|A3 _INITIAL_1|_AND|Q3  1.2e-12
L_INITIAL_1|_AND|B1 _INITIAL_1|B1_SYNC _INITIAL_1|_AND|B1  2.067833848e-12
L_INITIAL_1|_AND|B2 _INITIAL_1|_AND|B1 _INITIAL_1|_AND|B2  4.135667696e-12
L_INITIAL_1|_AND|B3 _INITIAL_1|_AND|B3 _INITIAL_1|_AND|Q3  1.2e-12
L_INITIAL_1|_AND|Q3 _INITIAL_1|_AND|Q3 _INITIAL_1|_AND|Q2  4.135667696e-12
L_INITIAL_1|_AND|Q2 _INITIAL_1|_AND|Q2 _INITIAL_1|_AND|Q1  4.135667696e-12
L_INITIAL_1|_AND|Q1 _INITIAL_1|_AND|Q1 IG1_0  2.067833848e-12
L_SPL_P0|I_D1|B _SPL_P0|D1 _SPL_P0|I_D1|MID  2e-12
I_SPL_P0|I_D1|B 0 _SPL_P0|I_D1|MID  0.000175
L_SPL_P0|I_D2|B _SPL_P0|D2 _SPL_P0|I_D2|MID  2e-12
I_SPL_P0|I_D2|B 0 _SPL_P0|I_D2|MID  0.000245
L_SPL_P0|I_Q1|B _SPL_P0|QA1 _SPL_P0|I_Q1|MID  2e-12
I_SPL_P0|I_Q1|B 0 _SPL_P0|I_Q1|MID  0.000175
L_SPL_P0|I_Q2|B _SPL_P0|QB1 _SPL_P0|I_Q2|MID  2e-12
I_SPL_P0|I_Q2|B 0 _SPL_P0|I_Q2|MID  0.000175
B_SPL_P0|1|1 _SPL_P0|D1 _SPL_P0|1|MID_SERIES JJMIT AREA=2.5
L_SPL_P0|1|P _SPL_P0|1|MID_SERIES 0  2e-13
R_SPL_P0|1|B _SPL_P0|D1 _SPL_P0|1|MID_SHUNT  2.7439617672
L_SPL_P0|1|RB _SPL_P0|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_P0|2|1 _SPL_P0|D2 _SPL_P0|2|MID_SERIES JJMIT AREA=2.5
L_SPL_P0|2|P _SPL_P0|2|MID_SERIES 0  2e-13
R_SPL_P0|2|B _SPL_P0|D2 _SPL_P0|2|MID_SHUNT  2.7439617672
L_SPL_P0|2|RB _SPL_P0|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_P0|A|1 _SPL_P0|QA1 _SPL_P0|A|MID_SERIES JJMIT AREA=2.5
L_SPL_P0|A|P _SPL_P0|A|MID_SERIES 0  2e-13
R_SPL_P0|A|B _SPL_P0|QA1 _SPL_P0|A|MID_SHUNT  2.7439617672
L_SPL_P0|A|RB _SPL_P0|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_P0|B|1 _SPL_P0|QB1 _SPL_P0|B|MID_SERIES JJMIT AREA=2.5
L_SPL_P0|B|P _SPL_P0|B|MID_SERIES 0  2e-13
R_SPL_P0|B|B _SPL_P0|QB1 _SPL_P0|B|MID_SHUNT  2.7439617672
L_SPL_P0|B|RB _SPL_P0|B|MID_SHUNT 0  1.550338398468e-12
L_SPL_G0|I_D1|B _SPL_G0|D1 _SPL_G0|I_D1|MID  2e-12
I_SPL_G0|I_D1|B 0 _SPL_G0|I_D1|MID  0.000175
L_SPL_G0|I_D2|B _SPL_G0|D2 _SPL_G0|I_D2|MID  2e-12
I_SPL_G0|I_D2|B 0 _SPL_G0|I_D2|MID  0.000245
L_SPL_G0|I_Q1|B _SPL_G0|QA1 _SPL_G0|I_Q1|MID  2e-12
I_SPL_G0|I_Q1|B 0 _SPL_G0|I_Q1|MID  0.000175
L_SPL_G0|I_Q2|B _SPL_G0|QB1 _SPL_G0|I_Q2|MID  2e-12
I_SPL_G0|I_Q2|B 0 _SPL_G0|I_Q2|MID  0.000175
B_SPL_G0|1|1 _SPL_G0|D1 _SPL_G0|1|MID_SERIES JJMIT AREA=2.5
L_SPL_G0|1|P _SPL_G0|1|MID_SERIES 0  2e-13
R_SPL_G0|1|B _SPL_G0|D1 _SPL_G0|1|MID_SHUNT  2.7439617672
L_SPL_G0|1|RB _SPL_G0|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_G0|2|1 _SPL_G0|D2 _SPL_G0|2|MID_SERIES JJMIT AREA=2.5
L_SPL_G0|2|P _SPL_G0|2|MID_SERIES 0  2e-13
R_SPL_G0|2|B _SPL_G0|D2 _SPL_G0|2|MID_SHUNT  2.7439617672
L_SPL_G0|2|RB _SPL_G0|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_G0|A|1 _SPL_G0|QA1 _SPL_G0|A|MID_SERIES JJMIT AREA=2.5
L_SPL_G0|A|P _SPL_G0|A|MID_SERIES 0  2e-13
R_SPL_G0|A|B _SPL_G0|QA1 _SPL_G0|A|MID_SHUNT  2.7439617672
L_SPL_G0|A|RB _SPL_G0|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_G0|B|1 _SPL_G0|QB1 _SPL_G0|B|MID_SERIES JJMIT AREA=2.5
L_SPL_G0|B|P _SPL_G0|B|MID_SERIES 0  2e-13
R_SPL_G0|B|B _SPL_G0|QB1 _SPL_G0|B|MID_SHUNT  2.7439617672
L_SPL_G0|B|RB _SPL_G0|B|MID_SHUNT 0  1.550338398468e-12
L_SPL_P1|I_D1|B _SPL_P1|D1 _SPL_P1|I_D1|MID  2e-12
I_SPL_P1|I_D1|B 0 _SPL_P1|I_D1|MID  0.000175
L_SPL_P1|I_D2|B _SPL_P1|D2 _SPL_P1|I_D2|MID  2e-12
I_SPL_P1|I_D2|B 0 _SPL_P1|I_D2|MID  0.000245
L_SPL_P1|I_Q1|B _SPL_P1|QA1 _SPL_P1|I_Q1|MID  2e-12
I_SPL_P1|I_Q1|B 0 _SPL_P1|I_Q1|MID  0.000175
L_SPL_P1|I_Q2|B _SPL_P1|QB1 _SPL_P1|I_Q2|MID  2e-12
I_SPL_P1|I_Q2|B 0 _SPL_P1|I_Q2|MID  0.000175
B_SPL_P1|1|1 _SPL_P1|D1 _SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_SPL_P1|1|P _SPL_P1|1|MID_SERIES 0  2e-13
R_SPL_P1|1|B _SPL_P1|D1 _SPL_P1|1|MID_SHUNT  2.7439617672
L_SPL_P1|1|RB _SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_P1|2|1 _SPL_P1|D2 _SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_SPL_P1|2|P _SPL_P1|2|MID_SERIES 0  2e-13
R_SPL_P1|2|B _SPL_P1|D2 _SPL_P1|2|MID_SHUNT  2.7439617672
L_SPL_P1|2|RB _SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_P1|A|1 _SPL_P1|QA1 _SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_SPL_P1|A|P _SPL_P1|A|MID_SERIES 0  2e-13
R_SPL_P1|A|B _SPL_P1|QA1 _SPL_P1|A|MID_SHUNT  2.7439617672
L_SPL_P1|A|RB _SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_P1|B|1 _SPL_P1|QB1 _SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_SPL_P1|B|P _SPL_P1|B|MID_SERIES 0  2e-13
R_SPL_P1|B|B _SPL_P1|QB1 _SPL_P1|B|MID_SHUNT  2.7439617672
L_SPL_P1|B|RB _SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_SPL_G1|I_D1|B _SPL_G1|D1 _SPL_G1|I_D1|MID  2e-12
I_SPL_G1|I_D1|B 0 _SPL_G1|I_D1|MID  0.000175
L_SPL_G1|I_D2|B _SPL_G1|D2 _SPL_G1|I_D2|MID  2e-12
I_SPL_G1|I_D2|B 0 _SPL_G1|I_D2|MID  0.000245
L_SPL_G1|I_Q1|B _SPL_G1|QA1 _SPL_G1|I_Q1|MID  2e-12
I_SPL_G1|I_Q1|B 0 _SPL_G1|I_Q1|MID  0.000175
L_SPL_G1|I_Q2|B _SPL_G1|QB1 _SPL_G1|I_Q2|MID  2e-12
I_SPL_G1|I_Q2|B 0 _SPL_G1|I_Q2|MID  0.000175
B_SPL_G1|1|1 _SPL_G1|D1 _SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_SPL_G1|1|P _SPL_G1|1|MID_SERIES 0  2e-13
R_SPL_G1|1|B _SPL_G1|D1 _SPL_G1|1|MID_SHUNT  2.7439617672
L_SPL_G1|1|RB _SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_SPL_G1|2|1 _SPL_G1|D2 _SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_SPL_G1|2|P _SPL_G1|2|MID_SERIES 0  2e-13
R_SPL_G1|2|B _SPL_G1|D2 _SPL_G1|2|MID_SHUNT  2.7439617672
L_SPL_G1|2|RB _SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_SPL_G1|A|1 _SPL_G1|QA1 _SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_SPL_G1|A|P _SPL_G1|A|MID_SERIES 0  2e-13
R_SPL_G1|A|B _SPL_G1|QA1 _SPL_G1|A|MID_SHUNT  2.7439617672
L_SPL_G1|A|RB _SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_SPL_G1|B|1 _SPL_G1|QB1 _SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_SPL_G1|B|P _SPL_G1|B|MID_SERIES 0  2e-13
R_SPL_G1|B|B _SPL_G1|QB1 _SPL_G1|B|MID_SHUNT  2.7439617672
L_SPL_G1|B|RB _SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_SPL_G1|1 IG1_0_B _PG_01|_SPL_G1|D1  2e-12
L_PG_01|_SPL_G1|2 _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|D2  4.135667696e-12
L_PG_01|_SPL_G1|3 _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|JCT  1.4770241771428573e-12
L_PG_01|_SPL_G1|4 _PG_01|_SPL_G1|JCT _PG_01|_SPL_G1|QA1  1.4770241771428573e-12
L_PG_01|_SPL_G1|5 _PG_01|_SPL_G1|QA1 _PG_01|G1_COPY_1  2e-12
L_PG_01|_SPL_G1|6 _PG_01|_SPL_G1|JCT _PG_01|_SPL_G1|QB1  1.4770241771428573e-12
L_PG_01|_SPL_G1|7 _PG_01|_SPL_G1|QB1 _PG_01|G1_COPY_2  2e-12
L_PG_01|_SPL_P1|1 IP1_0_B _PG_01|_SPL_P1|D1  2e-12
L_PG_01|_SPL_P1|2 _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|D2  4.135667696e-12
L_PG_01|_SPL_P1|3 _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|JCT  1.4770241771428573e-12
L_PG_01|_SPL_P1|4 _PG_01|_SPL_P1|JCT _PG_01|_SPL_P1|QA1  1.4770241771428573e-12
L_PG_01|_SPL_P1|5 _PG_01|_SPL_P1|QA1 _PG_01|P1_COPY_1  2e-12
L_PG_01|_SPL_P1|6 _PG_01|_SPL_P1|JCT _PG_01|_SPL_P1|QB1  1.4770241771428573e-12
L_PG_01|_SPL_P1|7 _PG_01|_SPL_P1|QB1 _PG_01|P1_COPY_2  2e-12
L_PG_01|_PG|A1 _PG_01|P1_COPY_1 _PG_01|_PG|A1  2.067833848e-12
L_PG_01|_PG|A2 _PG_01|_PG|A1 _PG_01|_PG|A2  4.135667696e-12
L_PG_01|_PG|A3 _PG_01|_PG|A3 _PG_01|_PG|Q3  1.2e-12
L_PG_01|_PG|B1 _PG_01|G1_COPY_1 _PG_01|_PG|B1  2.067833848e-12
L_PG_01|_PG|B2 _PG_01|_PG|B1 _PG_01|_PG|B2  4.135667696e-12
L_PG_01|_PG|B3 _PG_01|_PG|B3 _PG_01|_PG|Q3  1.2e-12
L_PG_01|_PG|Q3 _PG_01|_PG|Q3 _PG_01|_PG|Q2  4.135667696e-12
L_PG_01|_PG|Q2 _PG_01|_PG|Q2 _PG_01|_PG|Q1  4.135667696e-12
L_PG_01|_PG|Q1 _PG_01|_PG|Q1 _PG_01|PG  2.067833848e-12
L_PG_01|_GG|A1 IG0_0_B _PG_01|_GG|A1  2.067833848e-12
L_PG_01|_GG|A2 _PG_01|_GG|A1 _PG_01|_GG|A2  4.135667696e-12
L_PG_01|_GG|A3 _PG_01|_GG|A3 _PG_01|_GG|Q3  1.2e-12
L_PG_01|_GG|B1 _PG_01|G1_COPY_2 _PG_01|_GG|B1  2.067833848e-12
L_PG_01|_GG|B2 _PG_01|_GG|B1 _PG_01|_GG|B2  4.135667696e-12
L_PG_01|_GG|B3 _PG_01|_GG|B3 _PG_01|_GG|Q3  1.2e-12
L_PG_01|_GG|Q3 _PG_01|_GG|Q3 _PG_01|_GG|Q2  4.135667696e-12
L_PG_01|_GG|Q2 _PG_01|_GG|Q2 _PG_01|_GG|Q1  4.135667696e-12
L_PG_01|_GG|Q1 _PG_01|_GG|Q1 _PG_01|GG  2.067833848e-12
L_PG_01|_DFF_P0|1 IP0_0_B _PG_01|_DFF_P0|1  2.067833848e-12
L_PG_01|_DFF_P0|2 _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|2  4.135667696e-12
L_PG_01|_DFF_P0|3 _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|4  8.271335392e-12
L_PG_01|_DFF_P0|4 _PG_01|_DFF_P0|5 _PG_01|_DFF_P0|T1  4.135667696e-12
L_PG_01|_DFF_P0|T CLK3 _PG_01|_DFF_P0|T1  2.067833848e-12
L_PG_01|_DFF_P0|5 _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|6  4.135667696e-12
L_PG_01|_DFF_P0|6 _PG_01|_DFF_P0|6 _PG_01|P0_SYNC  2.067833848e-12
L_PG_01|_DFF_P1|1 _PG_01|P1_COPY_2 _PG_01|_DFF_P1|1  2.067833848e-12
L_PG_01|_DFF_P1|2 _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|2  4.135667696e-12
L_PG_01|_DFF_P1|3 _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|4  8.271335392e-12
L_PG_01|_DFF_P1|4 _PG_01|_DFF_P1|5 _PG_01|_DFF_P1|T1  4.135667696e-12
L_PG_01|_DFF_P1|T CLK3 _PG_01|_DFF_P1|T1  2.067833848e-12
L_PG_01|_DFF_P1|5 _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|6  4.135667696e-12
L_PG_01|_DFF_P1|6 _PG_01|_DFF_P1|6 _PG_01|P1_SYNC  2.067833848e-12
L_PG_01|_DFF_PG|1 _PG_01|PG _PG_01|_DFF_PG|1  2.067833848e-12
L_PG_01|_DFF_PG|2 _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|2  4.135667696e-12
L_PG_01|_DFF_PG|3 _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|4  8.271335392e-12
L_PG_01|_DFF_PG|4 _PG_01|_DFF_PG|5 _PG_01|_DFF_PG|T1  4.135667696e-12
L_PG_01|_DFF_PG|T CLK3 _PG_01|_DFF_PG|T1  2.067833848e-12
L_PG_01|_DFF_PG|5 _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|6  4.135667696e-12
L_PG_01|_DFF_PG|6 _PG_01|_DFF_PG|6 _PG_01|PG_SYNC  2.067833848e-12
L_PG_01|_DFF_GG|1 _PG_01|GG _PG_01|_DFF_GG|1  2.067833848e-12
L_PG_01|_DFF_GG|2 _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|2  4.135667696e-12
L_PG_01|_DFF_GG|3 _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|4  8.271335392e-12
L_PG_01|_DFF_GG|4 _PG_01|_DFF_GG|5 _PG_01|_DFF_GG|T1  4.135667696e-12
L_PG_01|_DFF_GG|T CLK3 _PG_01|_DFF_GG|T1  2.067833848e-12
L_PG_01|_DFF_GG|5 _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|6  4.135667696e-12
L_PG_01|_DFF_GG|6 _PG_01|_DFF_GG|6 _PG_01|GG_SYNC  2.067833848e-12
L_PG_01|_AND_G|A1 _PG_01|PG_SYNC _PG_01|_AND_G|A1  2.067833848e-12
L_PG_01|_AND_G|A2 _PG_01|_AND_G|A1 _PG_01|_AND_G|A2  4.135667696e-12
L_PG_01|_AND_G|A3 _PG_01|_AND_G|A3 _PG_01|_AND_G|Q3  1.2e-12
L_PG_01|_AND_G|B1 _PG_01|GG_SYNC _PG_01|_AND_G|B1  2.067833848e-12
L_PG_01|_AND_G|B2 _PG_01|_AND_G|B1 _PG_01|_AND_G|B2  4.135667696e-12
L_PG_01|_AND_G|B3 _PG_01|_AND_G|B3 _PG_01|_AND_G|Q3  1.2e-12
L_PG_01|_AND_G|Q3 _PG_01|_AND_G|Q3 _PG_01|_AND_G|Q2  4.135667696e-12
L_PG_01|_AND_G|Q2 _PG_01|_AND_G|Q2 _PG_01|_AND_G|Q1  4.135667696e-12
L_PG_01|_AND_G|Q1 _PG_01|_AND_G|Q1 G1_1  2.067833848e-12
L_PG_01|_AND_P|A1 _PG_01|P0_SYNC _PG_01|_AND_P|A1  2.067833848e-12
L_PG_01|_AND_P|A2 _PG_01|_AND_P|A1 _PG_01|_AND_P|A2  4.135667696e-12
L_PG_01|_AND_P|A3 _PG_01|_AND_P|A3 _PG_01|_AND_P|Q3  1.2e-12
L_PG_01|_AND_P|B1 _PG_01|P1_SYNC _PG_01|_AND_P|B1  2.067833848e-12
L_PG_01|_AND_P|B2 _PG_01|_AND_P|B1 _PG_01|_AND_P|B2  4.135667696e-12
L_PG_01|_AND_P|B3 _PG_01|_AND_P|B3 _PG_01|_AND_P|Q3  1.2e-12
L_PG_01|_AND_P|Q3 _PG_01|_AND_P|Q3 _PG_01|_AND_P|Q2  4.135667696e-12
L_PG_01|_AND_P|Q2 _PG_01|_AND_P|Q2 _PG_01|_AND_P|Q1  4.135667696e-12
L_PG_01|_AND_P|Q1 _PG_01|_AND_P|Q1 P1_1  2.067833848e-12
B_DFF_IP0_01|1|1 _DFF_IP0_01|1 _DFF_IP0_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_01|1|P _DFF_IP0_01|1|MID_SERIES 0  2e-13
R_DFF_IP0_01|1|B _DFF_IP0_01|1 _DFF_IP0_01|1|MID_SHUNT  2.7439617672
L_DFF_IP0_01|1|RB _DFF_IP0_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_01|23|1 _DFF_IP0_01|2 _DFF_IP0_01|3 JJMIT AREA=1.7857142857142858
R_DFF_IP0_01|23|B _DFF_IP0_01|2 _DFF_IP0_01|23|MID_SHUNT  3.84154647408
L_DFF_IP0_01|23|RB _DFF_IP0_01|23|MID_SHUNT _DFF_IP0_01|3  2.1704737578552e-12
B_DFF_IP0_01|3|1 _DFF_IP0_01|3 _DFF_IP0_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_01|3|P _DFF_IP0_01|3|MID_SERIES 0  2e-13
R_DFF_IP0_01|3|B _DFF_IP0_01|3 _DFF_IP0_01|3|MID_SHUNT  2.7439617672
L_DFF_IP0_01|3|RB _DFF_IP0_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_01|4|1 _DFF_IP0_01|4 _DFF_IP0_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_01|4|P _DFF_IP0_01|4|MID_SERIES 0  2e-13
R_DFF_IP0_01|4|B _DFF_IP0_01|4 _DFF_IP0_01|4|MID_SHUNT  2.7439617672
L_DFF_IP0_01|4|RB _DFF_IP0_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_01|45|1 _DFF_IP0_01|4 _DFF_IP0_01|5 JJMIT AREA=1.7857142857142858
R_DFF_IP0_01|45|B _DFF_IP0_01|4 _DFF_IP0_01|45|MID_SHUNT  3.84154647408
L_DFF_IP0_01|45|RB _DFF_IP0_01|45|MID_SHUNT _DFF_IP0_01|5  2.1704737578552e-12
B_DFF_IP0_01|T|1 _DFF_IP0_01|T1 _DFF_IP0_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_01|T|P _DFF_IP0_01|T|MID_SERIES 0  2e-13
R_DFF_IP0_01|T|B _DFF_IP0_01|T1 _DFF_IP0_01|T|MID_SHUNT  2.7439617672
L_DFF_IP0_01|T|RB _DFF_IP0_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_01|6|1 _DFF_IP0_01|6 _DFF_IP0_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_01|6|P _DFF_IP0_01|6|MID_SERIES 0  2e-13
R_DFF_IP0_01|6|B _DFF_IP0_01|6 _DFF_IP0_01|6|MID_SHUNT  2.7439617672
L_DFF_IP0_01|6|RB _DFF_IP0_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP0_01|I_1|B _DFF_IP0_01|1 _DFF_IP0_01|I_1|MID  2e-12
I_DFF_IP0_01|I_1|B 0 _DFF_IP0_01|I_1|MID  0.000175
L_DFF_IP0_01|I_3|B _DFF_IP0_01|3 _DFF_IP0_01|I_3|MID  2e-12
I_DFF_IP0_01|I_3|B 0 _DFF_IP0_01|I_3|MID  0.00025
L_DFF_IP0_01|I_T|B _DFF_IP0_01|T1 _DFF_IP0_01|I_T|MID  2e-12
I_DFF_IP0_01|I_T|B 0 _DFF_IP0_01|I_T|MID  0.000175
L_DFF_IP0_01|I_6|B _DFF_IP0_01|6 _DFF_IP0_01|I_6|MID  2e-12
I_DFF_IP0_01|I_6|B 0 _DFF_IP0_01|I_6|MID  0.000175
B_DFF_IP0_12|1|1 _DFF_IP0_12|1 _DFF_IP0_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_12|1|P _DFF_IP0_12|1|MID_SERIES 0  2e-13
R_DFF_IP0_12|1|B _DFF_IP0_12|1 _DFF_IP0_12|1|MID_SHUNT  2.7439617672
L_DFF_IP0_12|1|RB _DFF_IP0_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_12|23|1 _DFF_IP0_12|2 _DFF_IP0_12|3 JJMIT AREA=1.7857142857142858
R_DFF_IP0_12|23|B _DFF_IP0_12|2 _DFF_IP0_12|23|MID_SHUNT  3.84154647408
L_DFF_IP0_12|23|RB _DFF_IP0_12|23|MID_SHUNT _DFF_IP0_12|3  2.1704737578552e-12
B_DFF_IP0_12|3|1 _DFF_IP0_12|3 _DFF_IP0_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_12|3|P _DFF_IP0_12|3|MID_SERIES 0  2e-13
R_DFF_IP0_12|3|B _DFF_IP0_12|3 _DFF_IP0_12|3|MID_SHUNT  2.7439617672
L_DFF_IP0_12|3|RB _DFF_IP0_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_12|4|1 _DFF_IP0_12|4 _DFF_IP0_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_12|4|P _DFF_IP0_12|4|MID_SERIES 0  2e-13
R_DFF_IP0_12|4|B _DFF_IP0_12|4 _DFF_IP0_12|4|MID_SHUNT  2.7439617672
L_DFF_IP0_12|4|RB _DFF_IP0_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_12|45|1 _DFF_IP0_12|4 _DFF_IP0_12|5 JJMIT AREA=1.7857142857142858
R_DFF_IP0_12|45|B _DFF_IP0_12|4 _DFF_IP0_12|45|MID_SHUNT  3.84154647408
L_DFF_IP0_12|45|RB _DFF_IP0_12|45|MID_SHUNT _DFF_IP0_12|5  2.1704737578552e-12
B_DFF_IP0_12|T|1 _DFF_IP0_12|T1 _DFF_IP0_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_12|T|P _DFF_IP0_12|T|MID_SERIES 0  2e-13
R_DFF_IP0_12|T|B _DFF_IP0_12|T1 _DFF_IP0_12|T|MID_SHUNT  2.7439617672
L_DFF_IP0_12|T|RB _DFF_IP0_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP0_12|6|1 _DFF_IP0_12|6 _DFF_IP0_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP0_12|6|P _DFF_IP0_12|6|MID_SERIES 0  2e-13
R_DFF_IP0_12|6|B _DFF_IP0_12|6 _DFF_IP0_12|6|MID_SHUNT  2.7439617672
L_DFF_IP0_12|6|RB _DFF_IP0_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP0_12|I_1|B _DFF_IP0_12|1 _DFF_IP0_12|I_1|MID  2e-12
I_DFF_IP0_12|I_1|B 0 _DFF_IP0_12|I_1|MID  0.000175
L_DFF_IP0_12|I_3|B _DFF_IP0_12|3 _DFF_IP0_12|I_3|MID  2e-12
I_DFF_IP0_12|I_3|B 0 _DFF_IP0_12|I_3|MID  0.00025
L_DFF_IP0_12|I_T|B _DFF_IP0_12|T1 _DFF_IP0_12|I_T|MID  2e-12
I_DFF_IP0_12|I_T|B 0 _DFF_IP0_12|I_T|MID  0.000175
L_DFF_IP0_12|I_6|B _DFF_IP0_12|6 _DFF_IP0_12|I_6|MID  2e-12
I_DFF_IP0_12|I_6|B 0 _DFF_IP0_12|I_6|MID  0.000175
B_DFF_IG0_01|1|1 _DFF_IG0_01|1 _DFF_IG0_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IG0_01|1|P _DFF_IG0_01|1|MID_SERIES 0  2e-13
R_DFF_IG0_01|1|B _DFF_IG0_01|1 _DFF_IG0_01|1|MID_SHUNT  2.7439617672
L_DFF_IG0_01|1|RB _DFF_IG0_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG0_01|23|1 _DFF_IG0_01|2 _DFF_IG0_01|3 JJMIT AREA=1.7857142857142858
R_DFF_IG0_01|23|B _DFF_IG0_01|2 _DFF_IG0_01|23|MID_SHUNT  3.84154647408
L_DFF_IG0_01|23|RB _DFF_IG0_01|23|MID_SHUNT _DFF_IG0_01|3  2.1704737578552e-12
B_DFF_IG0_01|3|1 _DFF_IG0_01|3 _DFF_IG0_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IG0_01|3|P _DFF_IG0_01|3|MID_SERIES 0  2e-13
R_DFF_IG0_01|3|B _DFF_IG0_01|3 _DFF_IG0_01|3|MID_SHUNT  2.7439617672
L_DFF_IG0_01|3|RB _DFF_IG0_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG0_01|4|1 _DFF_IG0_01|4 _DFF_IG0_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IG0_01|4|P _DFF_IG0_01|4|MID_SERIES 0  2e-13
R_DFF_IG0_01|4|B _DFF_IG0_01|4 _DFF_IG0_01|4|MID_SHUNT  2.7439617672
L_DFF_IG0_01|4|RB _DFF_IG0_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG0_01|45|1 _DFF_IG0_01|4 _DFF_IG0_01|5 JJMIT AREA=1.7857142857142858
R_DFF_IG0_01|45|B _DFF_IG0_01|4 _DFF_IG0_01|45|MID_SHUNT  3.84154647408
L_DFF_IG0_01|45|RB _DFF_IG0_01|45|MID_SHUNT _DFF_IG0_01|5  2.1704737578552e-12
B_DFF_IG0_01|T|1 _DFF_IG0_01|T1 _DFF_IG0_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IG0_01|T|P _DFF_IG0_01|T|MID_SERIES 0  2e-13
R_DFF_IG0_01|T|B _DFF_IG0_01|T1 _DFF_IG0_01|T|MID_SHUNT  2.7439617672
L_DFF_IG0_01|T|RB _DFF_IG0_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG0_01|6|1 _DFF_IG0_01|6 _DFF_IG0_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IG0_01|6|P _DFF_IG0_01|6|MID_SERIES 0  2e-13
R_DFF_IG0_01|6|B _DFF_IG0_01|6 _DFF_IG0_01|6|MID_SHUNT  2.7439617672
L_DFF_IG0_01|6|RB _DFF_IG0_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IG0_01|I_1|B _DFF_IG0_01|1 _DFF_IG0_01|I_1|MID  2e-12
I_DFF_IG0_01|I_1|B 0 _DFF_IG0_01|I_1|MID  0.000175
L_DFF_IG0_01|I_3|B _DFF_IG0_01|3 _DFF_IG0_01|I_3|MID  2e-12
I_DFF_IG0_01|I_3|B 0 _DFF_IG0_01|I_3|MID  0.00025
L_DFF_IG0_01|I_T|B _DFF_IG0_01|T1 _DFF_IG0_01|I_T|MID  2e-12
I_DFF_IG0_01|I_T|B 0 _DFF_IG0_01|I_T|MID  0.000175
L_DFF_IG0_01|I_6|B _DFF_IG0_01|6 _DFF_IG0_01|I_6|MID  2e-12
I_DFF_IG0_01|I_6|B 0 _DFF_IG0_01|I_6|MID  0.000175
B_DFF_IP1_01|1|1 _DFF_IP1_01|1 _DFF_IP1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|1|P _DFF_IP1_01|1|MID_SERIES 0  2e-13
R_DFF_IP1_01|1|B _DFF_IP1_01|1 _DFF_IP1_01|1|MID_SHUNT  2.7439617672
L_DFF_IP1_01|1|RB _DFF_IP1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|23|1 _DFF_IP1_01|2 _DFF_IP1_01|3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|23|B _DFF_IP1_01|2 _DFF_IP1_01|23|MID_SHUNT  3.84154647408
L_DFF_IP1_01|23|RB _DFF_IP1_01|23|MID_SHUNT _DFF_IP1_01|3  2.1704737578552e-12
B_DFF_IP1_01|3|1 _DFF_IP1_01|3 _DFF_IP1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|3|P _DFF_IP1_01|3|MID_SERIES 0  2e-13
R_DFF_IP1_01|3|B _DFF_IP1_01|3 _DFF_IP1_01|3|MID_SHUNT  2.7439617672
L_DFF_IP1_01|3|RB _DFF_IP1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|4|1 _DFF_IP1_01|4 _DFF_IP1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|4|P _DFF_IP1_01|4|MID_SERIES 0  2e-13
R_DFF_IP1_01|4|B _DFF_IP1_01|4 _DFF_IP1_01|4|MID_SHUNT  2.7439617672
L_DFF_IP1_01|4|RB _DFF_IP1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|45|1 _DFF_IP1_01|4 _DFF_IP1_01|5 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|45|B _DFF_IP1_01|4 _DFF_IP1_01|45|MID_SHUNT  3.84154647408
L_DFF_IP1_01|45|RB _DFF_IP1_01|45|MID_SHUNT _DFF_IP1_01|5  2.1704737578552e-12
B_DFF_IP1_01|T|1 _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|T|P _DFF_IP1_01|T|MID_SERIES 0  2e-13
R_DFF_IP1_01|T|B _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SHUNT  2.7439617672
L_DFF_IP1_01|T|RB _DFF_IP1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|6|1 _DFF_IP1_01|6 _DFF_IP1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|6|P _DFF_IP1_01|6|MID_SERIES 0  2e-13
R_DFF_IP1_01|6|B _DFF_IP1_01|6 _DFF_IP1_01|6|MID_SHUNT  2.7439617672
L_DFF_IP1_01|6|RB _DFF_IP1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP1_01|I_1|B _DFF_IP1_01|1 _DFF_IP1_01|I_1|MID  2e-12
I_DFF_IP1_01|I_1|B 0 _DFF_IP1_01|I_1|MID  0.000175
L_DFF_IP1_01|I_3|B _DFF_IP1_01|3 _DFF_IP1_01|I_3|MID  2e-12
I_DFF_IP1_01|I_3|B 0 _DFF_IP1_01|I_3|MID  0.00025
L_DFF_IP1_01|I_T|B _DFF_IP1_01|T1 _DFF_IP1_01|I_T|MID  2e-12
I_DFF_IP1_01|I_T|B 0 _DFF_IP1_01|I_T|MID  0.000175
L_DFF_IP1_01|I_6|B _DFF_IP1_01|6 _DFF_IP1_01|I_6|MID  2e-12
I_DFF_IP1_01|I_6|B 0 _DFF_IP1_01|I_6|MID  0.000175
L_XOR_S1|I_A1|B _XOR_S1|A1 _XOR_S1|I_A1|MID  2e-12
I_XOR_S1|I_A1|B 0 _XOR_S1|I_A1|MID  0.000175
L_XOR_S1|I_A3|B _XOR_S1|A3 _XOR_S1|I_A3|MID  2e-12
I_XOR_S1|I_A3|B 0 _XOR_S1|I_A3|MID  0.000175
L_XOR_S1|I_B1|B _XOR_S1|B1 _XOR_S1|I_B1|MID  2e-12
I_XOR_S1|I_B1|B 0 _XOR_S1|I_B1|MID  0.000175
L_XOR_S1|I_B3|B _XOR_S1|B3 _XOR_S1|I_B3|MID  2e-12
I_XOR_S1|I_B3|B 0 _XOR_S1|I_B3|MID  0.000175
L_XOR_S1|I_T1|B _XOR_S1|T1 _XOR_S1|I_T1|MID  2e-12
I_XOR_S1|I_T1|B 0 _XOR_S1|I_T1|MID  0.000175
L_XOR_S1|I_Q1|B _XOR_S1|Q1 _XOR_S1|I_Q1|MID  2e-12
I_XOR_S1|I_Q1|B 0 _XOR_S1|I_Q1|MID  0.000175
B_XOR_S1|A1|1 _XOR_S1|A1 _XOR_S1|A1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|A1|P _XOR_S1|A1|MID_SERIES 0  5e-13
R_XOR_S1|A1|B _XOR_S1|A1 _XOR_S1|A1|MID_SHUNT  2.7439617672
L_XOR_S1|A1|RB _XOR_S1|A1|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|A2|1 _XOR_S1|A2 _XOR_S1|A2|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|A2|P _XOR_S1|A2|MID_SERIES 0  5e-13
R_XOR_S1|A2|B _XOR_S1|A2 _XOR_S1|A2|MID_SHUNT  2.7439617672
L_XOR_S1|A2|RB _XOR_S1|A2|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|A3|1 _XOR_S1|A2 _XOR_S1|A3|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|A3|P _XOR_S1|A3|MID_SERIES _XOR_S1|A3  1.2e-12
R_XOR_S1|A3|B _XOR_S1|A2 _XOR_S1|A3|MID_SHUNT  2.7439617672
L_XOR_S1|A3|RB _XOR_S1|A3|MID_SHUNT _XOR_S1|A3  2.050338398468e-12
B_XOR_S1|B1|1 _XOR_S1|B1 _XOR_S1|B1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|B1|P _XOR_S1|B1|MID_SERIES 0  5e-13
R_XOR_S1|B1|B _XOR_S1|B1 _XOR_S1|B1|MID_SHUNT  2.7439617672
L_XOR_S1|B1|RB _XOR_S1|B1|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|B2|1 _XOR_S1|B2 _XOR_S1|B2|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|B2|P _XOR_S1|B2|MID_SERIES 0  5e-13
R_XOR_S1|B2|B _XOR_S1|B2 _XOR_S1|B2|MID_SHUNT  2.7439617672
L_XOR_S1|B2|RB _XOR_S1|B2|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|B3|1 _XOR_S1|B2 _XOR_S1|B3|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|B3|P _XOR_S1|B3|MID_SERIES _XOR_S1|B3  1.2e-12
R_XOR_S1|B3|B _XOR_S1|B2 _XOR_S1|B3|MID_SHUNT  2.7439617672
L_XOR_S1|B3|RB _XOR_S1|B3|MID_SHUNT _XOR_S1|B3  2.050338398468e-12
B_XOR_S1|T1|1 _XOR_S1|T1 _XOR_S1|T1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|T1|P _XOR_S1|T1|MID_SERIES 0  5e-13
R_XOR_S1|T1|B _XOR_S1|T1 _XOR_S1|T1|MID_SHUNT  2.7439617672
L_XOR_S1|T1|RB _XOR_S1|T1|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|T2|1 _XOR_S1|T2 _XOR_S1|ABTQ JJMIT AREA=2.0
R_XOR_S1|T2|B _XOR_S1|T2 _XOR_S1|T2|MID_SHUNT  3.429952209
L_XOR_S1|T2|RB _XOR_S1|T2|MID_SHUNT _XOR_S1|ABTQ  2.437922998085e-12
B_XOR_S1|AB|1 _XOR_S1|AB _XOR_S1|AB|MID_SERIES JJMIT AREA=2.0
L_XOR_S1|AB|P _XOR_S1|AB|MID_SERIES _XOR_S1|ABTQ  1.2e-12
R_XOR_S1|AB|B _XOR_S1|AB _XOR_S1|AB|MID_SHUNT  3.429952209
L_XOR_S1|AB|RB _XOR_S1|AB|MID_SHUNT _XOR_S1|ABTQ  2.437922998085e-12
B_XOR_S1|ABTQ|1 _XOR_S1|ABTQ _XOR_S1|ABTQ|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|ABTQ|P _XOR_S1|ABTQ|MID_SERIES 0  5e-13
R_XOR_S1|ABTQ|B _XOR_S1|ABTQ _XOR_S1|ABTQ|MID_SHUNT  2.7439617672
L_XOR_S1|ABTQ|RB _XOR_S1|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_XOR_S1|Q1|1 _XOR_S1|Q1 _XOR_S1|Q1|MID_SERIES JJMIT AREA=2.5
L_XOR_S1|Q1|P _XOR_S1|Q1|MID_SERIES 0  5e-13
R_XOR_S1|Q1|B _XOR_S1|Q1 _XOR_S1|Q1|MID_SHUNT  2.7439617672
L_XOR_S1|Q1|RB _XOR_S1|Q1|MID_SHUNT 0  2.050338398468e-12
B_DFF_IG1_01|1|1 _DFF_IG1_01|1 _DFF_IG1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IG1_01|1|P _DFF_IG1_01|1|MID_SERIES 0  2e-13
R_DFF_IG1_01|1|B _DFF_IG1_01|1 _DFF_IG1_01|1|MID_SHUNT  2.7439617672
L_DFF_IG1_01|1|RB _DFF_IG1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG1_01|23|1 _DFF_IG1_01|2 _DFF_IG1_01|3 JJMIT AREA=1.7857142857142858
R_DFF_IG1_01|23|B _DFF_IG1_01|2 _DFF_IG1_01|23|MID_SHUNT  3.84154647408
L_DFF_IG1_01|23|RB _DFF_IG1_01|23|MID_SHUNT _DFF_IG1_01|3  2.1704737578552e-12
B_DFF_IG1_01|3|1 _DFF_IG1_01|3 _DFF_IG1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IG1_01|3|P _DFF_IG1_01|3|MID_SERIES 0  2e-13
R_DFF_IG1_01|3|B _DFF_IG1_01|3 _DFF_IG1_01|3|MID_SHUNT  2.7439617672
L_DFF_IG1_01|3|RB _DFF_IG1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG1_01|4|1 _DFF_IG1_01|4 _DFF_IG1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IG1_01|4|P _DFF_IG1_01|4|MID_SERIES 0  2e-13
R_DFF_IG1_01|4|B _DFF_IG1_01|4 _DFF_IG1_01|4|MID_SHUNT  2.7439617672
L_DFF_IG1_01|4|RB _DFF_IG1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG1_01|45|1 _DFF_IG1_01|4 _DFF_IG1_01|5 JJMIT AREA=1.7857142857142858
R_DFF_IG1_01|45|B _DFF_IG1_01|4 _DFF_IG1_01|45|MID_SHUNT  3.84154647408
L_DFF_IG1_01|45|RB _DFF_IG1_01|45|MID_SHUNT _DFF_IG1_01|5  2.1704737578552e-12
B_DFF_IG1_01|T|1 _DFF_IG1_01|T1 _DFF_IG1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IG1_01|T|P _DFF_IG1_01|T|MID_SERIES 0  2e-13
R_DFF_IG1_01|T|B _DFF_IG1_01|T1 _DFF_IG1_01|T|MID_SHUNT  2.7439617672
L_DFF_IG1_01|T|RB _DFF_IG1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IG1_01|6|1 _DFF_IG1_01|6 _DFF_IG1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IG1_01|6|P _DFF_IG1_01|6|MID_SERIES 0  2e-13
R_DFF_IG1_01|6|B _DFF_IG1_01|6 _DFF_IG1_01|6|MID_SHUNT  2.7439617672
L_DFF_IG1_01|6|RB _DFF_IG1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IG1_01|I_1|B _DFF_IG1_01|1 _DFF_IG1_01|I_1|MID  2e-12
I_DFF_IG1_01|I_1|B 0 _DFF_IG1_01|I_1|MID  0.000175
L_DFF_IG1_01|I_3|B _DFF_IG1_01|3 _DFF_IG1_01|I_3|MID  2e-12
I_DFF_IG1_01|I_3|B 0 _DFF_IG1_01|I_3|MID  0.00025
L_DFF_IG1_01|I_T|B _DFF_IG1_01|T1 _DFF_IG1_01|I_T|MID  2e-12
I_DFF_IG1_01|I_T|B 0 _DFF_IG1_01|I_T|MID  0.000175
L_DFF_IG1_01|I_6|B _DFF_IG1_01|6 _DFF_IG1_01|I_6|MID  2e-12
I_DFF_IG1_01|I_6|B 0 _DFF_IG1_01|I_6|MID  0.000175
B_DFF_S2|1|1 _DFF_S2|1 _DFF_S2|1|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|1|P _DFF_S2|1|MID_SERIES 0  2e-13
R_DFF_S2|1|B _DFF_S2|1 _DFF_S2|1|MID_SHUNT  2.7439617672
L_DFF_S2|1|RB _DFF_S2|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|23|1 _DFF_S2|2 _DFF_S2|3 JJMIT AREA=1.7857142857142858
R_DFF_S2|23|B _DFF_S2|2 _DFF_S2|23|MID_SHUNT  3.84154647408
L_DFF_S2|23|RB _DFF_S2|23|MID_SHUNT _DFF_S2|3  2.1704737578552e-12
B_DFF_S2|3|1 _DFF_S2|3 _DFF_S2|3|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|3|P _DFF_S2|3|MID_SERIES 0  2e-13
R_DFF_S2|3|B _DFF_S2|3 _DFF_S2|3|MID_SHUNT  2.7439617672
L_DFF_S2|3|RB _DFF_S2|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|4|1 _DFF_S2|4 _DFF_S2|4|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|4|P _DFF_S2|4|MID_SERIES 0  2e-13
R_DFF_S2|4|B _DFF_S2|4 _DFF_S2|4|MID_SHUNT  2.7439617672
L_DFF_S2|4|RB _DFF_S2|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|45|1 _DFF_S2|4 _DFF_S2|5 JJMIT AREA=1.7857142857142858
R_DFF_S2|45|B _DFF_S2|4 _DFF_S2|45|MID_SHUNT  3.84154647408
L_DFF_S2|45|RB _DFF_S2|45|MID_SHUNT _DFF_S2|5  2.1704737578552e-12
B_DFF_S2|T|1 _DFF_S2|T1 _DFF_S2|T|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|T|P _DFF_S2|T|MID_SERIES 0  2e-13
R_DFF_S2|T|B _DFF_S2|T1 _DFF_S2|T|MID_SHUNT  2.7439617672
L_DFF_S2|T|RB _DFF_S2|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_S2|6|1 _DFF_S2|6 _DFF_S2|6|MID_SERIES JJMIT AREA=2.5
L_DFF_S2|6|P _DFF_S2|6|MID_SERIES 0  2e-13
R_DFF_S2|6|B _DFF_S2|6 _DFF_S2|6|MID_SHUNT  2.7439617672
L_DFF_S2|6|RB _DFF_S2|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_S2|I_1|B _DFF_S2|1 _DFF_S2|I_1|MID  2e-12
I_DFF_S2|I_1|B 0 _DFF_S2|I_1|MID  0.000175
L_DFF_S2|I_3|B _DFF_S2|3 _DFF_S2|I_3|MID  2e-12
I_DFF_S2|I_3|B 0 _DFF_S2|I_3|MID  0.00025
L_DFF_S2|I_T|B _DFF_S2|T1 _DFF_S2|I_T|MID  2e-12
I_DFF_S2|I_T|B 0 _DFF_S2|I_T|MID  0.000175
L_DFF_S2|I_6|B _DFF_S2|6 _DFF_S2|I_6|MID  2e-12
I_DFF_S2|I_6|B 0 _DFF_S2|I_6|MID  0.000175
L_INITIAL_0|_SPL_A|I_D1|B _INITIAL_0|_SPL_A|D1 _INITIAL_0|_SPL_A|I_D1|MID  2e-12
I_INITIAL_0|_SPL_A|I_D1|B 0 _INITIAL_0|_SPL_A|I_D1|MID  0.000175
L_INITIAL_0|_SPL_A|I_D2|B _INITIAL_0|_SPL_A|D2 _INITIAL_0|_SPL_A|I_D2|MID  2e-12
I_INITIAL_0|_SPL_A|I_D2|B 0 _INITIAL_0|_SPL_A|I_D2|MID  0.000245
L_INITIAL_0|_SPL_A|I_Q1|B _INITIAL_0|_SPL_A|QA1 _INITIAL_0|_SPL_A|I_Q1|MID  2e-12
I_INITIAL_0|_SPL_A|I_Q1|B 0 _INITIAL_0|_SPL_A|I_Q1|MID  0.000175
L_INITIAL_0|_SPL_A|I_Q2|B _INITIAL_0|_SPL_A|QB1 _INITIAL_0|_SPL_A|I_Q2|MID  2e-12
I_INITIAL_0|_SPL_A|I_Q2|B 0 _INITIAL_0|_SPL_A|I_Q2|MID  0.000175
B_INITIAL_0|_SPL_A|1|1 _INITIAL_0|_SPL_A|D1 _INITIAL_0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_A|1|P _INITIAL_0|_SPL_A|1|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_A|1|B _INITIAL_0|_SPL_A|D1 _INITIAL_0|_SPL_A|1|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_A|1|RB _INITIAL_0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_SPL_A|2|1 _INITIAL_0|_SPL_A|D2 _INITIAL_0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_A|2|P _INITIAL_0|_SPL_A|2|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_A|2|B _INITIAL_0|_SPL_A|D2 _INITIAL_0|_SPL_A|2|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_A|2|RB _INITIAL_0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_SPL_A|A|1 _INITIAL_0|_SPL_A|QA1 _INITIAL_0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_A|A|P _INITIAL_0|_SPL_A|A|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_A|A|B _INITIAL_0|_SPL_A|QA1 _INITIAL_0|_SPL_A|A|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_A|A|RB _INITIAL_0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_SPL_A|B|1 _INITIAL_0|_SPL_A|QB1 _INITIAL_0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_A|B|P _INITIAL_0|_SPL_A|B|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_A|B|B _INITIAL_0|_SPL_A|QB1 _INITIAL_0|_SPL_A|B|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_A|B|RB _INITIAL_0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_0|_SPL_B|I_D1|B _INITIAL_0|_SPL_B|D1 _INITIAL_0|_SPL_B|I_D1|MID  2e-12
I_INITIAL_0|_SPL_B|I_D1|B 0 _INITIAL_0|_SPL_B|I_D1|MID  0.000175
L_INITIAL_0|_SPL_B|I_D2|B _INITIAL_0|_SPL_B|D2 _INITIAL_0|_SPL_B|I_D2|MID  2e-12
I_INITIAL_0|_SPL_B|I_D2|B 0 _INITIAL_0|_SPL_B|I_D2|MID  0.000245
L_INITIAL_0|_SPL_B|I_Q1|B _INITIAL_0|_SPL_B|QA1 _INITIAL_0|_SPL_B|I_Q1|MID  2e-12
I_INITIAL_0|_SPL_B|I_Q1|B 0 _INITIAL_0|_SPL_B|I_Q1|MID  0.000175
L_INITIAL_0|_SPL_B|I_Q2|B _INITIAL_0|_SPL_B|QB1 _INITIAL_0|_SPL_B|I_Q2|MID  2e-12
I_INITIAL_0|_SPL_B|I_Q2|B 0 _INITIAL_0|_SPL_B|I_Q2|MID  0.000175
B_INITIAL_0|_SPL_B|1|1 _INITIAL_0|_SPL_B|D1 _INITIAL_0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_B|1|P _INITIAL_0|_SPL_B|1|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_B|1|B _INITIAL_0|_SPL_B|D1 _INITIAL_0|_SPL_B|1|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_B|1|RB _INITIAL_0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_SPL_B|2|1 _INITIAL_0|_SPL_B|D2 _INITIAL_0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_B|2|P _INITIAL_0|_SPL_B|2|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_B|2|B _INITIAL_0|_SPL_B|D2 _INITIAL_0|_SPL_B|2|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_B|2|RB _INITIAL_0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_SPL_B|A|1 _INITIAL_0|_SPL_B|QA1 _INITIAL_0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_B|A|P _INITIAL_0|_SPL_B|A|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_B|A|B _INITIAL_0|_SPL_B|QA1 _INITIAL_0|_SPL_B|A|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_B|A|RB _INITIAL_0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_SPL_B|B|1 _INITIAL_0|_SPL_B|QB1 _INITIAL_0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_SPL_B|B|P _INITIAL_0|_SPL_B|B|MID_SERIES 0  2e-13
R_INITIAL_0|_SPL_B|B|B _INITIAL_0|_SPL_B|QB1 _INITIAL_0|_SPL_B|B|MID_SHUNT  2.7439617672
L_INITIAL_0|_SPL_B|B|RB _INITIAL_0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_A|1|1 _INITIAL_0|_DFF_A|1 _INITIAL_0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_A|1|P _INITIAL_0|_DFF_A|1|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_A|1|B _INITIAL_0|_DFF_A|1 _INITIAL_0|_DFF_A|1|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_A|1|RB _INITIAL_0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_A|23|1 _INITIAL_0|_DFF_A|2 _INITIAL_0|_DFF_A|3 JJMIT AREA=1.7857142857142858
R_INITIAL_0|_DFF_A|23|B _INITIAL_0|_DFF_A|2 _INITIAL_0|_DFF_A|23|MID_SHUNT  3.84154647408
L_INITIAL_0|_DFF_A|23|RB _INITIAL_0|_DFF_A|23|MID_SHUNT _INITIAL_0|_DFF_A|3  2.1704737578552e-12
B_INITIAL_0|_DFF_A|3|1 _INITIAL_0|_DFF_A|3 _INITIAL_0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_A|3|P _INITIAL_0|_DFF_A|3|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_A|3|B _INITIAL_0|_DFF_A|3 _INITIAL_0|_DFF_A|3|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_A|3|RB _INITIAL_0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_A|4|1 _INITIAL_0|_DFF_A|4 _INITIAL_0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_A|4|P _INITIAL_0|_DFF_A|4|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_A|4|B _INITIAL_0|_DFF_A|4 _INITIAL_0|_DFF_A|4|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_A|4|RB _INITIAL_0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_A|45|1 _INITIAL_0|_DFF_A|4 _INITIAL_0|_DFF_A|5 JJMIT AREA=1.7857142857142858
R_INITIAL_0|_DFF_A|45|B _INITIAL_0|_DFF_A|4 _INITIAL_0|_DFF_A|45|MID_SHUNT  3.84154647408
L_INITIAL_0|_DFF_A|45|RB _INITIAL_0|_DFF_A|45|MID_SHUNT _INITIAL_0|_DFF_A|5  2.1704737578552e-12
B_INITIAL_0|_DFF_A|T|1 _INITIAL_0|_DFF_A|T1 _INITIAL_0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_A|T|P _INITIAL_0|_DFF_A|T|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_A|T|B _INITIAL_0|_DFF_A|T1 _INITIAL_0|_DFF_A|T|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_A|T|RB _INITIAL_0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_A|6|1 _INITIAL_0|_DFF_A|6 _INITIAL_0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_A|6|P _INITIAL_0|_DFF_A|6|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_A|6|B _INITIAL_0|_DFF_A|6 _INITIAL_0|_DFF_A|6|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_A|6|RB _INITIAL_0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_0|_DFF_A|I_1|B _INITIAL_0|_DFF_A|1 _INITIAL_0|_DFF_A|I_1|MID  2e-12
I_INITIAL_0|_DFF_A|I_1|B 0 _INITIAL_0|_DFF_A|I_1|MID  0.000175
L_INITIAL_0|_DFF_A|I_3|B _INITIAL_0|_DFF_A|3 _INITIAL_0|_DFF_A|I_3|MID  2e-12
I_INITIAL_0|_DFF_A|I_3|B 0 _INITIAL_0|_DFF_A|I_3|MID  0.00025
L_INITIAL_0|_DFF_A|I_T|B _INITIAL_0|_DFF_A|T1 _INITIAL_0|_DFF_A|I_T|MID  2e-12
I_INITIAL_0|_DFF_A|I_T|B 0 _INITIAL_0|_DFF_A|I_T|MID  0.000175
L_INITIAL_0|_DFF_A|I_6|B _INITIAL_0|_DFF_A|6 _INITIAL_0|_DFF_A|I_6|MID  2e-12
I_INITIAL_0|_DFF_A|I_6|B 0 _INITIAL_0|_DFF_A|I_6|MID  0.000175
B_INITIAL_0|_DFF_B|1|1 _INITIAL_0|_DFF_B|1 _INITIAL_0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_B|1|P _INITIAL_0|_DFF_B|1|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_B|1|B _INITIAL_0|_DFF_B|1 _INITIAL_0|_DFF_B|1|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_B|1|RB _INITIAL_0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_B|23|1 _INITIAL_0|_DFF_B|2 _INITIAL_0|_DFF_B|3 JJMIT AREA=1.7857142857142858
R_INITIAL_0|_DFF_B|23|B _INITIAL_0|_DFF_B|2 _INITIAL_0|_DFF_B|23|MID_SHUNT  3.84154647408
L_INITIAL_0|_DFF_B|23|RB _INITIAL_0|_DFF_B|23|MID_SHUNT _INITIAL_0|_DFF_B|3  2.1704737578552e-12
B_INITIAL_0|_DFF_B|3|1 _INITIAL_0|_DFF_B|3 _INITIAL_0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_B|3|P _INITIAL_0|_DFF_B|3|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_B|3|B _INITIAL_0|_DFF_B|3 _INITIAL_0|_DFF_B|3|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_B|3|RB _INITIAL_0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_B|4|1 _INITIAL_0|_DFF_B|4 _INITIAL_0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_B|4|P _INITIAL_0|_DFF_B|4|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_B|4|B _INITIAL_0|_DFF_B|4 _INITIAL_0|_DFF_B|4|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_B|4|RB _INITIAL_0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_B|45|1 _INITIAL_0|_DFF_B|4 _INITIAL_0|_DFF_B|5 JJMIT AREA=1.7857142857142858
R_INITIAL_0|_DFF_B|45|B _INITIAL_0|_DFF_B|4 _INITIAL_0|_DFF_B|45|MID_SHUNT  3.84154647408
L_INITIAL_0|_DFF_B|45|RB _INITIAL_0|_DFF_B|45|MID_SHUNT _INITIAL_0|_DFF_B|5  2.1704737578552e-12
B_INITIAL_0|_DFF_B|T|1 _INITIAL_0|_DFF_B|T1 _INITIAL_0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_B|T|P _INITIAL_0|_DFF_B|T|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_B|T|B _INITIAL_0|_DFF_B|T1 _INITIAL_0|_DFF_B|T|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_B|T|RB _INITIAL_0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_DFF_B|6|1 _INITIAL_0|_DFF_B|6 _INITIAL_0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_DFF_B|6|P _INITIAL_0|_DFF_B|6|MID_SERIES 0  2e-13
R_INITIAL_0|_DFF_B|6|B _INITIAL_0|_DFF_B|6 _INITIAL_0|_DFF_B|6|MID_SHUNT  2.7439617672
L_INITIAL_0|_DFF_B|6|RB _INITIAL_0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_0|_DFF_B|I_1|B _INITIAL_0|_DFF_B|1 _INITIAL_0|_DFF_B|I_1|MID  2e-12
I_INITIAL_0|_DFF_B|I_1|B 0 _INITIAL_0|_DFF_B|I_1|MID  0.000175
L_INITIAL_0|_DFF_B|I_3|B _INITIAL_0|_DFF_B|3 _INITIAL_0|_DFF_B|I_3|MID  2e-12
I_INITIAL_0|_DFF_B|I_3|B 0 _INITIAL_0|_DFF_B|I_3|MID  0.00025
L_INITIAL_0|_DFF_B|I_T|B _INITIAL_0|_DFF_B|T1 _INITIAL_0|_DFF_B|I_T|MID  2e-12
I_INITIAL_0|_DFF_B|I_T|B 0 _INITIAL_0|_DFF_B|I_T|MID  0.000175
L_INITIAL_0|_DFF_B|I_6|B _INITIAL_0|_DFF_B|6 _INITIAL_0|_DFF_B|I_6|MID  2e-12
I_INITIAL_0|_DFF_B|I_6|B 0 _INITIAL_0|_DFF_B|I_6|MID  0.000175
L_INITIAL_0|_XOR|I_A1|B _INITIAL_0|_XOR|A1 _INITIAL_0|_XOR|I_A1|MID  2e-12
I_INITIAL_0|_XOR|I_A1|B 0 _INITIAL_0|_XOR|I_A1|MID  0.000175
L_INITIAL_0|_XOR|I_A3|B _INITIAL_0|_XOR|A3 _INITIAL_0|_XOR|I_A3|MID  2e-12
I_INITIAL_0|_XOR|I_A3|B 0 _INITIAL_0|_XOR|I_A3|MID  0.000175
L_INITIAL_0|_XOR|I_B1|B _INITIAL_0|_XOR|B1 _INITIAL_0|_XOR|I_B1|MID  2e-12
I_INITIAL_0|_XOR|I_B1|B 0 _INITIAL_0|_XOR|I_B1|MID  0.000175
L_INITIAL_0|_XOR|I_B3|B _INITIAL_0|_XOR|B3 _INITIAL_0|_XOR|I_B3|MID  2e-12
I_INITIAL_0|_XOR|I_B3|B 0 _INITIAL_0|_XOR|I_B3|MID  0.000175
L_INITIAL_0|_XOR|I_T1|B _INITIAL_0|_XOR|T1 _INITIAL_0|_XOR|I_T1|MID  2e-12
I_INITIAL_0|_XOR|I_T1|B 0 _INITIAL_0|_XOR|I_T1|MID  0.000175
L_INITIAL_0|_XOR|I_Q1|B _INITIAL_0|_XOR|Q1 _INITIAL_0|_XOR|I_Q1|MID  2e-12
I_INITIAL_0|_XOR|I_Q1|B 0 _INITIAL_0|_XOR|I_Q1|MID  0.000175
B_INITIAL_0|_XOR|A1|1 _INITIAL_0|_XOR|A1 _INITIAL_0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|A1|P _INITIAL_0|_XOR|A1|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|A1|B _INITIAL_0|_XOR|A1 _INITIAL_0|_XOR|A1|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|A1|RB _INITIAL_0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_0|_XOR|A2|1 _INITIAL_0|_XOR|A2 _INITIAL_0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|A2|P _INITIAL_0|_XOR|A2|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|A2|B _INITIAL_0|_XOR|A2 _INITIAL_0|_XOR|A2|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|A2|RB _INITIAL_0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_0|_XOR|A3|1 _INITIAL_0|_XOR|A2 _INITIAL_0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|A3|P _INITIAL_0|_XOR|A3|MID_SERIES _INITIAL_0|_XOR|A3  1.2e-12
R_INITIAL_0|_XOR|A3|B _INITIAL_0|_XOR|A2 _INITIAL_0|_XOR|A3|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|A3|RB _INITIAL_0|_XOR|A3|MID_SHUNT _INITIAL_0|_XOR|A3  2.050338398468e-12
B_INITIAL_0|_XOR|B1|1 _INITIAL_0|_XOR|B1 _INITIAL_0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|B1|P _INITIAL_0|_XOR|B1|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|B1|B _INITIAL_0|_XOR|B1 _INITIAL_0|_XOR|B1|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|B1|RB _INITIAL_0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_0|_XOR|B2|1 _INITIAL_0|_XOR|B2 _INITIAL_0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|B2|P _INITIAL_0|_XOR|B2|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|B2|B _INITIAL_0|_XOR|B2 _INITIAL_0|_XOR|B2|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|B2|RB _INITIAL_0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_0|_XOR|B3|1 _INITIAL_0|_XOR|B2 _INITIAL_0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|B3|P _INITIAL_0|_XOR|B3|MID_SERIES _INITIAL_0|_XOR|B3  1.2e-12
R_INITIAL_0|_XOR|B3|B _INITIAL_0|_XOR|B2 _INITIAL_0|_XOR|B3|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|B3|RB _INITIAL_0|_XOR|B3|MID_SHUNT _INITIAL_0|_XOR|B3  2.050338398468e-12
B_INITIAL_0|_XOR|T1|1 _INITIAL_0|_XOR|T1 _INITIAL_0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|T1|P _INITIAL_0|_XOR|T1|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|T1|B _INITIAL_0|_XOR|T1 _INITIAL_0|_XOR|T1|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|T1|RB _INITIAL_0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_0|_XOR|T2|1 _INITIAL_0|_XOR|T2 _INITIAL_0|_XOR|ABTQ JJMIT AREA=2.0
R_INITIAL_0|_XOR|T2|B _INITIAL_0|_XOR|T2 _INITIAL_0|_XOR|T2|MID_SHUNT  3.429952209
L_INITIAL_0|_XOR|T2|RB _INITIAL_0|_XOR|T2|MID_SHUNT _INITIAL_0|_XOR|ABTQ  2.437922998085e-12
B_INITIAL_0|_XOR|AB|1 _INITIAL_0|_XOR|AB _INITIAL_0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
L_INITIAL_0|_XOR|AB|P _INITIAL_0|_XOR|AB|MID_SERIES _INITIAL_0|_XOR|ABTQ  1.2e-12
R_INITIAL_0|_XOR|AB|B _INITIAL_0|_XOR|AB _INITIAL_0|_XOR|AB|MID_SHUNT  3.429952209
L_INITIAL_0|_XOR|AB|RB _INITIAL_0|_XOR|AB|MID_SHUNT _INITIAL_0|_XOR|ABTQ  2.437922998085e-12
B_INITIAL_0|_XOR|ABTQ|1 _INITIAL_0|_XOR|ABTQ _INITIAL_0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|ABTQ|P _INITIAL_0|_XOR|ABTQ|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|ABTQ|B _INITIAL_0|_XOR|ABTQ _INITIAL_0|_XOR|ABTQ|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|ABTQ|RB _INITIAL_0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_0|_XOR|Q1|1 _INITIAL_0|_XOR|Q1 _INITIAL_0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_XOR|Q1|P _INITIAL_0|_XOR|Q1|MID_SERIES 0  5e-13
R_INITIAL_0|_XOR|Q1|B _INITIAL_0|_XOR|Q1 _INITIAL_0|_XOR|Q1|MID_SHUNT  2.7439617672
L_INITIAL_0|_XOR|Q1|RB _INITIAL_0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
L_INITIAL_0|_AND|I_A1|B _INITIAL_0|_AND|A1 _INITIAL_0|_AND|I_A1|MID  2e-12
I_INITIAL_0|_AND|I_A1|B 0 _INITIAL_0|_AND|I_A1|MID  0.000175
L_INITIAL_0|_AND|I_B1|B _INITIAL_0|_AND|B1 _INITIAL_0|_AND|I_B1|MID  2e-12
I_INITIAL_0|_AND|I_B1|B 0 _INITIAL_0|_AND|I_B1|MID  0.000175
L_INITIAL_0|_AND|I_Q3|B _INITIAL_0|_AND|Q3 _INITIAL_0|_AND|I_Q3|MID  2e-12
I_INITIAL_0|_AND|I_Q3|B 0 _INITIAL_0|_AND|I_Q3|MID  5e-05
L_INITIAL_0|_AND|I_Q2|B _INITIAL_0|_AND|Q2 _INITIAL_0|_AND|I_Q2|MID  2e-12
I_INITIAL_0|_AND|I_Q2|B 0 _INITIAL_0|_AND|I_Q2|MID  0.000175
L_INITIAL_0|_AND|I_Q1|B _INITIAL_0|_AND|Q1 _INITIAL_0|_AND|I_Q1|MID  2e-12
I_INITIAL_0|_AND|I_Q1|B 0 _INITIAL_0|_AND|I_Q1|MID  0.000175
B_INITIAL_0|_AND|A1|1 _INITIAL_0|_AND|A1 _INITIAL_0|_AND|A1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_AND|A1|P _INITIAL_0|_AND|A1|MID_SERIES 0  2e-13
R_INITIAL_0|_AND|A1|B _INITIAL_0|_AND|A1 _INITIAL_0|_AND|A1|MID_SHUNT  2.7439617672
L_INITIAL_0|_AND|A1|RB _INITIAL_0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_AND|A2|1 _INITIAL_0|_AND|A2 _INITIAL_0|_AND|A2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_AND|A2|P _INITIAL_0|_AND|A2|MID_SERIES 0  2e-13
R_INITIAL_0|_AND|A2|B _INITIAL_0|_AND|A2 _INITIAL_0|_AND|A2|MID_SHUNT  2.7439617672
L_INITIAL_0|_AND|A2|RB _INITIAL_0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_AND|A12|1 _INITIAL_0|_AND|A2 _INITIAL_0|_AND|A3 JJMIT AREA=1.7857142857142858
R_INITIAL_0|_AND|A12|B _INITIAL_0|_AND|A2 _INITIAL_0|_AND|A12|MID_SHUNT  3.84154647408
L_INITIAL_0|_AND|A12|RB _INITIAL_0|_AND|A12|MID_SHUNT _INITIAL_0|_AND|A3  2.1704737578552e-12
B_INITIAL_0|_AND|B1|1 _INITIAL_0|_AND|B1 _INITIAL_0|_AND|B1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_AND|B1|P _INITIAL_0|_AND|B1|MID_SERIES 0  2e-13
R_INITIAL_0|_AND|B1|B _INITIAL_0|_AND|B1 _INITIAL_0|_AND|B1|MID_SHUNT  2.7439617672
L_INITIAL_0|_AND|B1|RB _INITIAL_0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_AND|B2|1 _INITIAL_0|_AND|B2 _INITIAL_0|_AND|B2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_AND|B2|P _INITIAL_0|_AND|B2|MID_SERIES 0  2e-13
R_INITIAL_0|_AND|B2|B _INITIAL_0|_AND|B2 _INITIAL_0|_AND|B2|MID_SHUNT  2.7439617672
L_INITIAL_0|_AND|B2|RB _INITIAL_0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_AND|B12|1 _INITIAL_0|_AND|B2 _INITIAL_0|_AND|B3 JJMIT AREA=1.7857142857142858
R_INITIAL_0|_AND|B12|B _INITIAL_0|_AND|B2 _INITIAL_0|_AND|B12|MID_SHUNT  3.84154647408
L_INITIAL_0|_AND|B12|RB _INITIAL_0|_AND|B12|MID_SHUNT _INITIAL_0|_AND|B3  2.1704737578552e-12
B_INITIAL_0|_AND|Q2|1 _INITIAL_0|_AND|Q2 _INITIAL_0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_AND|Q2|P _INITIAL_0|_AND|Q2|MID_SERIES 0  2e-13
R_INITIAL_0|_AND|Q2|B _INITIAL_0|_AND|Q2 _INITIAL_0|_AND|Q2|MID_SHUNT  2.7439617672
L_INITIAL_0|_AND|Q2|RB _INITIAL_0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_0|_AND|Q1|1 _INITIAL_0|_AND|Q1 _INITIAL_0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_0|_AND|Q1|P _INITIAL_0|_AND|Q1|MID_SERIES 0  2e-13
R_INITIAL_0|_AND|Q1|B _INITIAL_0|_AND|Q1 _INITIAL_0|_AND|Q1|MID_SHUNT  2.7439617672
L_INITIAL_0|_AND|Q1|RB _INITIAL_0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_1|_SPL_A|I_D1|B _INITIAL_1|_SPL_A|D1 _INITIAL_1|_SPL_A|I_D1|MID  2e-12
I_INITIAL_1|_SPL_A|I_D1|B 0 _INITIAL_1|_SPL_A|I_D1|MID  0.000175
L_INITIAL_1|_SPL_A|I_D2|B _INITIAL_1|_SPL_A|D2 _INITIAL_1|_SPL_A|I_D2|MID  2e-12
I_INITIAL_1|_SPL_A|I_D2|B 0 _INITIAL_1|_SPL_A|I_D2|MID  0.000245
L_INITIAL_1|_SPL_A|I_Q1|B _INITIAL_1|_SPL_A|QA1 _INITIAL_1|_SPL_A|I_Q1|MID  2e-12
I_INITIAL_1|_SPL_A|I_Q1|B 0 _INITIAL_1|_SPL_A|I_Q1|MID  0.000175
L_INITIAL_1|_SPL_A|I_Q2|B _INITIAL_1|_SPL_A|QB1 _INITIAL_1|_SPL_A|I_Q2|MID  2e-12
I_INITIAL_1|_SPL_A|I_Q2|B 0 _INITIAL_1|_SPL_A|I_Q2|MID  0.000175
B_INITIAL_1|_SPL_A|1|1 _INITIAL_1|_SPL_A|D1 _INITIAL_1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_A|1|P _INITIAL_1|_SPL_A|1|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_A|1|B _INITIAL_1|_SPL_A|D1 _INITIAL_1|_SPL_A|1|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_A|1|RB _INITIAL_1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_SPL_A|2|1 _INITIAL_1|_SPL_A|D2 _INITIAL_1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_A|2|P _INITIAL_1|_SPL_A|2|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_A|2|B _INITIAL_1|_SPL_A|D2 _INITIAL_1|_SPL_A|2|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_A|2|RB _INITIAL_1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_SPL_A|A|1 _INITIAL_1|_SPL_A|QA1 _INITIAL_1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_A|A|P _INITIAL_1|_SPL_A|A|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_A|A|B _INITIAL_1|_SPL_A|QA1 _INITIAL_1|_SPL_A|A|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_A|A|RB _INITIAL_1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_SPL_A|B|1 _INITIAL_1|_SPL_A|QB1 _INITIAL_1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_A|B|P _INITIAL_1|_SPL_A|B|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_A|B|B _INITIAL_1|_SPL_A|QB1 _INITIAL_1|_SPL_A|B|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_A|B|RB _INITIAL_1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_1|_SPL_B|I_D1|B _INITIAL_1|_SPL_B|D1 _INITIAL_1|_SPL_B|I_D1|MID  2e-12
I_INITIAL_1|_SPL_B|I_D1|B 0 _INITIAL_1|_SPL_B|I_D1|MID  0.000175
L_INITIAL_1|_SPL_B|I_D2|B _INITIAL_1|_SPL_B|D2 _INITIAL_1|_SPL_B|I_D2|MID  2e-12
I_INITIAL_1|_SPL_B|I_D2|B 0 _INITIAL_1|_SPL_B|I_D2|MID  0.000245
L_INITIAL_1|_SPL_B|I_Q1|B _INITIAL_1|_SPL_B|QA1 _INITIAL_1|_SPL_B|I_Q1|MID  2e-12
I_INITIAL_1|_SPL_B|I_Q1|B 0 _INITIAL_1|_SPL_B|I_Q1|MID  0.000175
L_INITIAL_1|_SPL_B|I_Q2|B _INITIAL_1|_SPL_B|QB1 _INITIAL_1|_SPL_B|I_Q2|MID  2e-12
I_INITIAL_1|_SPL_B|I_Q2|B 0 _INITIAL_1|_SPL_B|I_Q2|MID  0.000175
B_INITIAL_1|_SPL_B|1|1 _INITIAL_1|_SPL_B|D1 _INITIAL_1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_B|1|P _INITIAL_1|_SPL_B|1|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_B|1|B _INITIAL_1|_SPL_B|D1 _INITIAL_1|_SPL_B|1|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_B|1|RB _INITIAL_1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_SPL_B|2|1 _INITIAL_1|_SPL_B|D2 _INITIAL_1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_B|2|P _INITIAL_1|_SPL_B|2|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_B|2|B _INITIAL_1|_SPL_B|D2 _INITIAL_1|_SPL_B|2|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_B|2|RB _INITIAL_1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_SPL_B|A|1 _INITIAL_1|_SPL_B|QA1 _INITIAL_1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_B|A|P _INITIAL_1|_SPL_B|A|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_B|A|B _INITIAL_1|_SPL_B|QA1 _INITIAL_1|_SPL_B|A|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_B|A|RB _INITIAL_1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_SPL_B|B|1 _INITIAL_1|_SPL_B|QB1 _INITIAL_1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_SPL_B|B|P _INITIAL_1|_SPL_B|B|MID_SERIES 0  2e-13
R_INITIAL_1|_SPL_B|B|B _INITIAL_1|_SPL_B|QB1 _INITIAL_1|_SPL_B|B|MID_SHUNT  2.7439617672
L_INITIAL_1|_SPL_B|B|RB _INITIAL_1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_A|1|1 _INITIAL_1|_DFF_A|1 _INITIAL_1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_A|1|P _INITIAL_1|_DFF_A|1|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_A|1|B _INITIAL_1|_DFF_A|1 _INITIAL_1|_DFF_A|1|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_A|1|RB _INITIAL_1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_A|23|1 _INITIAL_1|_DFF_A|2 _INITIAL_1|_DFF_A|3 JJMIT AREA=1.7857142857142858
R_INITIAL_1|_DFF_A|23|B _INITIAL_1|_DFF_A|2 _INITIAL_1|_DFF_A|23|MID_SHUNT  3.84154647408
L_INITIAL_1|_DFF_A|23|RB _INITIAL_1|_DFF_A|23|MID_SHUNT _INITIAL_1|_DFF_A|3  2.1704737578552e-12
B_INITIAL_1|_DFF_A|3|1 _INITIAL_1|_DFF_A|3 _INITIAL_1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_A|3|P _INITIAL_1|_DFF_A|3|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_A|3|B _INITIAL_1|_DFF_A|3 _INITIAL_1|_DFF_A|3|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_A|3|RB _INITIAL_1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_A|4|1 _INITIAL_1|_DFF_A|4 _INITIAL_1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_A|4|P _INITIAL_1|_DFF_A|4|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_A|4|B _INITIAL_1|_DFF_A|4 _INITIAL_1|_DFF_A|4|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_A|4|RB _INITIAL_1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_A|45|1 _INITIAL_1|_DFF_A|4 _INITIAL_1|_DFF_A|5 JJMIT AREA=1.7857142857142858
R_INITIAL_1|_DFF_A|45|B _INITIAL_1|_DFF_A|4 _INITIAL_1|_DFF_A|45|MID_SHUNT  3.84154647408
L_INITIAL_1|_DFF_A|45|RB _INITIAL_1|_DFF_A|45|MID_SHUNT _INITIAL_1|_DFF_A|5  2.1704737578552e-12
B_INITIAL_1|_DFF_A|T|1 _INITIAL_1|_DFF_A|T1 _INITIAL_1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_A|T|P _INITIAL_1|_DFF_A|T|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_A|T|B _INITIAL_1|_DFF_A|T1 _INITIAL_1|_DFF_A|T|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_A|T|RB _INITIAL_1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_A|6|1 _INITIAL_1|_DFF_A|6 _INITIAL_1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_A|6|P _INITIAL_1|_DFF_A|6|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_A|6|B _INITIAL_1|_DFF_A|6 _INITIAL_1|_DFF_A|6|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_A|6|RB _INITIAL_1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_1|_DFF_A|I_1|B _INITIAL_1|_DFF_A|1 _INITIAL_1|_DFF_A|I_1|MID  2e-12
I_INITIAL_1|_DFF_A|I_1|B 0 _INITIAL_1|_DFF_A|I_1|MID  0.000175
L_INITIAL_1|_DFF_A|I_3|B _INITIAL_1|_DFF_A|3 _INITIAL_1|_DFF_A|I_3|MID  2e-12
I_INITIAL_1|_DFF_A|I_3|B 0 _INITIAL_1|_DFF_A|I_3|MID  0.00025
L_INITIAL_1|_DFF_A|I_T|B _INITIAL_1|_DFF_A|T1 _INITIAL_1|_DFF_A|I_T|MID  2e-12
I_INITIAL_1|_DFF_A|I_T|B 0 _INITIAL_1|_DFF_A|I_T|MID  0.000175
L_INITIAL_1|_DFF_A|I_6|B _INITIAL_1|_DFF_A|6 _INITIAL_1|_DFF_A|I_6|MID  2e-12
I_INITIAL_1|_DFF_A|I_6|B 0 _INITIAL_1|_DFF_A|I_6|MID  0.000175
B_INITIAL_1|_DFF_B|1|1 _INITIAL_1|_DFF_B|1 _INITIAL_1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_B|1|P _INITIAL_1|_DFF_B|1|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_B|1|B _INITIAL_1|_DFF_B|1 _INITIAL_1|_DFF_B|1|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_B|1|RB _INITIAL_1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_B|23|1 _INITIAL_1|_DFF_B|2 _INITIAL_1|_DFF_B|3 JJMIT AREA=1.7857142857142858
R_INITIAL_1|_DFF_B|23|B _INITIAL_1|_DFF_B|2 _INITIAL_1|_DFF_B|23|MID_SHUNT  3.84154647408
L_INITIAL_1|_DFF_B|23|RB _INITIAL_1|_DFF_B|23|MID_SHUNT _INITIAL_1|_DFF_B|3  2.1704737578552e-12
B_INITIAL_1|_DFF_B|3|1 _INITIAL_1|_DFF_B|3 _INITIAL_1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_B|3|P _INITIAL_1|_DFF_B|3|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_B|3|B _INITIAL_1|_DFF_B|3 _INITIAL_1|_DFF_B|3|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_B|3|RB _INITIAL_1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_B|4|1 _INITIAL_1|_DFF_B|4 _INITIAL_1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_B|4|P _INITIAL_1|_DFF_B|4|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_B|4|B _INITIAL_1|_DFF_B|4 _INITIAL_1|_DFF_B|4|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_B|4|RB _INITIAL_1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_B|45|1 _INITIAL_1|_DFF_B|4 _INITIAL_1|_DFF_B|5 JJMIT AREA=1.7857142857142858
R_INITIAL_1|_DFF_B|45|B _INITIAL_1|_DFF_B|4 _INITIAL_1|_DFF_B|45|MID_SHUNT  3.84154647408
L_INITIAL_1|_DFF_B|45|RB _INITIAL_1|_DFF_B|45|MID_SHUNT _INITIAL_1|_DFF_B|5  2.1704737578552e-12
B_INITIAL_1|_DFF_B|T|1 _INITIAL_1|_DFF_B|T1 _INITIAL_1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_B|T|P _INITIAL_1|_DFF_B|T|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_B|T|B _INITIAL_1|_DFF_B|T1 _INITIAL_1|_DFF_B|T|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_B|T|RB _INITIAL_1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_DFF_B|6|1 _INITIAL_1|_DFF_B|6 _INITIAL_1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_DFF_B|6|P _INITIAL_1|_DFF_B|6|MID_SERIES 0  2e-13
R_INITIAL_1|_DFF_B|6|B _INITIAL_1|_DFF_B|6 _INITIAL_1|_DFF_B|6|MID_SHUNT  2.7439617672
L_INITIAL_1|_DFF_B|6|RB _INITIAL_1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
L_INITIAL_1|_DFF_B|I_1|B _INITIAL_1|_DFF_B|1 _INITIAL_1|_DFF_B|I_1|MID  2e-12
I_INITIAL_1|_DFF_B|I_1|B 0 _INITIAL_1|_DFF_B|I_1|MID  0.000175
L_INITIAL_1|_DFF_B|I_3|B _INITIAL_1|_DFF_B|3 _INITIAL_1|_DFF_B|I_3|MID  2e-12
I_INITIAL_1|_DFF_B|I_3|B 0 _INITIAL_1|_DFF_B|I_3|MID  0.00025
L_INITIAL_1|_DFF_B|I_T|B _INITIAL_1|_DFF_B|T1 _INITIAL_1|_DFF_B|I_T|MID  2e-12
I_INITIAL_1|_DFF_B|I_T|B 0 _INITIAL_1|_DFF_B|I_T|MID  0.000175
L_INITIAL_1|_DFF_B|I_6|B _INITIAL_1|_DFF_B|6 _INITIAL_1|_DFF_B|I_6|MID  2e-12
I_INITIAL_1|_DFF_B|I_6|B 0 _INITIAL_1|_DFF_B|I_6|MID  0.000175
L_INITIAL_1|_XOR|I_A1|B _INITIAL_1|_XOR|A1 _INITIAL_1|_XOR|I_A1|MID  2e-12
I_INITIAL_1|_XOR|I_A1|B 0 _INITIAL_1|_XOR|I_A1|MID  0.000175
L_INITIAL_1|_XOR|I_A3|B _INITIAL_1|_XOR|A3 _INITIAL_1|_XOR|I_A3|MID  2e-12
I_INITIAL_1|_XOR|I_A3|B 0 _INITIAL_1|_XOR|I_A3|MID  0.000175
L_INITIAL_1|_XOR|I_B1|B _INITIAL_1|_XOR|B1 _INITIAL_1|_XOR|I_B1|MID  2e-12
I_INITIAL_1|_XOR|I_B1|B 0 _INITIAL_1|_XOR|I_B1|MID  0.000175
L_INITIAL_1|_XOR|I_B3|B _INITIAL_1|_XOR|B3 _INITIAL_1|_XOR|I_B3|MID  2e-12
I_INITIAL_1|_XOR|I_B3|B 0 _INITIAL_1|_XOR|I_B3|MID  0.000175
L_INITIAL_1|_XOR|I_T1|B _INITIAL_1|_XOR|T1 _INITIAL_1|_XOR|I_T1|MID  2e-12
I_INITIAL_1|_XOR|I_T1|B 0 _INITIAL_1|_XOR|I_T1|MID  0.000175
L_INITIAL_1|_XOR|I_Q1|B _INITIAL_1|_XOR|Q1 _INITIAL_1|_XOR|I_Q1|MID  2e-12
I_INITIAL_1|_XOR|I_Q1|B 0 _INITIAL_1|_XOR|I_Q1|MID  0.000175
B_INITIAL_1|_XOR|A1|1 _INITIAL_1|_XOR|A1 _INITIAL_1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|A1|P _INITIAL_1|_XOR|A1|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|A1|B _INITIAL_1|_XOR|A1 _INITIAL_1|_XOR|A1|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|A1|RB _INITIAL_1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_1|_XOR|A2|1 _INITIAL_1|_XOR|A2 _INITIAL_1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|A2|P _INITIAL_1|_XOR|A2|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|A2|B _INITIAL_1|_XOR|A2 _INITIAL_1|_XOR|A2|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|A2|RB _INITIAL_1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_1|_XOR|A3|1 _INITIAL_1|_XOR|A2 _INITIAL_1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|A3|P _INITIAL_1|_XOR|A3|MID_SERIES _INITIAL_1|_XOR|A3  1.2e-12
R_INITIAL_1|_XOR|A3|B _INITIAL_1|_XOR|A2 _INITIAL_1|_XOR|A3|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|A3|RB _INITIAL_1|_XOR|A3|MID_SHUNT _INITIAL_1|_XOR|A3  2.050338398468e-12
B_INITIAL_1|_XOR|B1|1 _INITIAL_1|_XOR|B1 _INITIAL_1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|B1|P _INITIAL_1|_XOR|B1|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|B1|B _INITIAL_1|_XOR|B1 _INITIAL_1|_XOR|B1|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|B1|RB _INITIAL_1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_1|_XOR|B2|1 _INITIAL_1|_XOR|B2 _INITIAL_1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|B2|P _INITIAL_1|_XOR|B2|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|B2|B _INITIAL_1|_XOR|B2 _INITIAL_1|_XOR|B2|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|B2|RB _INITIAL_1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_1|_XOR|B3|1 _INITIAL_1|_XOR|B2 _INITIAL_1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|B3|P _INITIAL_1|_XOR|B3|MID_SERIES _INITIAL_1|_XOR|B3  1.2e-12
R_INITIAL_1|_XOR|B3|B _INITIAL_1|_XOR|B2 _INITIAL_1|_XOR|B3|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|B3|RB _INITIAL_1|_XOR|B3|MID_SHUNT _INITIAL_1|_XOR|B3  2.050338398468e-12
B_INITIAL_1|_XOR|T1|1 _INITIAL_1|_XOR|T1 _INITIAL_1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|T1|P _INITIAL_1|_XOR|T1|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|T1|B _INITIAL_1|_XOR|T1 _INITIAL_1|_XOR|T1|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|T1|RB _INITIAL_1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_1|_XOR|T2|1 _INITIAL_1|_XOR|T2 _INITIAL_1|_XOR|ABTQ JJMIT AREA=2.0
R_INITIAL_1|_XOR|T2|B _INITIAL_1|_XOR|T2 _INITIAL_1|_XOR|T2|MID_SHUNT  3.429952209
L_INITIAL_1|_XOR|T2|RB _INITIAL_1|_XOR|T2|MID_SHUNT _INITIAL_1|_XOR|ABTQ  2.437922998085e-12
B_INITIAL_1|_XOR|AB|1 _INITIAL_1|_XOR|AB _INITIAL_1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
L_INITIAL_1|_XOR|AB|P _INITIAL_1|_XOR|AB|MID_SERIES _INITIAL_1|_XOR|ABTQ  1.2e-12
R_INITIAL_1|_XOR|AB|B _INITIAL_1|_XOR|AB _INITIAL_1|_XOR|AB|MID_SHUNT  3.429952209
L_INITIAL_1|_XOR|AB|RB _INITIAL_1|_XOR|AB|MID_SHUNT _INITIAL_1|_XOR|ABTQ  2.437922998085e-12
B_INITIAL_1|_XOR|ABTQ|1 _INITIAL_1|_XOR|ABTQ _INITIAL_1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|ABTQ|P _INITIAL_1|_XOR|ABTQ|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|ABTQ|B _INITIAL_1|_XOR|ABTQ _INITIAL_1|_XOR|ABTQ|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|ABTQ|RB _INITIAL_1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_INITIAL_1|_XOR|Q1|1 _INITIAL_1|_XOR|Q1 _INITIAL_1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_XOR|Q1|P _INITIAL_1|_XOR|Q1|MID_SERIES 0  5e-13
R_INITIAL_1|_XOR|Q1|B _INITIAL_1|_XOR|Q1 _INITIAL_1|_XOR|Q1|MID_SHUNT  2.7439617672
L_INITIAL_1|_XOR|Q1|RB _INITIAL_1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
L_INITIAL_1|_AND|I_A1|B _INITIAL_1|_AND|A1 _INITIAL_1|_AND|I_A1|MID  2e-12
I_INITIAL_1|_AND|I_A1|B 0 _INITIAL_1|_AND|I_A1|MID  0.000175
L_INITIAL_1|_AND|I_B1|B _INITIAL_1|_AND|B1 _INITIAL_1|_AND|I_B1|MID  2e-12
I_INITIAL_1|_AND|I_B1|B 0 _INITIAL_1|_AND|I_B1|MID  0.000175
L_INITIAL_1|_AND|I_Q3|B _INITIAL_1|_AND|Q3 _INITIAL_1|_AND|I_Q3|MID  2e-12
I_INITIAL_1|_AND|I_Q3|B 0 _INITIAL_1|_AND|I_Q3|MID  5e-05
L_INITIAL_1|_AND|I_Q2|B _INITIAL_1|_AND|Q2 _INITIAL_1|_AND|I_Q2|MID  2e-12
I_INITIAL_1|_AND|I_Q2|B 0 _INITIAL_1|_AND|I_Q2|MID  0.000175
L_INITIAL_1|_AND|I_Q1|B _INITIAL_1|_AND|Q1 _INITIAL_1|_AND|I_Q1|MID  2e-12
I_INITIAL_1|_AND|I_Q1|B 0 _INITIAL_1|_AND|I_Q1|MID  0.000175
B_INITIAL_1|_AND|A1|1 _INITIAL_1|_AND|A1 _INITIAL_1|_AND|A1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_AND|A1|P _INITIAL_1|_AND|A1|MID_SERIES 0  2e-13
R_INITIAL_1|_AND|A1|B _INITIAL_1|_AND|A1 _INITIAL_1|_AND|A1|MID_SHUNT  2.7439617672
L_INITIAL_1|_AND|A1|RB _INITIAL_1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_AND|A2|1 _INITIAL_1|_AND|A2 _INITIAL_1|_AND|A2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_AND|A2|P _INITIAL_1|_AND|A2|MID_SERIES 0  2e-13
R_INITIAL_1|_AND|A2|B _INITIAL_1|_AND|A2 _INITIAL_1|_AND|A2|MID_SHUNT  2.7439617672
L_INITIAL_1|_AND|A2|RB _INITIAL_1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_AND|A12|1 _INITIAL_1|_AND|A2 _INITIAL_1|_AND|A3 JJMIT AREA=1.7857142857142858
R_INITIAL_1|_AND|A12|B _INITIAL_1|_AND|A2 _INITIAL_1|_AND|A12|MID_SHUNT  3.84154647408
L_INITIAL_1|_AND|A12|RB _INITIAL_1|_AND|A12|MID_SHUNT _INITIAL_1|_AND|A3  2.1704737578552e-12
B_INITIAL_1|_AND|B1|1 _INITIAL_1|_AND|B1 _INITIAL_1|_AND|B1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_AND|B1|P _INITIAL_1|_AND|B1|MID_SERIES 0  2e-13
R_INITIAL_1|_AND|B1|B _INITIAL_1|_AND|B1 _INITIAL_1|_AND|B1|MID_SHUNT  2.7439617672
L_INITIAL_1|_AND|B1|RB _INITIAL_1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_AND|B2|1 _INITIAL_1|_AND|B2 _INITIAL_1|_AND|B2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_AND|B2|P _INITIAL_1|_AND|B2|MID_SERIES 0  2e-13
R_INITIAL_1|_AND|B2|B _INITIAL_1|_AND|B2 _INITIAL_1|_AND|B2|MID_SHUNT  2.7439617672
L_INITIAL_1|_AND|B2|RB _INITIAL_1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_AND|B12|1 _INITIAL_1|_AND|B2 _INITIAL_1|_AND|B3 JJMIT AREA=1.7857142857142858
R_INITIAL_1|_AND|B12|B _INITIAL_1|_AND|B2 _INITIAL_1|_AND|B12|MID_SHUNT  3.84154647408
L_INITIAL_1|_AND|B12|RB _INITIAL_1|_AND|B12|MID_SHUNT _INITIAL_1|_AND|B3  2.1704737578552e-12
B_INITIAL_1|_AND|Q2|1 _INITIAL_1|_AND|Q2 _INITIAL_1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_AND|Q2|P _INITIAL_1|_AND|Q2|MID_SERIES 0  2e-13
R_INITIAL_1|_AND|Q2|B _INITIAL_1|_AND|Q2 _INITIAL_1|_AND|Q2|MID_SHUNT  2.7439617672
L_INITIAL_1|_AND|Q2|RB _INITIAL_1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
B_INITIAL_1|_AND|Q1|1 _INITIAL_1|_AND|Q1 _INITIAL_1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
L_INITIAL_1|_AND|Q1|P _INITIAL_1|_AND|Q1|MID_SERIES 0  2e-13
R_INITIAL_1|_AND|Q1|B _INITIAL_1|_AND|Q1 _INITIAL_1|_AND|Q1|MID_SHUNT  2.7439617672
L_INITIAL_1|_AND|Q1|RB _INITIAL_1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_SPL_G1|I_D1|B _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|I_D1|MID  2e-12
I_PG_01|_SPL_G1|I_D1|B 0 _PG_01|_SPL_G1|I_D1|MID  0.000175
L_PG_01|_SPL_G1|I_D2|B _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|I_D2|MID  2e-12
I_PG_01|_SPL_G1|I_D2|B 0 _PG_01|_SPL_G1|I_D2|MID  0.000245
L_PG_01|_SPL_G1|I_Q1|B _PG_01|_SPL_G1|QA1 _PG_01|_SPL_G1|I_Q1|MID  2e-12
I_PG_01|_SPL_G1|I_Q1|B 0 _PG_01|_SPL_G1|I_Q1|MID  0.000175
L_PG_01|_SPL_G1|I_Q2|B _PG_01|_SPL_G1|QB1 _PG_01|_SPL_G1|I_Q2|MID  2e-12
I_PG_01|_SPL_G1|I_Q2|B 0 _PG_01|_SPL_G1|I_Q2|MID  0.000175
B_PG_01|_SPL_G1|1|1 _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|1|P _PG_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|1|B _PG_01|_SPL_G1|D1 _PG_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|1|RB _PG_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_G1|2|1 _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|2|P _PG_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|2|B _PG_01|_SPL_G1|D2 _PG_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|2|RB _PG_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_G1|A|1 _PG_01|_SPL_G1|QA1 _PG_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|A|P _PG_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|A|B _PG_01|_SPL_G1|QA1 _PG_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|A|RB _PG_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_G1|B|1 _PG_01|_SPL_G1|QB1 _PG_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_G1|B|P _PG_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG_01|_SPL_G1|B|B _PG_01|_SPL_G1|QB1 _PG_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG_01|_SPL_G1|B|RB _PG_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_SPL_P1|I_D1|B _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|I_D1|MID  2e-12
I_PG_01|_SPL_P1|I_D1|B 0 _PG_01|_SPL_P1|I_D1|MID  0.000175
L_PG_01|_SPL_P1|I_D2|B _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|I_D2|MID  2e-12
I_PG_01|_SPL_P1|I_D2|B 0 _PG_01|_SPL_P1|I_D2|MID  0.000245
L_PG_01|_SPL_P1|I_Q1|B _PG_01|_SPL_P1|QA1 _PG_01|_SPL_P1|I_Q1|MID  2e-12
I_PG_01|_SPL_P1|I_Q1|B 0 _PG_01|_SPL_P1|I_Q1|MID  0.000175
L_PG_01|_SPL_P1|I_Q2|B _PG_01|_SPL_P1|QB1 _PG_01|_SPL_P1|I_Q2|MID  2e-12
I_PG_01|_SPL_P1|I_Q2|B 0 _PG_01|_SPL_P1|I_Q2|MID  0.000175
B_PG_01|_SPL_P1|1|1 _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|1|P _PG_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|1|B _PG_01|_SPL_P1|D1 _PG_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|1|RB _PG_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_P1|2|1 _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|2|P _PG_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|2|B _PG_01|_SPL_P1|D2 _PG_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|2|RB _PG_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_P1|A|1 _PG_01|_SPL_P1|QA1 _PG_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|A|P _PG_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|A|B _PG_01|_SPL_P1|QA1 _PG_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|A|RB _PG_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_SPL_P1|B|1 _PG_01|_SPL_P1|QB1 _PG_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG_01|_SPL_P1|B|P _PG_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG_01|_SPL_P1|B|B _PG_01|_SPL_P1|QB1 _PG_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG_01|_SPL_P1|B|RB _PG_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_PG|I_A1|B _PG_01|_PG|A1 _PG_01|_PG|I_A1|MID  2e-12
I_PG_01|_PG|I_A1|B 0 _PG_01|_PG|I_A1|MID  0.000175
L_PG_01|_PG|I_B1|B _PG_01|_PG|B1 _PG_01|_PG|I_B1|MID  2e-12
I_PG_01|_PG|I_B1|B 0 _PG_01|_PG|I_B1|MID  0.000175
L_PG_01|_PG|I_Q3|B _PG_01|_PG|Q3 _PG_01|_PG|I_Q3|MID  2e-12
I_PG_01|_PG|I_Q3|B 0 _PG_01|_PG|I_Q3|MID  0.00025
L_PG_01|_PG|I_Q2|B _PG_01|_PG|Q2 _PG_01|_PG|I_Q2|MID  2e-12
I_PG_01|_PG|I_Q2|B 0 _PG_01|_PG|I_Q2|MID  0.000175
L_PG_01|_PG|I_Q1|B _PG_01|_PG|Q1 _PG_01|_PG|I_Q1|MID  2e-12
I_PG_01|_PG|I_Q1|B 0 _PG_01|_PG|I_Q1|MID  0.000175
B_PG_01|_PG|A1|1 _PG_01|_PG|A1 _PG_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|A1|P _PG_01|_PG|A1|MID_SERIES 0  2e-13
R_PG_01|_PG|A1|B _PG_01|_PG|A1 _PG_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG_01|_PG|A1|RB _PG_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|A2|1 _PG_01|_PG|A2 _PG_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|A2|P _PG_01|_PG|A2|MID_SERIES 0  2e-13
R_PG_01|_PG|A2|B _PG_01|_PG|A2 _PG_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG_01|_PG|A2|RB _PG_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|A12|1 _PG_01|_PG|A2 _PG_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_PG|A12|B _PG_01|_PG|A2 _PG_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG_01|_PG|A12|RB _PG_01|_PG|A12|MID_SHUNT _PG_01|_PG|A3  2.1704737578552e-12
B_PG_01|_PG|B1|1 _PG_01|_PG|B1 _PG_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|B1|P _PG_01|_PG|B1|MID_SERIES 0  2e-13
R_PG_01|_PG|B1|B _PG_01|_PG|B1 _PG_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG_01|_PG|B1|RB _PG_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|B2|1 _PG_01|_PG|B2 _PG_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|B2|P _PG_01|_PG|B2|MID_SERIES 0  2e-13
R_PG_01|_PG|B2|B _PG_01|_PG|B2 _PG_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG_01|_PG|B2|RB _PG_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|B12|1 _PG_01|_PG|B2 _PG_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_PG|B12|B _PG_01|_PG|B2 _PG_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG_01|_PG|B12|RB _PG_01|_PG|B12|MID_SHUNT _PG_01|_PG|B3  2.1704737578552e-12
B_PG_01|_PG|Q2|1 _PG_01|_PG|Q2 _PG_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|Q2|P _PG_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG_01|_PG|Q2|B _PG_01|_PG|Q2 _PG_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG_01|_PG|Q2|RB _PG_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_PG|Q1|1 _PG_01|_PG|Q1 _PG_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_PG|Q1|P _PG_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG_01|_PG|Q1|B _PG_01|_PG|Q1 _PG_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG_01|_PG|Q1|RB _PG_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_GG|I_A1|B _PG_01|_GG|A1 _PG_01|_GG|I_A1|MID  2e-12
I_PG_01|_GG|I_A1|B 0 _PG_01|_GG|I_A1|MID  0.000175
L_PG_01|_GG|I_B1|B _PG_01|_GG|B1 _PG_01|_GG|I_B1|MID  2e-12
I_PG_01|_GG|I_B1|B 0 _PG_01|_GG|I_B1|MID  0.000175
L_PG_01|_GG|I_Q3|B _PG_01|_GG|Q3 _PG_01|_GG|I_Q3|MID  2e-12
I_PG_01|_GG|I_Q3|B 0 _PG_01|_GG|I_Q3|MID  0.00025
L_PG_01|_GG|I_Q2|B _PG_01|_GG|Q2 _PG_01|_GG|I_Q2|MID  2e-12
I_PG_01|_GG|I_Q2|B 0 _PG_01|_GG|I_Q2|MID  0.000175
L_PG_01|_GG|I_Q1|B _PG_01|_GG|Q1 _PG_01|_GG|I_Q1|MID  2e-12
I_PG_01|_GG|I_Q1|B 0 _PG_01|_GG|I_Q1|MID  0.000175
B_PG_01|_GG|A1|1 _PG_01|_GG|A1 _PG_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|A1|P _PG_01|_GG|A1|MID_SERIES 0  2e-13
R_PG_01|_GG|A1|B _PG_01|_GG|A1 _PG_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG_01|_GG|A1|RB _PG_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|A2|1 _PG_01|_GG|A2 _PG_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|A2|P _PG_01|_GG|A2|MID_SERIES 0  2e-13
R_PG_01|_GG|A2|B _PG_01|_GG|A2 _PG_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG_01|_GG|A2|RB _PG_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|A12|1 _PG_01|_GG|A2 _PG_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_GG|A12|B _PG_01|_GG|A2 _PG_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG_01|_GG|A12|RB _PG_01|_GG|A12|MID_SHUNT _PG_01|_GG|A3  2.1704737578552e-12
B_PG_01|_GG|B1|1 _PG_01|_GG|B1 _PG_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|B1|P _PG_01|_GG|B1|MID_SERIES 0  2e-13
R_PG_01|_GG|B1|B _PG_01|_GG|B1 _PG_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG_01|_GG|B1|RB _PG_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|B2|1 _PG_01|_GG|B2 _PG_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|B2|P _PG_01|_GG|B2|MID_SERIES 0  2e-13
R_PG_01|_GG|B2|B _PG_01|_GG|B2 _PG_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG_01|_GG|B2|RB _PG_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|B12|1 _PG_01|_GG|B2 _PG_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_GG|B12|B _PG_01|_GG|B2 _PG_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG_01|_GG|B12|RB _PG_01|_GG|B12|MID_SHUNT _PG_01|_GG|B3  2.1704737578552e-12
B_PG_01|_GG|Q2|1 _PG_01|_GG|Q2 _PG_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|Q2|P _PG_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG_01|_GG|Q2|B _PG_01|_GG|Q2 _PG_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG_01|_GG|Q2|RB _PG_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_GG|Q1|1 _PG_01|_GG|Q1 _PG_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_GG|Q1|P _PG_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG_01|_GG|Q1|B _PG_01|_GG|Q1 _PG_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG_01|_GG|Q1|RB _PG_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|1|1 _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|1|P _PG_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|1|B _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|1|RB _PG_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|23|1 _PG_01|_DFF_P0|2 _PG_01|_DFF_P0|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P0|23|B _PG_01|_DFF_P0|2 _PG_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P0|23|RB _PG_01|_DFF_P0|23|MID_SHUNT _PG_01|_DFF_P0|3  2.1704737578552e-12
B_PG_01|_DFF_P0|3|1 _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|3|P _PG_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|3|B _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|3|RB _PG_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|4|1 _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|4|P _PG_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|4|B _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|4|RB _PG_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|45|1 _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P0|45|B _PG_01|_DFF_P0|4 _PG_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P0|45|RB _PG_01|_DFF_P0|45|MID_SHUNT _PG_01|_DFF_P0|5  2.1704737578552e-12
B_PG_01|_DFF_P0|T|1 _PG_01|_DFF_P0|T1 _PG_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|T|P _PG_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|T|B _PG_01|_DFF_P0|T1 _PG_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|T|RB _PG_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P0|6|1 _PG_01|_DFF_P0|6 _PG_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P0|6|P _PG_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_P0|6|B _PG_01|_DFF_P0|6 _PG_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P0|6|RB _PG_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_P0|I_1|B _PG_01|_DFF_P0|1 _PG_01|_DFF_P0|I_1|MID  2e-12
I_PG_01|_DFF_P0|I_1|B 0 _PG_01|_DFF_P0|I_1|MID  0.000175
L_PG_01|_DFF_P0|I_3|B _PG_01|_DFF_P0|3 _PG_01|_DFF_P0|I_3|MID  2e-12
I_PG_01|_DFF_P0|I_3|B 0 _PG_01|_DFF_P0|I_3|MID  0.00025
L_PG_01|_DFF_P0|I_T|B _PG_01|_DFF_P0|T1 _PG_01|_DFF_P0|I_T|MID  2e-12
I_PG_01|_DFF_P0|I_T|B 0 _PG_01|_DFF_P0|I_T|MID  0.000175
L_PG_01|_DFF_P0|I_6|B _PG_01|_DFF_P0|6 _PG_01|_DFF_P0|I_6|MID  2e-12
I_PG_01|_DFF_P0|I_6|B 0 _PG_01|_DFF_P0|I_6|MID  0.000175
B_PG_01|_DFF_P1|1|1 _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|1|P _PG_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|1|B _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|1|RB _PG_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|23|1 _PG_01|_DFF_P1|2 _PG_01|_DFF_P1|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P1|23|B _PG_01|_DFF_P1|2 _PG_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P1|23|RB _PG_01|_DFF_P1|23|MID_SHUNT _PG_01|_DFF_P1|3  2.1704737578552e-12
B_PG_01|_DFF_P1|3|1 _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|3|P _PG_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|3|B _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|3|RB _PG_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|4|1 _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|4|P _PG_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|4|B _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|4|RB _PG_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|45|1 _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_P1|45|B _PG_01|_DFF_P1|4 _PG_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_P1|45|RB _PG_01|_DFF_P1|45|MID_SHUNT _PG_01|_DFF_P1|5  2.1704737578552e-12
B_PG_01|_DFF_P1|T|1 _PG_01|_DFF_P1|T1 _PG_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|T|P _PG_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|T|B _PG_01|_DFF_P1|T1 _PG_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|T|RB _PG_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_P1|6|1 _PG_01|_DFF_P1|6 _PG_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_P1|6|P _PG_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_P1|6|B _PG_01|_DFF_P1|6 _PG_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_P1|6|RB _PG_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_P1|I_1|B _PG_01|_DFF_P1|1 _PG_01|_DFF_P1|I_1|MID  2e-12
I_PG_01|_DFF_P1|I_1|B 0 _PG_01|_DFF_P1|I_1|MID  0.000175
L_PG_01|_DFF_P1|I_3|B _PG_01|_DFF_P1|3 _PG_01|_DFF_P1|I_3|MID  2e-12
I_PG_01|_DFF_P1|I_3|B 0 _PG_01|_DFF_P1|I_3|MID  0.00025
L_PG_01|_DFF_P1|I_T|B _PG_01|_DFF_P1|T1 _PG_01|_DFF_P1|I_T|MID  2e-12
I_PG_01|_DFF_P1|I_T|B 0 _PG_01|_DFF_P1|I_T|MID  0.000175
L_PG_01|_DFF_P1|I_6|B _PG_01|_DFF_P1|6 _PG_01|_DFF_P1|I_6|MID  2e-12
I_PG_01|_DFF_P1|I_6|B 0 _PG_01|_DFF_P1|I_6|MID  0.000175
B_PG_01|_DFF_PG|1|1 _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|1|P _PG_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|1|B _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|1|RB _PG_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|23|1 _PG_01|_DFF_PG|2 _PG_01|_DFF_PG|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_PG|23|B _PG_01|_DFF_PG|2 _PG_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_PG|23|RB _PG_01|_DFF_PG|23|MID_SHUNT _PG_01|_DFF_PG|3  2.1704737578552e-12
B_PG_01|_DFF_PG|3|1 _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|3|P _PG_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|3|B _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|3|RB _PG_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|4|1 _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|4|P _PG_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|4|B _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|4|RB _PG_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|45|1 _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_PG|45|B _PG_01|_DFF_PG|4 _PG_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_PG|45|RB _PG_01|_DFF_PG|45|MID_SHUNT _PG_01|_DFF_PG|5  2.1704737578552e-12
B_PG_01|_DFF_PG|T|1 _PG_01|_DFF_PG|T1 _PG_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|T|P _PG_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|T|B _PG_01|_DFF_PG|T1 _PG_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|T|RB _PG_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_PG|6|1 _PG_01|_DFF_PG|6 _PG_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_PG|6|P _PG_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_PG|6|B _PG_01|_DFF_PG|6 _PG_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_PG|6|RB _PG_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_PG|I_1|B _PG_01|_DFF_PG|1 _PG_01|_DFF_PG|I_1|MID  2e-12
I_PG_01|_DFF_PG|I_1|B 0 _PG_01|_DFF_PG|I_1|MID  0.000175
L_PG_01|_DFF_PG|I_3|B _PG_01|_DFF_PG|3 _PG_01|_DFF_PG|I_3|MID  2e-12
I_PG_01|_DFF_PG|I_3|B 0 _PG_01|_DFF_PG|I_3|MID  0.00025
L_PG_01|_DFF_PG|I_T|B _PG_01|_DFF_PG|T1 _PG_01|_DFF_PG|I_T|MID  2e-12
I_PG_01|_DFF_PG|I_T|B 0 _PG_01|_DFF_PG|I_T|MID  0.000175
L_PG_01|_DFF_PG|I_6|B _PG_01|_DFF_PG|6 _PG_01|_DFF_PG|I_6|MID  2e-12
I_PG_01|_DFF_PG|I_6|B 0 _PG_01|_DFF_PG|I_6|MID  0.000175
B_PG_01|_DFF_GG|1|1 _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|1|P _PG_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|1|B _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|1|RB _PG_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|23|1 _PG_01|_DFF_GG|2 _PG_01|_DFF_GG|3 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_GG|23|B _PG_01|_DFF_GG|2 _PG_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG_01|_DFF_GG|23|RB _PG_01|_DFF_GG|23|MID_SHUNT _PG_01|_DFF_GG|3  2.1704737578552e-12
B_PG_01|_DFF_GG|3|1 _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|3|P _PG_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|3|B _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|3|RB _PG_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|4|1 _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|4|P _PG_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|4|B _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|4|RB _PG_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|45|1 _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|5 JJMIT AREA=1.7857142857142858
R_PG_01|_DFF_GG|45|B _PG_01|_DFF_GG|4 _PG_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG_01|_DFF_GG|45|RB _PG_01|_DFF_GG|45|MID_SHUNT _PG_01|_DFF_GG|5  2.1704737578552e-12
B_PG_01|_DFF_GG|T|1 _PG_01|_DFF_GG|T1 _PG_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|T|P _PG_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|T|B _PG_01|_DFF_GG|T1 _PG_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|T|RB _PG_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_DFF_GG|6|1 _PG_01|_DFF_GG|6 _PG_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG_01|_DFF_GG|6|P _PG_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG_01|_DFF_GG|6|B _PG_01|_DFF_GG|6 _PG_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG_01|_DFF_GG|6|RB _PG_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_DFF_GG|I_1|B _PG_01|_DFF_GG|1 _PG_01|_DFF_GG|I_1|MID  2e-12
I_PG_01|_DFF_GG|I_1|B 0 _PG_01|_DFF_GG|I_1|MID  0.000175
L_PG_01|_DFF_GG|I_3|B _PG_01|_DFF_GG|3 _PG_01|_DFF_GG|I_3|MID  2e-12
I_PG_01|_DFF_GG|I_3|B 0 _PG_01|_DFF_GG|I_3|MID  0.00025
L_PG_01|_DFF_GG|I_T|B _PG_01|_DFF_GG|T1 _PG_01|_DFF_GG|I_T|MID  2e-12
I_PG_01|_DFF_GG|I_T|B 0 _PG_01|_DFF_GG|I_T|MID  0.000175
L_PG_01|_DFF_GG|I_6|B _PG_01|_DFF_GG|6 _PG_01|_DFF_GG|I_6|MID  2e-12
I_PG_01|_DFF_GG|I_6|B 0 _PG_01|_DFF_GG|I_6|MID  0.000175
L_PG_01|_AND_G|I_A1|B _PG_01|_AND_G|A1 _PG_01|_AND_G|I_A1|MID  2e-12
I_PG_01|_AND_G|I_A1|B 0 _PG_01|_AND_G|I_A1|MID  0.000175
L_PG_01|_AND_G|I_B1|B _PG_01|_AND_G|B1 _PG_01|_AND_G|I_B1|MID  2e-12
I_PG_01|_AND_G|I_B1|B 0 _PG_01|_AND_G|I_B1|MID  0.000175
L_PG_01|_AND_G|I_Q3|B _PG_01|_AND_G|Q3 _PG_01|_AND_G|I_Q3|MID  2e-12
I_PG_01|_AND_G|I_Q3|B 0 _PG_01|_AND_G|I_Q3|MID  5e-05
L_PG_01|_AND_G|I_Q2|B _PG_01|_AND_G|Q2 _PG_01|_AND_G|I_Q2|MID  2e-12
I_PG_01|_AND_G|I_Q2|B 0 _PG_01|_AND_G|I_Q2|MID  0.000175
L_PG_01|_AND_G|I_Q1|B _PG_01|_AND_G|Q1 _PG_01|_AND_G|I_Q1|MID  2e-12
I_PG_01|_AND_G|I_Q1|B 0 _PG_01|_AND_G|I_Q1|MID  0.000175
B_PG_01|_AND_G|A1|1 _PG_01|_AND_G|A1 _PG_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|A1|P _PG_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG_01|_AND_G|A1|B _PG_01|_AND_G|A1 _PG_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|A1|RB _PG_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|A2|1 _PG_01|_AND_G|A2 _PG_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|A2|P _PG_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG_01|_AND_G|A2|B _PG_01|_AND_G|A2 _PG_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|A2|RB _PG_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|A12|1 _PG_01|_AND_G|A2 _PG_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_G|A12|B _PG_01|_AND_G|A2 _PG_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG_01|_AND_G|A12|RB _PG_01|_AND_G|A12|MID_SHUNT _PG_01|_AND_G|A3  2.1704737578552e-12
B_PG_01|_AND_G|B1|1 _PG_01|_AND_G|B1 _PG_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|B1|P _PG_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG_01|_AND_G|B1|B _PG_01|_AND_G|B1 _PG_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|B1|RB _PG_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|B2|1 _PG_01|_AND_G|B2 _PG_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|B2|P _PG_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG_01|_AND_G|B2|B _PG_01|_AND_G|B2 _PG_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|B2|RB _PG_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|B12|1 _PG_01|_AND_G|B2 _PG_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_G|B12|B _PG_01|_AND_G|B2 _PG_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG_01|_AND_G|B12|RB _PG_01|_AND_G|B12|MID_SHUNT _PG_01|_AND_G|B3  2.1704737578552e-12
B_PG_01|_AND_G|Q2|1 _PG_01|_AND_G|Q2 _PG_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|Q2|P _PG_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG_01|_AND_G|Q2|B _PG_01|_AND_G|Q2 _PG_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|Q2|RB _PG_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_G|Q1|1 _PG_01|_AND_G|Q1 _PG_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_G|Q1|P _PG_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG_01|_AND_G|Q1|B _PG_01|_AND_G|Q1 _PG_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG_01|_AND_G|Q1|RB _PG_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG_01|_AND_P|I_A1|B _PG_01|_AND_P|A1 _PG_01|_AND_P|I_A1|MID  2e-12
I_PG_01|_AND_P|I_A1|B 0 _PG_01|_AND_P|I_A1|MID  0.000175
L_PG_01|_AND_P|I_B1|B _PG_01|_AND_P|B1 _PG_01|_AND_P|I_B1|MID  2e-12
I_PG_01|_AND_P|I_B1|B 0 _PG_01|_AND_P|I_B1|MID  0.000175
L_PG_01|_AND_P|I_Q3|B _PG_01|_AND_P|Q3 _PG_01|_AND_P|I_Q3|MID  2e-12
I_PG_01|_AND_P|I_Q3|B 0 _PG_01|_AND_P|I_Q3|MID  5e-05
L_PG_01|_AND_P|I_Q2|B _PG_01|_AND_P|Q2 _PG_01|_AND_P|I_Q2|MID  2e-12
I_PG_01|_AND_P|I_Q2|B 0 _PG_01|_AND_P|I_Q2|MID  0.000175
L_PG_01|_AND_P|I_Q1|B _PG_01|_AND_P|Q1 _PG_01|_AND_P|I_Q1|MID  2e-12
I_PG_01|_AND_P|I_Q1|B 0 _PG_01|_AND_P|I_Q1|MID  0.000175
B_PG_01|_AND_P|A1|1 _PG_01|_AND_P|A1 _PG_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|A1|P _PG_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG_01|_AND_P|A1|B _PG_01|_AND_P|A1 _PG_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|A1|RB _PG_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|A2|1 _PG_01|_AND_P|A2 _PG_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|A2|P _PG_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG_01|_AND_P|A2|B _PG_01|_AND_P|A2 _PG_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|A2|RB _PG_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|A12|1 _PG_01|_AND_P|A2 _PG_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_P|A12|B _PG_01|_AND_P|A2 _PG_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG_01|_AND_P|A12|RB _PG_01|_AND_P|A12|MID_SHUNT _PG_01|_AND_P|A3  2.1704737578552e-12
B_PG_01|_AND_P|B1|1 _PG_01|_AND_P|B1 _PG_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|B1|P _PG_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG_01|_AND_P|B1|B _PG_01|_AND_P|B1 _PG_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|B1|RB _PG_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|B2|1 _PG_01|_AND_P|B2 _PG_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|B2|P _PG_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG_01|_AND_P|B2|B _PG_01|_AND_P|B2 _PG_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|B2|RB _PG_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|B12|1 _PG_01|_AND_P|B2 _PG_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG_01|_AND_P|B12|B _PG_01|_AND_P|B2 _PG_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG_01|_AND_P|B12|RB _PG_01|_AND_P|B12|MID_SHUNT _PG_01|_AND_P|B3  2.1704737578552e-12
B_PG_01|_AND_P|Q2|1 _PG_01|_AND_P|Q2 _PG_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|Q2|P _PG_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG_01|_AND_P|Q2|B _PG_01|_AND_P|Q2 _PG_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|Q2|RB _PG_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG_01|_AND_P|Q1|1 _PG_01|_AND_P|Q1 _PG_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG_01|_AND_P|Q1|P _PG_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG_01|_AND_P|Q1|B _PG_01|_AND_P|Q1 _PG_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG_01|_AND_P|Q1|RB _PG_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI RS0
.print DEVI RS1
.print DEVI RIG1
.print DEVI RS2
.print DEVI RP1
.print DEVI RG1
.print DEVI IDATA_A0|A
.print DEVI IDATA_B0|B
.print DEVI IDATA_A1|C
.print DEVI IDATA_B1|D
.print DEVI IT1|T
.print DEVI IT2|T
.print DEVI L_SPL_P0|1
.print DEVI L_SPL_P0|2
.print DEVI L_SPL_P0|3
.print DEVI L_SPL_P0|4
.print DEVI L_SPL_P0|5
.print DEVI L_SPL_P0|6
.print DEVI L_SPL_P0|7
.print DEVI L_SPL_G0|1
.print DEVI L_SPL_G0|2
.print DEVI L_SPL_G0|3
.print DEVI L_SPL_G0|4
.print DEVI L_SPL_G0|5
.print DEVI L_SPL_G0|6
.print DEVI L_SPL_G0|7
.print DEVI L_SPL_P1|1
.print DEVI L_SPL_P1|2
.print DEVI L_SPL_P1|3
.print DEVI L_SPL_P1|4
.print DEVI L_SPL_P1|5
.print DEVI L_SPL_P1|6
.print DEVI L_SPL_P1|7
.print DEVI L_SPL_G1|1
.print DEVI L_SPL_G1|2
.print DEVI L_SPL_G1|3
.print DEVI L_SPL_G1|4
.print DEVI L_SPL_G1|5
.print DEVI L_SPL_G1|6
.print DEVI L_SPL_G1|7
.print DEVI IT3|T
.print DEVI IT4|T
.print DEVI L_DFF_IP0_01|1
.print DEVI L_DFF_IP0_01|2
.print DEVI L_DFF_IP0_01|3
.print DEVI L_DFF_IP0_01|4
.print DEVI L_DFF_IP0_01|T
.print DEVI L_DFF_IP0_01|5
.print DEVI L_DFF_IP0_01|6
.print DEVI IT5|T
.print DEVI L_DFF_IP0_12|1
.print DEVI L_DFF_IP0_12|2
.print DEVI L_DFF_IP0_12|3
.print DEVI L_DFF_IP0_12|4
.print DEVI L_DFF_IP0_12|T
.print DEVI L_DFF_IP0_12|5
.print DEVI L_DFF_IP0_12|6
.print DEVI IT6|T
.print DEVI L_DFF_IG0_01|1
.print DEVI L_DFF_IG0_01|2
.print DEVI L_DFF_IG0_01|3
.print DEVI L_DFF_IG0_01|4
.print DEVI L_DFF_IG0_01|T
.print DEVI L_DFF_IG0_01|5
.print DEVI L_DFF_IG0_01|6
.print DEVI IT7|T
.print DEVI L_DFF_IP1_01|1
.print DEVI L_DFF_IP1_01|2
.print DEVI L_DFF_IP1_01|3
.print DEVI L_DFF_IP1_01|4
.print DEVI L_DFF_IP1_01|T
.print DEVI L_DFF_IP1_01|5
.print DEVI L_DFF_IP1_01|6
.print DEVI IT8|T
.print DEVI L_XOR_S1|A1
.print DEVI L_XOR_S1|A2
.print DEVI L_XOR_S1|A3
.print DEVI L_XOR_S1|B1
.print DEVI L_XOR_S1|B2
.print DEVI L_XOR_S1|B3
.print DEVI L_XOR_S1|T1
.print DEVI L_XOR_S1|T2
.print DEVI L_XOR_S1|Q2
.print DEVI L_XOR_S1|Q1
.print DEVI IT9|T
.print DEVI L_DFF_IG1_01|1
.print DEVI L_DFF_IG1_01|2
.print DEVI L_DFF_IG1_01|3
.print DEVI L_DFF_IG1_01|4
.print DEVI L_DFF_IG1_01|T
.print DEVI L_DFF_IG1_01|5
.print DEVI L_DFF_IG1_01|6
.print DEVI IT10|T
.print DEVI L_DFF_S2|1
.print DEVI L_DFF_S2|2
.print DEVI L_DFF_S2|3
.print DEVI L_DFF_S2|4
.print DEVI L_DFF_S2|T
.print DEVI L_DFF_S2|5
.print DEVI L_DFF_S2|6
.print V _PG_01|GG
.print V _SPL_P1|QB1
.print V _SPL_P1|D1
.print V _DFF_IG0_01|T1
.print V _DFF_IP0_12|6
.print V _DFF_IP0_01|5
.print V IP1_0
.print V _DFF_IP1_01|3
.print V _XOR_S1|A2
.print V _INITIAL_1|B1_SYNC
.print V IP0_0_B
.print V _DFF_IP1_01|5
.print V _PG_01|P1_SYNC
.print V _PG_01|G1_COPY_2
.print V IG1_1
.print V P1_1
.print V CLK5
.print V _PG_01|P0_SYNC
.print V _SPL_G0|D1
.print V _XOR_S1|A3
.print V _SPL_G1|D2
.print V A0
.print V _SPL_P0|D1
.print V _DFF_IP0_01|2
.print V _DFF_IP1_01|1
.print V _DFF_S2|T1
.print V _DFF_IP0_01|6
.print V CLK1
.print V _XOR_S1|B2
.print V _XOR_S1|T2
.print V _PG_01|PG
.print V _DFF_IP0_01|4
.print V IP0_1
.print V _DFF_S2|2
.print V _SPL_G0|QA1
.print V _PG_01|G1_COPY_1
.print V _DFF_S2|6
.print V _DFF_S2|1
.print V CLK2
.print V B0
.print V _DFF_S2|3
.print V _INITIAL_1|A1_SYNC
.print V _DFF_IG1_01|2
.print V IG0_0_W
.print V G1_1
.print V _SPL_P1|JCT
.print V _DFF_S2|4
.print V _DFF_IP0_12|T1
.print V CLK9
.print V _SPL_G0|JCT
.print V _SPL_P0|QB1
.print V _DFF_IP0_12|1
.print V _INITIAL_0|B1_SYNC
.print V _DFF_S2|5
.print V _DFF_IP0_12|5
.print V IP0_0_W
.print V _INITIAL_1|A1
.print V _DFF_IP0_12|4
.print V _DFF_IG0_01|4
.print V _INITIAL_0|A1_SYNC
.print V _SPL_G1|QA1
.print V _PG_01|P1_COPY_2
.print V _DFF_IG0_01|3
.print V _DFF_IP0_01|3
.print V _XOR_S1|B1
.print V _SPL_G0|QB1
.print V CLK3
.print V _XOR_S1|Q1
.print V B1
.print V _XOR_S1|AB
.print V _DFF_IG1_01|6
.print V A1
.print V _XOR_S1|T1
.print V _SPL_G1|JCT
.print V _INITIAL_0|A2
.print V _DFF_IP1_01|6
.print V _XOR_S1|B3
.print V _SPL_P0|JCT
.print V _DFF_IP0_12|2
.print V _INITIAL_0|B2
.print V IP0_0
.print V _DFF_IP0_01|1
.print V S2
.print V _SPL_P0|D2
.print V IG1_0_W
.print V IG1_0_B
.print V IP1_0_B
.print V _INITIAL_0|B1
.print V _DFF_IG0_01|2
.print V _SPL_P0|QA1
.print V CLK8
.print V _DFF_IG1_01|5
.print V _SPL_G1|QB1
.print V _PG_01|GG_SYNC
.print V CLK7
.print V _DFF_IG1_01|4
.print V _DFF_IP0_12|3
.print V IG0_1
.print V _DFF_IG1_01|1
.print V IG0_0_B
.print V _XOR_S1|ABTQ
.print V _SPL_P1|D2
.print V _PG_01|P1_COPY_1
.print V IG0_0
.print V _DFF_IG0_01|5
.print V _DFF_IP1_01|T1
.print V _SPL_G0|D2
.print V CLK4
.print V S0
.print V S1
.print V IP1_1
.print V _DFF_IG1_01|T1
.print V _PG_01|PG_SYNC
.print V _DFF_IG0_01|1
.print V CLK10
.print V CLK6
.print V _DFF_IG1_01|3
.print V IG1_0
.print V _SPL_P1|QA1
.print V _DFF_IP0_01|T1
.print V _INITIAL_1|B2
.print V _INITIAL_0|A1
.print V _INITIAL_1|B1
.print V IP1_0_W
.print V _SPL_G1|D1
.print V _INITIAL_1|A2
.print V _DFF_IP1_01|4
.print V _XOR_S1|A1
.print V _DFF_IP1_01|2
.print V _DFF_IG0_01|6
