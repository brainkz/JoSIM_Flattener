*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=0
.PARAM TCLOCK=1e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.1E-12 0.45E-09
ROUT Q 0  1
IT1|T 0 CLK  PWL(0 0 -3e-12 0 0 0.0005 3e-12 0 9.7e-11 0 1e-10 0.0005 1.03e-10 0 1.97e-10 0 2e-10 0.0005 2.03e-10 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 3.97e-10 0 4e-10 0.0005 4.03e-10 0 4.97e-10 0 5e-10 0.0005 5.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 6.97e-10 0 7e-10 0.0005 7.03e-10 0 7.97e-10 0 8e-10 0.0005 8.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 9.97e-10 0 1e-09 0.0005 1.003e-09 0 1.097e-09 0 1.1e-09 0.0005 1.103e-09 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.297e-09 0 1.3e-09 0.0005 1.303e-09 0 1.397e-09 0 1.4e-09 0.0005 1.403e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.597e-09 0 1.6e-09 0.0005 1.603e-09 0 1.697e-09 0 1.7e-09 0.0005 1.703e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 1.897e-09 0 1.9e-09 0.0005 1.903e-09 0 1.997e-09 0 2e-09 0.0005 2.003e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.197e-09 0 2.2e-09 0.0005 2.203e-09 0 2.297e-09 0 2.3e-09 0.0005 2.303e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.497e-09 0 2.5e-09 0.0005 2.503e-09 0 2.597e-09 0 2.6e-09 0.0005 2.603e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.797e-09 0 2.8e-09 0.0005 2.803e-09 0 2.897e-09 0 2.9e-09 0.0005 2.903e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.097e-09 0 3.1e-09 0.0005 3.103e-09 0 3.197e-09 0 3.2e-09 0.0005 3.203e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.397e-09 0 3.4e-09 0.0005 3.403e-09 0 3.497e-09 0 3.5e-09 0.0005 3.503e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.697e-09 0 3.7e-09 0.0005 3.703e-09 0 3.797e-09 0 3.8e-09 0.0005 3.803e-09 0)
IDATA_A1|A 0 A  PWL(0 0 1.07e-10 0 1.1e-10 0.0005 1.13e-10 0 3.07e-10 0 3.1e-10 0.0005 3.13e-10 0 5.07e-10 0 5.1e-10 0.0005 5.13e-10 0 7.07e-10 0 7.1e-10 0.0005 7.13e-10 0 9.07e-10 0 9.1e-10 0.0005 9.13e-10 0 1.107e-09 0 1.11e-09 0.0005 1.113e-09 0 1.307e-09 0 1.31e-09 0.0005 1.313e-09 0 1.507e-09 0 1.51e-09 0.0005 1.513e-09 0 1.707e-09 0 1.71e-09 0.0005 1.713e-09 0 1.907e-09 0 1.91e-09 0.0005 1.913e-09 0 2.107e-09 0 2.11e-09 0.0005 2.113e-09 0 2.307e-09 0 2.31e-09 0.0005 2.313e-09 0 2.507e-09 0 2.51e-09 0.0005 2.513e-09 0 2.707e-09 0 2.71e-09 0.0005 2.713e-09 0 2.907e-09 0 2.91e-09 0.0005 2.913e-09 0 3.107e-09 0 3.11e-09 0.0005 3.113e-09 0 3.307e-09 0 3.31e-09 0.0005 3.313e-09 0 3.507e-09 0 3.51e-09 0.0005 3.513e-09 0 3.707e-09 0 3.71e-09 0.0005 3.713e-09 0)
IDATA_B1|B 0 B  PWL(0 0 2.67e-10 0 2.7e-10 0.0005 2.73e-10 0 3.67e-10 0 3.7e-10 0.0005 3.73e-10 0 6.67e-10 0 6.7e-10 0.0005 6.73e-10 0 7.67e-10 0 7.7e-10 0.0005 7.73e-10 0 1.067e-09 0 1.07e-09 0.0005 1.073e-09 0 1.167e-09 0 1.17e-09 0.0005 1.173e-09 0 1.467e-09 0 1.47e-09 0.0005 1.473e-09 0 1.567e-09 0 1.57e-09 0.0005 1.573e-09 0 1.867e-09 0 1.87e-09 0.0005 1.873e-09 0 1.967e-09 0 1.97e-09 0.0005 1.973e-09 0 2.267e-09 0 2.27e-09 0.0005 2.273e-09 0 2.367e-09 0 2.37e-09 0.0005 2.373e-09 0 2.667e-09 0 2.67e-09 0.0005 2.673e-09 0 2.767e-09 0 2.77e-09 0.0005 2.773e-09 0 3.067e-09 0 3.07e-09 0.0005 3.073e-09 0 3.167e-09 0 3.17e-09 0.0005 3.173e-09 0 3.467e-09 0 3.47e-09 0.0005 3.473e-09 0 3.567e-09 0 3.57e-09 0.0005 3.573e-09 0 3.867e-09 0 3.87e-09 0.0005 3.873e-09 0)
IDATA_C1|C 0 C  PWL(0 0 3.7e-11 0 4e-11 0.0005 4.3e-11 0 1.37e-10 0 1.4e-10 0.0005 1.43e-10 0 2.37e-10 0 2.4e-10 0.0005 2.43e-10 0 3.37e-10 0 3.4e-10 0.0005 3.43e-10 0 8.37e-10 0 8.4e-10 0.0005 8.43e-10 0 9.37e-10 0 9.4e-10 0.0005 9.43e-10 0 1.037e-09 0 1.04e-09 0.0005 1.043e-09 0 1.137e-09 0 1.14e-09 0.0005 1.143e-09 0 1.637e-09 0 1.64e-09 0.0005 1.643e-09 0 1.737e-09 0 1.74e-09 0.0005 1.743e-09 0 1.837e-09 0 1.84e-09 0.0005 1.843e-09 0 1.937e-09 0 1.94e-09 0.0005 1.943e-09 0 2.437e-09 0 2.44e-09 0.0005 2.443e-09 0 2.537e-09 0 2.54e-09 0.0005 2.543e-09 0 2.637e-09 0 2.64e-09 0.0005 2.643e-09 0 2.737e-09 0 2.74e-09 0.0005 2.743e-09 0 3.237e-09 0 3.24e-09 0.0005 3.243e-09 0 3.337e-09 0 3.34e-09 0.0005 3.343e-09 0 3.437e-09 0 3.44e-09 0.0005 3.443e-09 0 3.537e-09 0 3.54e-09 0.0005 3.543e-09 0)
L_MERGE|A1 A _MERGE|A1  2.067833848e-12
L_MERGE|A2 _MERGE|A1 _MERGE|A2  4.135667696e-12
L_MERGE|A3 _MERGE|A3 _MERGE|Q3  1.2e-12
L_MERGE|B1 B _MERGE|B1  2.067833848e-12
L_MERGE|B2 _MERGE|B1 _MERGE|B2  4.135667696e-12
L_MERGE|B3 _MERGE|B3 _MERGE|Q3  1.2e-12
L_MERGE|Q3 _MERGE|Q3 _MERGE|Q2  4.135667696e-12
L_MERGE|Q2 _MERGE|Q2 _MERGE|Q1  4.135667696e-12
L_MERGE|Q1 _MERGE|Q1 A_OR_B  2.067833848e-12
L_XOR|A1 A_OR_B _XOR|A1  2.067833848e-12
L_XOR|A2 _XOR|A1 _XOR|A2  4.135667696e-12
L_XOR|A3 _XOR|A3 _XOR|AB  8.271335392e-12
L_XOR|B1 C _XOR|B1  2.067833848e-12
L_XOR|B2 _XOR|B1 _XOR|B2  4.135667696e-12
L_XOR|B3 _XOR|B3 _XOR|AB  8.271335392e-12
L_XOR|T1 CLK _XOR|T1  2.067833848e-12
L_XOR|T2 _XOR|T1 _XOR|T2  4.135667696e-12
L_XOR|Q2 _XOR|ABTQ _XOR|Q1  4.135667696e-12
L_XOR|Q1 _XOR|Q1 Q  2.067833848e-12
L_MERGE|I_A1|B _MERGE|A1 _MERGE|I_A1|MID  2e-12
I_MERGE|I_A1|B 0 _MERGE|I_A1|MID  0.000175
L_MERGE|I_B1|B _MERGE|B1 _MERGE|I_B1|MID  2e-12
I_MERGE|I_B1|B 0 _MERGE|I_B1|MID  0.000175
L_MERGE|I_Q3|B _MERGE|Q3 _MERGE|I_Q3|MID  2e-12
I_MERGE|I_Q3|B 0 _MERGE|I_Q3|MID  0.00025
L_MERGE|I_Q2|B _MERGE|Q2 _MERGE|I_Q2|MID  2e-12
I_MERGE|I_Q2|B 0 _MERGE|I_Q2|MID  0.000175
L_MERGE|I_Q1|B _MERGE|Q1 _MERGE|I_Q1|MID  2e-12
I_MERGE|I_Q1|B 0 _MERGE|I_Q1|MID  0.000175
B_MERGE|A1|1 _MERGE|A1 _MERGE|A1|MID_SERIES JJMIT AREA=2.5
L_MERGE|A1|P _MERGE|A1|MID_SERIES 0  2e-13
R_MERGE|A1|B _MERGE|A1 _MERGE|A1|MID_SHUNT  2.7439617672
L_MERGE|A1|RB _MERGE|A1|MID_SHUNT 0  1.550338398468e-12
B_MERGE|A2|1 _MERGE|A2 _MERGE|A2|MID_SERIES JJMIT AREA=2.5
L_MERGE|A2|P _MERGE|A2|MID_SERIES 0  2e-13
R_MERGE|A2|B _MERGE|A2 _MERGE|A2|MID_SHUNT  2.7439617672
L_MERGE|A2|RB _MERGE|A2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|A12|1 _MERGE|A2 _MERGE|A3 JJMIT AREA=1.7857142857142858
R_MERGE|A12|B _MERGE|A2 _MERGE|A12|MID_SHUNT  3.84154647408
L_MERGE|A12|RB _MERGE|A12|MID_SHUNT _MERGE|A3  2.1704737578552e-12
B_MERGE|B1|1 _MERGE|B1 _MERGE|B1|MID_SERIES JJMIT AREA=2.5
L_MERGE|B1|P _MERGE|B1|MID_SERIES 0  2e-13
R_MERGE|B1|B _MERGE|B1 _MERGE|B1|MID_SHUNT  2.7439617672
L_MERGE|B1|RB _MERGE|B1|MID_SHUNT 0  1.550338398468e-12
B_MERGE|B2|1 _MERGE|B2 _MERGE|B2|MID_SERIES JJMIT AREA=2.5
L_MERGE|B2|P _MERGE|B2|MID_SERIES 0  2e-13
R_MERGE|B2|B _MERGE|B2 _MERGE|B2|MID_SHUNT  2.7439617672
L_MERGE|B2|RB _MERGE|B2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|B12|1 _MERGE|B2 _MERGE|B3 JJMIT AREA=1.7857142857142858
R_MERGE|B12|B _MERGE|B2 _MERGE|B12|MID_SHUNT  3.84154647408
L_MERGE|B12|RB _MERGE|B12|MID_SHUNT _MERGE|B3  2.1704737578552e-12
B_MERGE|Q2|1 _MERGE|Q2 _MERGE|Q2|MID_SERIES JJMIT AREA=2.5
L_MERGE|Q2|P _MERGE|Q2|MID_SERIES 0  2e-13
R_MERGE|Q2|B _MERGE|Q2 _MERGE|Q2|MID_SHUNT  2.7439617672
L_MERGE|Q2|RB _MERGE|Q2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|Q1|1 _MERGE|Q1 _MERGE|Q1|MID_SERIES JJMIT AREA=2.5
L_MERGE|Q1|P _MERGE|Q1|MID_SERIES 0  2e-13
R_MERGE|Q1|B _MERGE|Q1 _MERGE|Q1|MID_SHUNT  2.7439617672
L_MERGE|Q1|RB _MERGE|Q1|MID_SHUNT 0  1.550338398468e-12
L_XOR|I_A1|B _XOR|A1 _XOR|I_A1|MID  2e-12
I_XOR|I_A1|B 0 _XOR|I_A1|MID  0.000175
L_XOR|I_A3|B _XOR|A3 _XOR|I_A3|MID  2e-12
I_XOR|I_A3|B 0 _XOR|I_A3|MID  0.000175
L_XOR|I_B1|B _XOR|B1 _XOR|I_B1|MID  2e-12
I_XOR|I_B1|B 0 _XOR|I_B1|MID  0.000175
L_XOR|I_B3|B _XOR|B3 _XOR|I_B3|MID  2e-12
I_XOR|I_B3|B 0 _XOR|I_B3|MID  0.000175
L_XOR|I_T1|B _XOR|T1 _XOR|I_T1|MID  2e-12
I_XOR|I_T1|B 0 _XOR|I_T1|MID  0.000175
L_XOR|I_Q1|B _XOR|Q1 _XOR|I_Q1|MID  2e-12
I_XOR|I_Q1|B 0 _XOR|I_Q1|MID  0.000175
B_XOR|A1|1 _XOR|A1 _XOR|A1|MID_SERIES JJMIT AREA=2.5
L_XOR|A1|P _XOR|A1|MID_SERIES 0  5e-13
R_XOR|A1|B _XOR|A1 _XOR|A1|MID_SHUNT  2.7439617672
L_XOR|A1|RB _XOR|A1|MID_SHUNT 0  2.050338398468e-12
B_XOR|A2|1 _XOR|A2 _XOR|A2|MID_SERIES JJMIT AREA=2.5
L_XOR|A2|P _XOR|A2|MID_SERIES 0  5e-13
R_XOR|A2|B _XOR|A2 _XOR|A2|MID_SHUNT  2.7439617672
L_XOR|A2|RB _XOR|A2|MID_SHUNT 0  2.050338398468e-12
B_XOR|A3|1 _XOR|A2 _XOR|A3|MID_SERIES JJMIT AREA=2.5
L_XOR|A3|P _XOR|A3|MID_SERIES _XOR|A3  1.2e-12
R_XOR|A3|B _XOR|A2 _XOR|A3|MID_SHUNT  2.7439617672
L_XOR|A3|RB _XOR|A3|MID_SHUNT _XOR|A3  2.050338398468e-12
B_XOR|B1|1 _XOR|B1 _XOR|B1|MID_SERIES JJMIT AREA=2.5
L_XOR|B1|P _XOR|B1|MID_SERIES 0  5e-13
R_XOR|B1|B _XOR|B1 _XOR|B1|MID_SHUNT  2.7439617672
L_XOR|B1|RB _XOR|B1|MID_SHUNT 0  2.050338398468e-12
B_XOR|B2|1 _XOR|B2 _XOR|B2|MID_SERIES JJMIT AREA=2.5
L_XOR|B2|P _XOR|B2|MID_SERIES 0  5e-13
R_XOR|B2|B _XOR|B2 _XOR|B2|MID_SHUNT  2.7439617672
L_XOR|B2|RB _XOR|B2|MID_SHUNT 0  2.050338398468e-12
B_XOR|B3|1 _XOR|B2 _XOR|B3|MID_SERIES JJMIT AREA=2.5
L_XOR|B3|P _XOR|B3|MID_SERIES _XOR|B3  1.2e-12
R_XOR|B3|B _XOR|B2 _XOR|B3|MID_SHUNT  2.7439617672
L_XOR|B3|RB _XOR|B3|MID_SHUNT _XOR|B3  2.050338398468e-12
B_XOR|T1|1 _XOR|T1 _XOR|T1|MID_SERIES JJMIT AREA=2.5
L_XOR|T1|P _XOR|T1|MID_SERIES 0  5e-13
R_XOR|T1|B _XOR|T1 _XOR|T1|MID_SHUNT  2.7439617672
L_XOR|T1|RB _XOR|T1|MID_SHUNT 0  2.050338398468e-12
B_XOR|T2|1 _XOR|T2 _XOR|ABTQ JJMIT AREA=2.0
R_XOR|T2|B _XOR|T2 _XOR|T2|MID_SHUNT  3.429952209
L_XOR|T2|RB _XOR|T2|MID_SHUNT _XOR|ABTQ  2.437922998085e-12
B_XOR|AB|1 _XOR|AB _XOR|AB|MID_SERIES JJMIT AREA=2.0
L_XOR|AB|P _XOR|AB|MID_SERIES _XOR|ABTQ  1.2e-12
R_XOR|AB|B _XOR|AB _XOR|AB|MID_SHUNT  3.429952209
L_XOR|AB|RB _XOR|AB|MID_SHUNT _XOR|ABTQ  2.437922998085e-12
B_XOR|ABTQ|1 _XOR|ABTQ _XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
L_XOR|ABTQ|P _XOR|ABTQ|MID_SERIES 0  5e-13
R_XOR|ABTQ|B _XOR|ABTQ _XOR|ABTQ|MID_SHUNT  2.7439617672
L_XOR|ABTQ|RB _XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
B_XOR|Q1|1 _XOR|Q1 _XOR|Q1|MID_SERIES JJMIT AREA=2.5
L_XOR|Q1|P _XOR|Q1|MID_SERIES 0  5e-13
R_XOR|Q1|B _XOR|Q1 _XOR|Q1|MID_SHUNT  2.7439617672
L_XOR|Q1|RB _XOR|Q1|MID_SHUNT 0  2.050338398468e-12
.print DEVI ROUT
.print DEVI IT1|T
.print DEVI IDATA_A1|A
.print DEVI IDATA_B1|B
.print DEVI IDATA_C1|C
.print DEVI L_MERGE|A1
.print DEVI L_MERGE|A2
.print DEVI L_MERGE|A3
.print DEVI L_MERGE|B1
.print DEVI L_MERGE|B2
.print DEVI L_MERGE|B3
.print DEVI L_MERGE|Q3
.print DEVI L_MERGE|Q2
.print DEVI L_MERGE|Q1
.print DEVI L_XOR|A1
.print DEVI L_XOR|A2
.print DEVI L_XOR|A3
.print DEVI L_XOR|B1
.print DEVI L_XOR|B2
.print DEVI L_XOR|B3
.print DEVI L_XOR|T1
.print DEVI L_XOR|T2
.print DEVI L_XOR|Q2
.print DEVI L_XOR|Q1
.print DEVI L_MERGE|I_A1|B
.print DEVI I_MERGE|I_A1|B
.print DEVI L_MERGE|I_B1|B
.print DEVI I_MERGE|I_B1|B
.print DEVI L_MERGE|I_Q3|B
.print DEVI I_MERGE|I_Q3|B
.print DEVI L_MERGE|I_Q2|B
.print DEVI I_MERGE|I_Q2|B
.print DEVI L_MERGE|I_Q1|B
.print DEVI I_MERGE|I_Q1|B
.print DEVI B_MERGE|A1|1
.print DEVI L_MERGE|A1|P
.print DEVI R_MERGE|A1|B
.print DEVI L_MERGE|A1|RB
.print DEVI B_MERGE|A2|1
.print DEVI L_MERGE|A2|P
.print DEVI R_MERGE|A2|B
.print DEVI L_MERGE|A2|RB
.print DEVI B_MERGE|A12|1
.print DEVI R_MERGE|A12|B
.print DEVI L_MERGE|A12|RB
.print DEVI B_MERGE|B1|1
.print DEVI L_MERGE|B1|P
.print DEVI R_MERGE|B1|B
.print DEVI L_MERGE|B1|RB
.print DEVI B_MERGE|B2|1
.print DEVI L_MERGE|B2|P
.print DEVI R_MERGE|B2|B
.print DEVI L_MERGE|B2|RB
.print DEVI B_MERGE|B12|1
.print DEVI R_MERGE|B12|B
.print DEVI L_MERGE|B12|RB
.print DEVI B_MERGE|Q2|1
.print DEVI L_MERGE|Q2|P
.print DEVI R_MERGE|Q2|B
.print DEVI L_MERGE|Q2|RB
.print DEVI B_MERGE|Q1|1
.print DEVI L_MERGE|Q1|P
.print DEVI R_MERGE|Q1|B
.print DEVI L_MERGE|Q1|RB
.print DEVI L_XOR|I_A1|B
.print DEVI I_XOR|I_A1|B
.print DEVI L_XOR|I_A3|B
.print DEVI I_XOR|I_A3|B
.print DEVI L_XOR|I_B1|B
.print DEVI I_XOR|I_B1|B
.print DEVI L_XOR|I_B3|B
.print DEVI I_XOR|I_B3|B
.print DEVI L_XOR|I_T1|B
.print DEVI I_XOR|I_T1|B
.print DEVI L_XOR|I_Q1|B
.print DEVI I_XOR|I_Q1|B
.print DEVI B_XOR|A1|1
.print DEVI L_XOR|A1|P
.print DEVI R_XOR|A1|B
.print DEVI L_XOR|A1|RB
.print DEVI B_XOR|A2|1
.print DEVI L_XOR|A2|P
.print DEVI R_XOR|A2|B
.print DEVI L_XOR|A2|RB
.print DEVI B_XOR|A3|1
.print DEVI L_XOR|A3|P
.print DEVI R_XOR|A3|B
.print DEVI L_XOR|A3|RB
.print DEVI B_XOR|B1|1
.print DEVI L_XOR|B1|P
.print DEVI R_XOR|B1|B
.print DEVI L_XOR|B1|RB
.print DEVI B_XOR|B2|1
.print DEVI L_XOR|B2|P
.print DEVI R_XOR|B2|B
.print DEVI L_XOR|B2|RB
.print DEVI B_XOR|B3|1
.print DEVI L_XOR|B3|P
.print DEVI R_XOR|B3|B
.print DEVI L_XOR|B3|RB
.print DEVI B_XOR|T1|1
.print DEVI L_XOR|T1|P
.print DEVI R_XOR|T1|B
.print DEVI L_XOR|T1|RB
.print DEVI B_XOR|T2|1
.print DEVI R_XOR|T2|B
.print DEVI L_XOR|T2|RB
.print DEVI B_XOR|AB|1
.print DEVI L_XOR|AB|P
.print DEVI R_XOR|AB|B
.print DEVI L_XOR|AB|RB
.print DEVI B_XOR|ABTQ|1
.print DEVI L_XOR|ABTQ|P
.print DEVI R_XOR|ABTQ|B
.print DEVI L_XOR|ABTQ|RB
.print DEVI B_XOR|Q1|1
.print DEVI L_XOR|Q1|P
.print DEVI R_XOR|Q1|B
.print DEVI L_XOR|Q1|RB
.print V _XOR|B2
.print V _MERGE|A1|MID_SHUNT
.print V CLK
.print V _XOR|B3
.print V _XOR|B2|MID_SHUNT
.print V _MERGE|B1|MID_SHUNT
.print V _MERGE|B2
.print V _XOR|A2|MID_SERIES
.print V _MERGE|A2|MID_SERIES
.print V _MERGE|B2|MID_SERIES
.print V _XOR|A1
.print V _XOR|I_A3|MID
.print V _XOR|I_B1|MID
.print V _XOR|A2|MID_SHUNT
.print V _XOR|B3|MID_SHUNT
.print V _XOR|A1|MID_SERIES
.print V _XOR|A1|MID_SHUNT
.print V _XOR|B2|MID_SERIES
.print V _MERGE|B1
.print V _XOR|A3
.print V _MERGE|Q1|MID_SERIES
.print V _XOR|I_B3|MID
.print V _XOR|Q1|MID_SERIES
.print V _MERGE|I_B1|MID
.print V _XOR|A2
.print V _MERGE|I_Q1|MID
.print V _XOR|T1|MID_SHUNT
.print V _MERGE|A2|MID_SHUNT
.print V _MERGE|A1
.print V A
.print V _XOR|AB|MID_SERIES
.print V _MERGE|A3
.print V _MERGE|A1|MID_SERIES
.print V _XOR|T1|MID_SERIES
.print V _MERGE|Q2|MID_SERIES
.print V _XOR|Q1|MID_SHUNT
.print V Q
.print V A_OR_B
.print V _XOR|ABTQ|MID_SERIES
.print V _XOR|I_A1|MID
.print V _XOR|AB|MID_SHUNT
.print V _XOR|AB
.print V _XOR|T2
.print V _XOR|B3|MID_SERIES
.print V _MERGE|A2
.print V _XOR|B1
.print V _XOR|B1|MID_SHUNT
.print V _MERGE|I_Q3|MID
.print V _MERGE|B2|MID_SHUNT
.print V _MERGE|B12|MID_SHUNT
.print V _MERGE|B3
.print V _XOR|A3|MID_SERIES
.print V _XOR|A3|MID_SHUNT
.print V _MERGE|A12|MID_SHUNT
.print V B
.print V _MERGE|I_A1|MID
.print V _XOR|Q1
.print V _MERGE|B1|MID_SERIES
.print V C
.print V _MERGE|Q2
.print V _MERGE|Q1|MID_SHUNT
.print V _XOR|I_Q1|MID
.print V _XOR|T2|MID_SHUNT
.print V _XOR|ABTQ
.print V _XOR|T1
.print V _MERGE|Q2|MID_SHUNT
.print V _XOR|I_T1|MID
.print V _XOR|B1|MID_SERIES
.print V _MERGE|Q3
.print V _MERGE|I_Q2|MID
.print V _XOR|ABTQ|MID_SHUNT
.print V _MERGE|Q1
.print DEVP B_MERGE|A1|1
.print DEVP B_MERGE|A2|1
.print DEVP B_MERGE|A12|1
.print DEVP B_MERGE|B1|1
.print DEVP B_MERGE|B2|1
.print DEVP B_MERGE|B12|1
.print DEVP B_MERGE|Q2|1
.print DEVP B_MERGE|Q1|1
.print DEVP B_XOR|A1|1
.print DEVP B_XOR|A2|1
.print DEVP B_XOR|A3|1
.print DEVP B_XOR|B1|1
.print DEVP B_XOR|B2|1
.print DEVP B_XOR|B3|1
.print DEVP B_XOR|T1|1
.print DEVP B_XOR|T2|1
.print DEVP B_XOR|AB|1
.print DEVP B_XOR|ABTQ|1
.print DEVP B_XOR|Q1|1
