*
.include /Users/brainkz/Documents/GitHub/SFQ_gate_Exploration/jj_library.cir
.include /Users/brainkz/Documents/GitHub/SFQ/sunmagnetics_library.cir

* x_and a b t1 ab0 LSMITLL_AND_opt
* xjtl1  ab0 ab jtl
* x_xor ab c t2 abxc0 LSmitll_XOR_opt
* xjtl2  abxc0 abxc jtl
* ROUT  abxc  0  1  


.param offset1=5e-11
.param period=3e-10

Xt1      t1 clk_signal Tclk=period clk_offset=offset1 factor=4
Xdata_a  a  data_signal_a Tclk=period clk_offset=offset1
Xdata_b  b  data_signal_b Tclk=period clk_offset=offset1
Xdata_c  c  data_signal_c Tclk=period clk_offset=offset1+period


x_and_1 a b t1 ab0 LSMITLL_AND2
* Xc_delay c t1 cd0 dff

xd1 ab0 ab1 LSMITLL_BUFF
* xd2 cd0 cd1 LSMITLL_BUFF
xd3 ab1 ab  LSMITLL_JTL
* xd4 cd1 cd  LSMITLL_JTL

Xt2 t2 clk_signal clk_offset=0
x_xor ab c t2 abxc0 LSmitll_XOR_2
xjtlout  abxc0 abxc jtl
ROUT  abxc  0  1  


* Xc_delay c t1 c1 dff
* x_and a b t1 ab LSMITLL_AND_opt
* * xjtl1  ab0 ab1 jtl
* * xjtl2  ab1 ab2 jtl
* * xjtl3  ab2 ab3 jtl
* * xjtl4  ab1 ab  jtl
* x_xor ab c1 t2 abxc0 LSmitll_XOR_2
* xjtlout  abxc0 abxc jtl
* ROUT  abxc  0  1  

* Xt1 t1 clk_signal clk_offset=1e-10 factor=2
* Xdata_a  a data_signal_a clk_offset=1e-10
* Xdata_b  b data_signal_b clk_offset=1e-10

* Xt3 t2 clk_signal clk_offset=0
* Xdata_c  c data_signal_c clk_offset=1e-10

* * x_and a b t1 ab0 LSMITLL_AND_opt
* * xjtl1  ab0 ab jtl
* x_xor a b t1 ab0 xor 
* *LSmitll_XOR
* xjtl1  ab0 ab jtl
* ROUT  ab  0  1  

* .print DEVI ROUT

.tran 0.5e-12 6e-09

.end
* Ia   0    a    pwl(0 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 7.97e-10 0 8e-10 0.0005 8.03e-10 0 1.297e-09 0 1.3e-09 0.0005 1.303e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 2.297e-09 0 2.3e-09 0.0005 2.303e-09 0 2.797e-09 0 2.8e-09 0.0005 2.803e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.797e-09 0 3.8e-09 0.0005 3.803e-09 0 4.297e-09 0 4.3e-09 0.0005 4.303e-09 0 4.797e-09 0 4.8e-09 0.0005 4.803e-09 0 5.297e-09 0 5.3e-09 0.0005 5.303e-09 0 5.797e-09 0 5.8e-09 0.0005 5.803e-09 0 6.297e-09 0 6.3e-09 0.0005 6.303e-09 0 6.797e-09 0 6.8e-09 0.0005 6.803e-09 0 7.297e-09 0 7.3e-09 0.0005 7.303e-09 0 7.797e-09 0 7.8e-09 0.0005 7.803e-09 0)
* .print DEVI Ia

* Ib   0    b    pwl(0 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 8.47e-10 0 8.5e-10 0.0005 8.53e-10 0 1.597e-09 0 1.6e-09 0.0005 1.603e-09 0 1.847e-09 0 1.85e-09 0.0005 1.853e-09 0 2.597e-09 0 2.6e-09 0.0005 2.603e-09 0 2.847e-09 0 2.85e-09 0.0005 2.853e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.847e-09 0 3.85e-09 0.0005 3.853e-09 0 4.597e-09 0 4.6e-09 0.0005 4.603e-09 0 4.847e-09 0 4.85e-09 0.0005 4.853e-09 0 5.597e-09 0 5.6e-09 0.0005 5.603e-09 0 5.847e-09 0 5.85e-09 0.0005 5.853e-09 0 6.597e-09 0 6.6e-09 0.0005 6.603e-09 0 6.847e-09 0 6.85e-09 0.0005 6.853e-09 0 7.597e-09 0 7.6e-09 0.0005 7.603e-09 0 7.847e-09 0 7.85e-09 0.0005 7.853e-09 0)
* .print DEVI Ib

* Ic   0    c    pwl(0 0 1.147e-09 0 1.15e-09 0.0005 1.153e-09 0 1.397e-09 0 1.4e-09 0.0005 1.403e-09 0 1.647e-09 0 1.65e-09 0.0005 1.653e-09 0 1.897e-09 0 1.9e-09 0.0005 1.903e-09 0 3.147e-09 0 3.15e-09 0.0005 3.153e-09 0 3.397e-09 0 3.4e-09 0.0005 3.403e-09 0 3.647e-09 0 3.65e-09 0.0005 3.653e-09 0 3.897e-09 0 3.9e-09 0.0005 3.903e-09 0 5.147e-09 0 5.15e-09 0.0005 5.153e-09 0 5.397e-09 0 5.4e-09 0.0005 5.403e-09 0 5.647e-09 0 5.65e-09 0.0005 5.653e-09 0 5.897e-09 0 5.9e-09 0.0005 5.903e-09 0 7.147e-09 0 7.15e-09 0.0005 7.153e-09 0 7.397e-09 0 7.4e-09 0.0005 7.403e-09 0 7.647e-09 0 7.65e-09 0.0005 7.653e-09 0 7.897e-09 0 7.9e-09 0.0005 7.903e-09 0)
* .print DEVI Ic

* Id   0    d    pwl(0 0  2.197e-09 0 2.2000000000000003e-09 0.0005 2.2030000000000004e-09 0 2.447e-09 0 2.45e-09 0.0005 2.453e-09 0 2.697e-09 0 2.7e-09 0.0005 2.7030000000000003e-09 0 2.9470000000000003e-09 0 2.9500000000000004e-09 0.0005 2.9530000000000005e-09 0 3.197e-09 0 3.2e-09 0.0005 3.2030000000000002e-09 0 3.447e-09 0 3.4500000000000003e-09 0.0005 3.4530000000000004e-09 0 3.6970000000000004e-09 0 3.7000000000000005e-09 0.0005 3.7030000000000006e-09 0 3.9470000000000005e-09 0 3.950000000000001e-09 0.0005 3.953000000000001e-09 0 6.197000000000001e-09 0 6.200000000000001e-09 0.0005 6.203000000000001e-09 0 6.447000000000001e-09 0 6.450000000000001e-09 0.0005 6.453000000000001e-09 0 6.697e-09 0 6.7000000000000004e-09 0.0005 6.7030000000000005e-09 0 6.947000000000001e-09 0 6.950000000000001e-09 0.0005 6.953000000000001e-09 0 7.197000000000001e-09 0 7.200000000000001e-09 0.0005 7.203000000000001e-09 0 7.447000000000001e-09 0 7.450000000000001e-09 0.0005 7.453e-09 0 7.697e-09 0 7.7e-09 0.0005 7.703e-09 0 7.947e-09 0 7.95e-09 0.0005 7.953e-09 0 )
* .print DEVI Id



