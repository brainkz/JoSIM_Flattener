*
.include /Users/brainkz/Documents/GitHub/SFQ_gate_Exploration/jj_library.cir
.include /Users/brainkz/Documents/GitHub/SFQ/sunmagnetics_library.cir

* .param offset1=1e-10

* Xt1       t1  clk_signal    clk_offset=offset1 factor=8
* Xt2       t2  clk_signal    clk_offset=0       factor=2

* Xdata_a1  a1  data_signal_a clk_offset=offset1
* Xdata_b1  b1  data_signal_b clk_offset=offset1
* Xdata_c1  c1  data_signal_c clk_offset=offset1
* Xdata_d1  d1  data_signal_d clk_offset=offset1

* Xdata_a2  a2  data_signal_a clk_offset=offset1
* Xdata_b2  b2  data_signal_b clk_offset=offset1
* Xdata_c2  c2  data_signal_c clk_offset=offset1
* Xdata_d2  d2  data_signal_d clk_offset=offset1

* x_and_a1b1 a1 b1 t1 a1b1_0 LSMITLL_AND2
* x_and_c1d1 c1 d1 t1 c1d1_0 LSMITLL_AND2

* xd1 a1b1_0 a1b1_1 LSMITLL_BUFF
* xd2 c1d1_0 c1d1_1 LSMITLL_BUFF
* xd3 a1b1_1 a1b1  LSMITLL_JTL
* xd4 c1d1_1 c1d1  LSMITLL_JTL

* x_xor a1b1 c1d1 t2 a1b1xc1d1_0 LSmitll_XOR_2
* xjtlout  a1b1xc1d1_0 a1b1xc1d1 jtl

.param offset1=1e-10

.subckt ab_xor_cd a b c d t1 t2 out1 out2
    x_and_ab a b t1 ab_0 and2_clocked
    x_and_cd c d t1 cd_0 and2_clocked

    xd1 ab_0 ab_1 LSMITLL_BUFF
    xd2 cd_0 cd_1 LSMITLL_BUFF
    xd3 ab_1 ab   LSMITLL_JTL
    xd4 cd_1 cd   LSMITLL_JTL

    x_ab_spl ab abx abn LSmitll_SPLIT

    x_xor abx cd t2 abxcd  xor
    x_not abn    t2 not_ab LSMITLL_NOT
    xjtlout1  abxcd  out1 jtl
    xjtlout2  not_ab out2 jtl
.ends

Xt1       t1  clk_signal    clk_offset=offset1 factor=2
Xt2       t2  clk_signal    clk_offset=0       factor=2

Xdata_a1  a1  data_signal_a clk_offset=offset1
*  do_factor=0.1
Xdata_b1  b1  data_signal_b clk_offset=offset1
*  do_factor=0.1
Xdata_c1  c1  data_signal_c clk_offset=offset1
*  do_factor=0.1
Xdata_d1  d1  data_signal_d clk_offset=offset1
*  do_factor=0.1

* Xdata_a2  a2  data_signal_a clk_offset=offset1
* *  do_factor=0.1
* Xdata_b2  b2  data_signal_b clk_offset=offset1
* *  do_factor=0.1
* Xdata_c2  c2  data_signal_c clk_offset=offset1
* *  do_factor=0.1
* Xdata_d2  d2  data_signal_d clk_offset=offset1
* *  do_factor=0.1

x1 a1 b1 c1 d1 t1 t2 ab_xor_cd_1 not_ab_1 ab_xor_cd 
* not_ab_1
* x2 a2 b2 c2 d2 ab_xor_cd_2
* x2 d2 c2 b2 a2 t1 ab_xor_cd_2 ab_xor_cd

* x3 ab_xor_cd_1 ab_xor_cd_2 t2 out and2_clocked


ROUT1 ab_xor_cd_1  0  1  
ROUT2 not_ab_1  0  1  

.tran 0.5e-12 12e-09

.end
