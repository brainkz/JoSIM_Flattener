*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=5e-11
.PARAM PERIOD=3e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.5E-12 6E-09
ROUT ABXC 0  1
IT1|T 0 T1  PWL(0 0 3.47e-10 0 3.5e-10 0.002 3.53e-10 0 6.47e-10 0 6.5e-10 0.002 6.53e-10 0 9.47e-10 0 9.5e-10 0.002 9.53e-10 0 1.247e-09 0 1.25e-09 0.002 1.253e-09 0 1.547e-09 0 1.55e-09 0.002 1.553e-09 0 1.847e-09 0 1.85e-09 0.002 1.853e-09 0 2.147e-09 0 2.15e-09 0.002 2.153e-09 0 2.447e-09 0 2.45e-09 0.002 2.453e-09 0 2.747e-09 0 2.75e-09 0.002 2.753e-09 0 3.047e-09 0 3.05e-09 0.002 3.053e-09 0 3.347e-09 0 3.35e-09 0.002 3.353e-09 0 3.647e-09 0 3.65e-09 0.002 3.653e-09 0 3.947e-09 0 3.95e-09 0.002 3.953e-09 0 4.247e-09 0 4.25e-09 0.002 4.253e-09 0 4.547e-09 0 4.55e-09 0.002 4.553e-09 0 4.847e-09 0 4.85e-09 0.002 4.853e-09 0 5.147e-09 0 5.15e-09 0.002 5.153e-09 0 5.447e-09 0 5.45e-09 0.002 5.453e-09 0 5.747e-09 0 5.75e-09 0.002 5.753e-09 0 6.047e-09 0 6.05e-09 0.002 6.053e-09 0 6.347e-09 0 6.35e-09 0.002 6.353e-09 0 6.647e-09 0 6.65e-09 0.002 6.653e-09 0 6.947e-09 0 6.95e-09 0.002 6.953e-09 0 7.247e-09 0 7.25e-09 0.002 7.253e-09 0 7.547e-09 0 7.55e-09 0.002 7.553e-09 0 7.847e-09 0 7.85e-09 0.002 7.853e-09 0 8.147e-09 0 8.15e-09 0.002 8.153e-09 0 8.447e-09 0 8.45e-09 0.002 8.453e-09 0 8.747e-09 0 8.75e-09 0.002 8.753e-09 0 9.047e-09 0 9.05e-09 0.002 9.053e-09 0 9.347e-09 0 9.35e-09 0.002 9.353e-09 0 9.647e-09 0 9.65e-09 0.002 9.653e-09 0 9.947e-09 0 9.95e-09 0.002 9.953e-09 0 1.0247e-08 0 1.025e-08 0.002 1.0253e-08 0 1.0547e-08 0 1.055e-08 0.002 1.0553e-08 0 1.0847e-08 0 1.085e-08 0.002 1.0853e-08 0 1.1147e-08 0 1.115e-08 0.002 1.1153e-08 0 1.1447e-08 0 1.145e-08 0.002 1.1453e-08 0 1.1747e-08 0 1.175e-08 0.002 1.1753e-08 0)
IDATA_A|A 0 A  PWL(0 0 7.07e-10 0 7.1e-10 0.0005 7.13e-10 0 1.307e-09 0 1.31e-09 0.0005 1.313e-09 0 1.907e-09 0 1.91e-09 0.0005 1.913e-09 0 2.507e-09 0 2.51e-09 0.0005 2.513e-09 0 3.107e-09 0 3.11e-09 0.0005 3.113e-09 0 3.707e-09 0 3.71e-09 0.0005 3.713e-09 0 4.307e-09 0 4.31e-09 0.0005 4.313e-09 0 4.907e-09 0 4.91e-09 0.0005 4.913e-09 0 5.507e-09 0 5.51e-09 0.0005 5.513e-09 0 6.107e-09 0 6.11e-09 0.0005 6.113e-09 0 6.707e-09 0 6.71e-09 0.0005 6.713e-09 0 7.307e-09 0 7.31e-09 0.0005 7.313e-09 0 7.907e-09 0 7.91e-09 0.0005 7.913e-09 0 8.507e-09 0 8.51e-09 0.0005 8.513e-09 0 9.107e-09 0 9.11e-09 0.0005 9.113e-09 0 9.707e-09 0 9.71e-09 0.0005 9.713e-09 0 1.0307e-08 0 1.031e-08 0.0005 1.0313e-08 0 1.0907e-08 0 1.091e-08 0.0005 1.0913e-08 0 1.1507e-08 0 1.151e-08 0.0005 1.1513e-08 0)
IDATA_B|B 0 B  PWL(0 0 1.067e-09 0 1.07e-09 0.0005 1.073e-09 0 1.367e-09 0 1.37e-09 0.0005 1.373e-09 0 2.267e-09 0 2.27e-09 0.0005 2.273e-09 0 2.567e-09 0 2.57e-09 0.0005 2.573e-09 0 3.467e-09 0 3.47e-09 0.0005 3.473e-09 0 3.767e-09 0 3.77e-09 0.0005 3.773e-09 0 4.667e-09 0 4.67e-09 0.0005 4.673e-09 0 4.967e-09 0 4.97e-09 0.0005 4.973e-09 0 5.867e-09 0 5.87e-09 0.0005 5.873e-09 0 6.167e-09 0 6.17e-09 0.0005 6.173e-09 0 7.067e-09 0 7.07e-09 0.0005 7.073e-09 0 7.367e-09 0 7.37e-09 0.0005 7.373e-09 0 8.267e-09 0 8.27e-09 0.0005 8.273e-09 0 8.567e-09 0 8.57e-09 0.0005 8.573e-09 0 9.467e-09 0 9.47e-09 0.0005 9.473e-09 0 9.767e-09 0 9.77e-09 0.0005 9.773e-09 0 1.0667e-08 0 1.067e-08 0.0005 1.0673e-08 0 1.0967e-08 0 1.097e-08 0.0005 1.0973e-08 0 1.1867e-08 0 1.187e-08 0.0005 1.1873e-08 0)
IDATA_C|T 0 C  PWL(0 0 2.027e-09 0 2.03e-09 0.0005 2.033e-09 0 2.327e-09 0 2.33e-09 0.0005 2.333e-09 0 2.627e-09 0 2.63e-09 0.0005 2.633e-09 0 2.927e-09 0 2.93e-09 0.0005 2.933e-09 0 4.427e-09 0 4.43e-09 0.0005 4.433e-09 0 4.727e-09 0 4.73e-09 0.0005 4.733e-09 0 5.027e-09 0 5.03e-09 0.0005 5.033e-09 0 5.327e-09 0 5.33e-09 0.0005 5.333e-09 0 6.827e-09 0 6.83e-09 0.0005 6.833e-09 0 7.127e-09 0 7.13e-09 0.0005 7.133e-09 0 7.427e-09 0 7.43e-09 0.0005 7.433e-09 0 7.727e-09 0 7.73e-09 0.0005 7.733e-09 0 9.227e-09 0 9.23e-09 0.0005 9.233e-09 0 9.527e-09 0 9.53e-09 0.0005 9.533e-09 0 9.827e-09 0 9.83e-09 0.0005 9.833e-09 0 1.0127e-08 0 1.013e-08 0.0005 1.0133e-08 0 1.1627e-08 0 1.163e-08 0.0005 1.1633e-08 0 1.1927e-08 0 1.193e-08 0.0005 1.1933e-08 0 1.2227e-08 0 1.223e-08 0.0005 1.2233e-08 0)
B_AND_1|1 _AND_1|1 _AND_1|2 JJMIT AREA=2.5
B_AND_1|2 _AND_1|4 _AND_1|5 JJMIT AREA=1.7857142857142858
B_AND_1|3 _AND_1|5 _AND_1|6 JJMIT AREA=2.5
B_AND_1|4 _AND_1|8 _AND_1|9 JJMIT AREA=1.7857142857142858
B_AND_1|5 _AND_1|8 _AND_1|11 JJMIT AREA=2.5
B_AND_1|6 _AND_1|12 _AND_1|13 JJMIT AREA=1.7857142857142858
B_AND_1|7 _AND_1|14 _AND_1|15 JJMIT AREA=2.5
B_AND_1|8 _AND_1|17 _AND_1|18 JJMIT AREA=1.7857142857142858
B_AND_1|9 _AND_1|18 _AND_1|19 JJMIT AREA=2.5
B_AND_1|10 _AND_1|21 _AND_1|22 JJMIT AREA=1.7857142857142858
B_AND_1|11 _AND_1|21 _AND_1|23 JJMIT AREA=2.5
B_AND_1|12 _AND_1|24 _AND_1|13 JJMIT AREA=1.7857142857142858
B_AND_1|13 _AND_1|25 _AND_1|26 JJMIT AREA=2.5
B_AND_1|14 _AND_1|31 _AND_1|32 JJMIT AREA=2.5
B_AND_1|15 _AND_1|28 _AND_1|29 JJMIT AREA=2.5
I_AND_1|B1 0 _AND_1|3  PWL(0 0 5e-12 0.000175)
I_AND_1|B2 0 _AND_1|7  PWL(0 0 5e-12 0.000175)
I_AND_1|B3 0 _AND_1|16  PWL(0 0 5e-12 0.000175)
I_AND_1|B4 0 _AND_1|20  PWL(0 0 5e-12 0.000175)
I_AND_1|B5 0 _AND_1|27  PWL(0 0 5e-12 0.000175)
I_AND_1|B6 0 _AND_1|33  PWL(0 0 5e-12 0.000175)
I_AND_1|B7 0 _AND_1|30  PWL(0 0 5e-12 0.000175)
L_AND_1|B1 _AND_1|3 _AND_1|1  2e-12
L_AND_1|B2 _AND_1|7 _AND_1|5  2e-12
L_AND_1|B3 _AND_1|16 _AND_1|14  2e-12
L_AND_1|B4 _AND_1|20 _AND_1|18  2e-12
L_AND_1|B5 _AND_1|27 _AND_1|25  2e-12
L_AND_1|B6 _AND_1|30 _AND_1|28  2e-12
L_AND_1|B7 _AND_1|33 _AND_1|31  2e-12
L_AND_1|P1 _AND_1|2 0  2e-13
L_AND_1|P3 _AND_1|6 0  2e-13
L_AND_1|P5 _AND_1|11 0  2e-13
L_AND_1|P7 _AND_1|15 0  2e-13
L_AND_1|P9 _AND_1|19 0  2e-13
L_AND_1|P11 _AND_1|23 0  2e-13
L_AND_1|P13 _AND_1|26 0  2e-13
L_AND_1|P14 _AND_1|32 0  2e-13
L_AND_1|P15 _AND_1|29 0  2e-13
L_AND_1|1 A _AND_1|1  2.067833848e-12
L_AND_1|2 _AND_1|1 _AND_1|4  4.135667696e-12
L_AND_1|3 _AND_1|5 _AND_1|8  8.271335392e-12
L_AND_1|4 _AND_1|9 _AND_1|10  1e-12
L_AND_1|5 _AND_1|8 _AND_1|12  4.135667696e-12
L_AND_1|6 B _AND_1|14  2.067833848e-12
L_AND_1|7 _AND_1|14 _AND_1|17  4.135667696e-12
L_AND_1|8 _AND_1|18 _AND_1|21  8.271335392e-12
L_AND_1|9 _AND_1|22 _AND_1|10  1e-12
L_AND_1|10 _AND_1|21 _AND_1|24  4.135667696e-12
L_AND_1|11 T1 _AND_1|25  2.067833848e-12
L_AND_1|12 _AND_1|25 _AND_1|31  4.135667696e-12
L_AND_1|13 _AND_1|31 _AND_1|10  1e-12
L_AND_1|14 _AND_1|13 _AND_1|28  1e-12
L_AND_1|15 _AND_1|28 AB0  2.067833848e-12
R_AND_1|B1 _AND_1|1 _AND_1|101  2.7439617672
L_AND_1|RB1 _AND_1|101 0  1.550338398468e-12
R_AND_1|B2 _AND_1|4 _AND_1|104  3.84154647408
L_AND_1|RB2 _AND_1|104 _AND_1|5  2.1704737578552e-12
R_AND_1|B3 _AND_1|5 _AND_1|105  2.7439617672
L_AND_1|RB3 _AND_1|105 0  1.550338398468e-12
R_AND_1|B4 _AND_1|8 _AND_1|109  3.84154647408
L_AND_1|RB4 _AND_1|109 _AND_1|9  2.1704737578552e-12
R_AND_1|B5 _AND_1|8 _AND_1|108  2.7439617672
L_AND_1|RB5 _AND_1|108 0  1.550338398468e-12
R_AND_1|B6 _AND_1|12 _AND_1|112  3.84154647408
L_AND_1|RB6 _AND_1|112 _AND_1|13  2.1704737578552e-12
R_AND_1|B7 _AND_1|14 _AND_1|114  2.7439617672
L_AND_1|RB7 _AND_1|114 0  1.550338398468e-12
R_AND_1|B8 _AND_1|17 _AND_1|117  3.84154647408
L_AND_1|RB8 _AND_1|117 _AND_1|18  2.1704737578552e-12
R_AND_1|B9 _AND_1|18 _AND_1|118  2.7439617672
L_AND_1|RB9 _AND_1|118 0  1.550338398468e-12
R_AND_1|B10 _AND_1|21 _AND_1|122  3.84154647408
L_AND_1|RB10 _AND_1|122 _AND_1|22  2.1704737578552e-12
R_AND_1|B11 _AND_1|21 _AND_1|121  2.7439617672
L_AND_1|RB11 _AND_1|121 0  1.550338398468e-12
R_AND_1|B12 _AND_1|24 _AND_1|124  3.84154647408
L_AND_1|RB12 _AND_1|124 _AND_1|13  2.1704737578552e-12
R_AND_1|B13 _AND_1|25 _AND_1|125  2.7439617672
L_AND_1|RB13 _AND_1|125 0  1.550338398468e-12
R_AND_1|B14 _AND_1|31 _AND_1|131  2.7439617672
L_AND_1|RB14 _AND_1|131 0  1.550338398468e-12
R_AND_1|B15 _AND_1|28 _AND_1|128  2.7439617672
L_AND_1|RB15 _AND_1|128 0  1.550338398468e-12
BD1|1 D1|1 D1|2 JJMIT AREA=2.5
BD1|2 D1|4 D1|5 JJMIT AREA=2.5
BD1|3 D1|7 D1|8 JJMIT AREA=2.5
BD1|4 D1|10 D1|11 JJMIT AREA=2.5
ID1|B1 0 D1|3  PWL(0 0 5e-12 0.000175)
ID1|B2 0 D1|6  PWL(0 0 5e-12 0.0002375)
ID1|B3 0 D1|9  PWL(0 0 5e-12 0.0002375)
ID1|B4 0 D1|12  PWL(0 0 5e-12 0.000175)
LD1|1 AB0 D1|1  2.067833848e-12
LD1|2 D1|1 D1|4  4.135667696e-12
LD1|3 D1|4 D1|7  4.135667696e-12
LD1|4 D1|7 D1|10  4.135667696e-12
LD1|5 D1|10 AB1  2.067833848e-12
LD1|P1 D1|2 0  5e-13
LD1|P2 D1|5 0  5e-13
LD1|P3 D1|8 0  5e-13
LD1|P4 D1|11 0  5e-13
LD1|B1 D1|1 D1|3  2e-12
LD1|B2 D1|4 D1|6  2e-12
LD1|B3 D1|7 D1|9  2e-12
LD1|B4 D1|10 D1|12  2e-12
RD1|B1 D1|1 D1|101  2.7439617672
RD1|B2 D1|4 D1|104  2.7439617672
RD1|B3 D1|7 D1|107  2.7439617672
RD1|B4 D1|10 D1|110  2.7439617672
LD1|RB1 D1|101 0  2.050338398468e-12
LD1|RB2 D1|104 0  2.050338398468e-12
LD1|RB3 D1|107 0  2.050338398468e-12
LD1|RB4 D1|110 0  2.050338398468e-12
BD3|1 D3|1 D3|2 JJMIT AREA=2.5
BD3|2 D3|6 D3|7 JJMIT AREA=2.5
ID3|B1 0 D3|5  0.00035
LD3|1 AB1 D3|1  2.067833848e-12
LD3|2 D3|1 D3|4  2.067833848e-12
LD3|3 D3|4 D3|6  2.067833848e-12
LD3|4 D3|6 AB  2.067833848e-12
LD3|P1 D3|2 0  2e-13
LD3|P2 D3|7 0  2e-13
LD3|B1 D3|5 D3|4  2e-12
RD3|B1 D3|1 D3|3  2.7439617672
RD3|B2 D3|6 D3|8  2.7439617672
LD3|RB1 D3|3 0  1.750338398468e-12
LD3|RB2 D3|8 0  1.750338398468e-12
IT2|T 0 T2  PWL(0 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.897e-09 0 3.9e-09 0.0005 3.903e-09 0 4.197e-09 0 4.2e-09 0.0005 4.203e-09 0 4.497e-09 0 4.5e-09 0.0005 4.503e-09 0 4.797e-09 0 4.8e-09 0.0005 4.803e-09 0 5.097e-09 0 5.1e-09 0.0005 5.103e-09 0 5.397e-09 0 5.4e-09 0.0005 5.403e-09 0 5.697e-09 0 5.7e-09 0.0005 5.703e-09 0 5.997e-09 0 6e-09 0.0005 6.003e-09 0 6.297e-09 0 6.3e-09 0.0005 6.303e-09 0 6.597e-09 0 6.6e-09 0.0005 6.603e-09 0 6.897e-09 0 6.9e-09 0.0005 6.903e-09 0 7.197e-09 0 7.2e-09 0.0005 7.203e-09 0 7.497e-09 0 7.5e-09 0.0005 7.503e-09 0 7.797e-09 0 7.8e-09 0.0005 7.803e-09 0 8.097e-09 0 8.1e-09 0.0005 8.103e-09 0 8.397e-09 0 8.4e-09 0.0005 8.403e-09 0 8.697e-09 0 8.7e-09 0.0005 8.703e-09 0 8.997e-09 0 9e-09 0.0005 9.003e-09 0 9.297e-09 0 9.3e-09 0.0005 9.303e-09 0 9.597e-09 0 9.6e-09 0.0005 9.603e-09 0 9.897e-09 0 9.9e-09 0.0005 9.903e-09 0 1.0197e-08 0 1.02e-08 0.0005 1.0203e-08 0 1.0497e-08 0 1.05e-08 0.0005 1.0503e-08 0 1.0797e-08 0 1.08e-08 0.0005 1.0803e-08 0 1.1097e-08 0 1.11e-08 0.0005 1.1103e-08 0 1.1397e-08 0 1.14e-08 0.0005 1.1403e-08 0 1.1697e-08 0 1.17e-08 0.0005 1.1703e-08 0)
B_XOR|1 _XOR|1 _XOR|2 JJMIT AREA=2.5
B_XOR|2 _XOR|4 _XOR|5 JJMIT AREA=2.5
B_XOR|3 _XOR|25 _XOR|6 JJMIT AREA=2.5
B_XOR|4 _XOR|9 _XOR|10 JJMIT AREA=2.5
B_XOR|5 _XOR|12 _XOR|13 JJMIT AREA=2.5
B_XOR|6 _XOR|26 _XOR|14 JJMIT AREA=2.5
B_XOR|7 _XOR|27 _XOR|16 JJMIT AREA=2.0
B_XOR|8 _XOR|17 _XOR|18 JJMIT AREA=2.5
B_XOR|9 _XOR|20 _XOR|16 JJMIT AREA=2.0
B_XOR|10 _XOR|16 _XOR|21 JJMIT AREA=2.5
B_XOR|11 _XOR|22 _XOR|23 JJMIT AREA=2.5
I_XOR|B1 0 _XOR|3  0.00017499999999999997
I_XOR|B2 0 _XOR|7  0.00017499999999999997
I_XOR|B3 0 _XOR|11  0.00017499999999999997
I_XOR|B4 0 _XOR|15  0.00017499999999999997
I_XOR|B5 0 _XOR|19  0.00017499999999999997
I_XOR|B6 0 _XOR|24  0.00017499999999999997
L_XOR|B1 _XOR|3 _XOR|1  2e-12
L_XOR|B2 _XOR|7 _XOR|6  2e-12
L_XOR|B3 _XOR|11 _XOR|9  2e-12
L_XOR|B4 _XOR|15 _XOR|14  2e-12
L_XOR|B5 _XOR|19 _XOR|17  2e-12
L_XOR|B6 _XOR|24 _XOR|22  2e-12
L_XOR|1 AB _XOR|1  2.067833848e-12
L_XOR|2 _XOR|1 _XOR|4  4.135667696e-12
L_XOR|3 _XOR|4 _XOR|25  1.2e-12
L_XOR|4 _XOR|6 _XOR|8  8.271335392e-12
L_XOR|5 C _XOR|9  2.067833848e-12
L_XOR|6 _XOR|9 _XOR|12  4.135667696e-12
L_XOR|7 _XOR|12 _XOR|26  1.2e-12
L_XOR|8 _XOR|14 _XOR|8  8.271335392e-12
L_XOR|9 _XOR|8 _XOR|27  1.2e-12
L_XOR|10 T2 _XOR|17  2.067833848e-12
L_XOR|11 _XOR|17 _XOR|20  4.135667696e-12
L_XOR|12 _XOR|16 _XOR|22  4.135667696e-12
L_XOR|13 _XOR|22 ABXC0  2.067833848e-12
L_XOR|P1 _XOR|2 0  5e-13
L_XOR|P2 _XOR|5 0  5e-13
L_XOR|P4 _XOR|10 0  5e-13
L_XOR|P5 _XOR|13 0  5e-13
L_XOR|P8 _XOR|18 0  5e-13
L_XOR|P10 _XOR|21 0  5e-13
L_XOR|P11 _XOR|23 0  5e-13
R_XOR|B1 _XOR|1 _XOR|101  2.7439617672
L_XOR|RB1 _XOR|101 0  2.050338398468e-12
R_XOR|B2 _XOR|4 _XOR|104  2.7439617672
L_XOR|RB2 _XOR|104 0  2.050338398468e-12
R_XOR|B3 _XOR|4 _XOR|106  2.7439617672
L_XOR|RB3 _XOR|106 _XOR|6  2.050338398468e-12
R_XOR|B4 _XOR|9 _XOR|109  2.7439617672
L_XOR|RB4 _XOR|109 0  2.050338398468e-12
R_XOR|B5 _XOR|12 _XOR|112  2.7439617672
L_XOR|RB5 _XOR|112 0  2.050338398468e-12
R_XOR|B6 _XOR|12 _XOR|114  2.7439617672
L_XOR|RB6 _XOR|114 _XOR|14  2.050338398468e-12
R_XOR|B7 _XOR|8 _XOR|108  3.429952209
L_XOR|RB7 _XOR|108 _XOR|16  2.437922998085e-12
R_XOR|B8 _XOR|17 _XOR|117  2.7439617672
L_XOR|RB8 _XOR|117 0  2.050338398468e-12
R_XOR|B9 _XOR|20 _XOR|120  3.429952209
L_XOR|RB9 _XOR|120 _XOR|16  2.437922998085e-12
R_XOR|B10 _XOR|16 _XOR|116  2.7439617672
L_XOR|RB10 _XOR|116 0  2.050338398468e-12
R_XOR|B11 _XOR|22 _XOR|122  2.7439617672
L_XOR|RB11 _XOR|122 0  2.050338398468e-12
LJTLOUT|1 ABXC0 JTLOUT|1  2.067833848e-12
LJTLOUT|2 JTLOUT|1 JTLOUT|4  2.067833848e-12
LJTLOUT|3 JTLOUT|4 JTLOUT|6  2.067833848e-12
LJTLOUT|4 JTLOUT|6 ABXC  2.067833848e-12
BJTLOUT|1|1 JTLOUT|1 JTLOUT|1|MID_SERIES JJMIT AREA=2.5
LJTLOUT|1|P JTLOUT|1|MID_SERIES 0  2e-13
RJTLOUT|1|B JTLOUT|1 JTLOUT|1|MID_SHUNT  2.7439617672
LJTLOUT|1|RB JTLOUT|1|MID_SHUNT 0  1.750338398468e-12
LJTLOUT|B|B JTLOUT|4 JTLOUT|B|MID  2e-12
IJTLOUT|B|B 0 JTLOUT|B|MID  0.0005
BJTLOUT|2|1 JTLOUT|6 JTLOUT|2|MID_SERIES JJMIT AREA=2.5
LJTLOUT|2|P JTLOUT|2|MID_SERIES 0  2e-13
RJTLOUT|2|B JTLOUT|6 JTLOUT|2|MID_SHUNT  2.7439617672
LJTLOUT|2|RB JTLOUT|2|MID_SHUNT 0  1.750338398468e-12
.print DEVI ROUT
.print DEVI IT1|T
.print DEVI IDATA_A|A
.print DEVI IDATA_B|B
.print DEVI IDATA_C|T
.print DEVI B_AND_1|1
.print DEVI B_AND_1|2
.print DEVI B_AND_1|3
.print DEVI B_AND_1|4
.print DEVI B_AND_1|5
.print DEVI B_AND_1|6
.print DEVI B_AND_1|7
.print DEVI B_AND_1|8
.print DEVI B_AND_1|9
.print DEVI B_AND_1|10
.print DEVI B_AND_1|11
.print DEVI B_AND_1|12
.print DEVI B_AND_1|13
.print DEVI B_AND_1|14
.print DEVI B_AND_1|15
.print DEVI I_AND_1|B1
.print DEVI I_AND_1|B2
.print DEVI I_AND_1|B3
.print DEVI I_AND_1|B4
.print DEVI I_AND_1|B5
.print DEVI I_AND_1|B6
.print DEVI I_AND_1|B7
.print DEVI L_AND_1|B1
.print DEVI L_AND_1|B2
.print DEVI L_AND_1|B3
.print DEVI L_AND_1|B4
.print DEVI L_AND_1|B5
.print DEVI L_AND_1|B6
.print DEVI L_AND_1|B7
.print DEVI L_AND_1|P1
.print DEVI L_AND_1|P3
.print DEVI L_AND_1|P5
.print DEVI L_AND_1|P7
.print DEVI L_AND_1|P9
.print DEVI L_AND_1|P11
.print DEVI L_AND_1|P13
.print DEVI L_AND_1|P14
.print DEVI L_AND_1|P15
.print DEVI L_AND_1|1
.print DEVI L_AND_1|2
.print DEVI L_AND_1|3
.print DEVI L_AND_1|4
.print DEVI L_AND_1|5
.print DEVI L_AND_1|6
.print DEVI L_AND_1|7
.print DEVI L_AND_1|8
.print DEVI L_AND_1|9
.print DEVI L_AND_1|10
.print DEVI L_AND_1|11
.print DEVI L_AND_1|12
.print DEVI L_AND_1|13
.print DEVI L_AND_1|14
.print DEVI L_AND_1|15
.print DEVI R_AND_1|B1
.print DEVI L_AND_1|RB1
.print DEVI R_AND_1|B2
.print DEVI L_AND_1|RB2
.print DEVI R_AND_1|B3
.print DEVI L_AND_1|RB3
.print DEVI R_AND_1|B4
.print DEVI L_AND_1|RB4
.print DEVI R_AND_1|B5
.print DEVI L_AND_1|RB5
.print DEVI R_AND_1|B6
.print DEVI L_AND_1|RB6
.print DEVI R_AND_1|B7
.print DEVI L_AND_1|RB7
.print DEVI R_AND_1|B8
.print DEVI L_AND_1|RB8
.print DEVI R_AND_1|B9
.print DEVI L_AND_1|RB9
.print DEVI R_AND_1|B10
.print DEVI L_AND_1|RB10
.print DEVI R_AND_1|B11
.print DEVI L_AND_1|RB11
.print DEVI R_AND_1|B12
.print DEVI L_AND_1|RB12
.print DEVI R_AND_1|B13
.print DEVI L_AND_1|RB13
.print DEVI R_AND_1|B14
.print DEVI L_AND_1|RB14
.print DEVI R_AND_1|B15
.print DEVI L_AND_1|RB15
.print DEVI BD1|1
.print DEVI BD1|2
.print DEVI BD1|3
.print DEVI BD1|4
.print DEVI ID1|B1
.print DEVI ID1|B2
.print DEVI ID1|B3
.print DEVI ID1|B4
.print DEVI LD1|1
.print DEVI LD1|2
.print DEVI LD1|3
.print DEVI LD1|4
.print DEVI LD1|5
.print DEVI LD1|P1
.print DEVI LD1|P2
.print DEVI LD1|P3
.print DEVI LD1|P4
.print DEVI LD1|B1
.print DEVI LD1|B2
.print DEVI LD1|B3
.print DEVI LD1|B4
.print DEVI RD1|B1
.print DEVI RD1|B2
.print DEVI RD1|B3
.print DEVI RD1|B4
.print DEVI LD1|RB1
.print DEVI LD1|RB2
.print DEVI LD1|RB3
.print DEVI LD1|RB4
.print DEVI BD3|1
.print DEVI BD3|2
.print DEVI ID3|B1
.print DEVI LD3|1
.print DEVI LD3|2
.print DEVI LD3|3
.print DEVI LD3|4
.print DEVI LD3|P1
.print DEVI LD3|P2
.print DEVI LD3|B1
.print DEVI RD3|B1
.print DEVI RD3|B2
.print DEVI LD3|RB1
.print DEVI LD3|RB2
.print DEVI IT2|T
.print DEVI B_XOR|1
.print DEVI B_XOR|2
.print DEVI B_XOR|3
.print DEVI B_XOR|4
.print DEVI B_XOR|5
.print DEVI B_XOR|6
.print DEVI B_XOR|7
.print DEVI B_XOR|8
.print DEVI B_XOR|9
.print DEVI B_XOR|10
.print DEVI B_XOR|11
.print DEVI I_XOR|B1
.print DEVI I_XOR|B2
.print DEVI I_XOR|B3
.print DEVI I_XOR|B4
.print DEVI I_XOR|B5
.print DEVI I_XOR|B6
.print DEVI L_XOR|B1
.print DEVI L_XOR|B2
.print DEVI L_XOR|B3
.print DEVI L_XOR|B4
.print DEVI L_XOR|B5
.print DEVI L_XOR|B6
.print DEVI L_XOR|1
.print DEVI L_XOR|2
.print DEVI L_XOR|3
.print DEVI L_XOR|4
.print DEVI L_XOR|5
.print DEVI L_XOR|6
.print DEVI L_XOR|7
.print DEVI L_XOR|8
.print DEVI L_XOR|9
.print DEVI L_XOR|10
.print DEVI L_XOR|11
.print DEVI L_XOR|12
.print DEVI L_XOR|13
.print DEVI L_XOR|P1
.print DEVI L_XOR|P2
.print DEVI L_XOR|P4
.print DEVI L_XOR|P5
.print DEVI L_XOR|P8
.print DEVI L_XOR|P10
.print DEVI L_XOR|P11
.print DEVI R_XOR|B1
.print DEVI L_XOR|RB1
.print DEVI R_XOR|B2
.print DEVI L_XOR|RB2
.print DEVI R_XOR|B3
.print DEVI L_XOR|RB3
.print DEVI R_XOR|B4
.print DEVI L_XOR|RB4
.print DEVI R_XOR|B5
.print DEVI L_XOR|RB5
.print DEVI R_XOR|B6
.print DEVI L_XOR|RB6
.print DEVI R_XOR|B7
.print DEVI L_XOR|RB7
.print DEVI R_XOR|B8
.print DEVI L_XOR|RB8
.print DEVI R_XOR|B9
.print DEVI L_XOR|RB9
.print DEVI R_XOR|B10
.print DEVI L_XOR|RB10
.print DEVI R_XOR|B11
.print DEVI L_XOR|RB11
.print DEVI LJTLOUT|1
.print DEVI LJTLOUT|2
.print DEVI LJTLOUT|3
.print DEVI LJTLOUT|4
.print DEVI BJTLOUT|1|1
.print DEVI LJTLOUT|1|P
.print DEVI RJTLOUT|1|B
.print DEVI LJTLOUT|1|RB
.print DEVI LJTLOUT|B|B
.print DEVI IJTLOUT|B|B
.print DEVI BJTLOUT|2|1
.print DEVI LJTLOUT|2|P
.print DEVI RJTLOUT|2|B
.print DEVI LJTLOUT|2|RB
.print V JTLOUT|1|MID_SERIES
.print V _XOR|25
.print V _XOR|8
.print V _XOR|27
.print V _AND_1|30
.print V _AND_1|118
.print V _XOR|6
.print V AB1
.print V ABXC0
.print V _AND_1|9
.print V _XOR|17
.print V _AND_1|117
.print V AB0
.print V A
.print V _XOR|19
.print V _XOR|117
.print V D3|6
.print V T1
.print V _AND_1|7
.print V _AND_1|21
.print V ABXC
.print V _XOR|108
.print V _AND_1|27
.print V D1|6
.print V JTLOUT|1
.print V _XOR|116
.print V _AND_1|8
.print V _AND_1|105
.print V _AND_1|131
.print V D1|1
.print V _XOR|9
.print V D1|110
.print V _XOR|10
.print V D1|101
.print V _XOR|26
.print V JTLOUT|4
.print V _AND_1|114
.print V _AND_1|11
.print V D1|4
.print V _XOR|24
.print V _AND_1|16
.print V C
.print V D1|5
.print V _AND_1|32
.print V _XOR|120
.print V _AND_1|124
.print V JTLOUT|2|MID_SHUNT
.print V _XOR|14
.print V _AND_1|125
.print V _XOR|101
.print V _XOR|16
.print V _XOR|22
.print V _AND_1|23
.print V _AND_1|14
.print V D1|12
.print V _AND_1|109
.print V _XOR|112
.print V T2
.print V D1|2
.print V D3|5
.print V _AND_1|29
.print V _XOR|13
.print V D3|3
.print V D1|107
.print V B
.print V D1|11
.print V _XOR|21
.print V _AND_1|24
.print V _XOR|15
.print V D3|4
.print V _AND_1|121
.print V AB
.print V _XOR|23
.print V _XOR|7
.print V _AND_1|28
.print V _XOR|5
.print V _AND_1|3
.print V _XOR|11
.print V _XOR|3
.print V JTLOUT|2|MID_SERIES
.print V _AND_1|4
.print V _AND_1|20
.print V _AND_1|128
.print V _AND_1|33
.print V D1|7
.print V _AND_1|2
.print V _XOR|106
.print V JTLOUT|B|MID
.print V _AND_1|13
.print V _AND_1|10
.print V _AND_1|101
.print V D1|3
.print V _XOR|20
.print V _AND_1|122
.print V _AND_1|17
.print V D1|8
.print V D3|1
.print V _XOR|122
.print V _AND_1|22
.print V _AND_1|104
.print V _XOR|18
.print V JTLOUT|1|MID_SHUNT
.print V _XOR|4
.print V D1|9
.print V D3|8
.print V _XOR|2
.print V _AND_1|31
.print V _XOR|114
.print V _AND_1|15
.print V _AND_1|19
.print V _AND_1|112
.print V D1|10
.print V _XOR|12
.print V _XOR|109
.print V _AND_1|25
.print V _AND_1|18
.print V _XOR|1
.print V JTLOUT|6
.print V _AND_1|5
.print V _AND_1|12
.print V _AND_1|26
.print V _XOR|104
.print V _AND_1|6
.print V D1|104
.print V D3|2
.print V D3|7
.print V _AND_1|108
.print V _AND_1|1
.print DEVP B_AND_1|1
.print DEVP B_AND_1|2
.print DEVP B_AND_1|3
.print DEVP B_AND_1|4
.print DEVP B_AND_1|5
.print DEVP B_AND_1|6
.print DEVP B_AND_1|7
.print DEVP B_AND_1|8
.print DEVP B_AND_1|9
.print DEVP B_AND_1|10
.print DEVP B_AND_1|11
.print DEVP B_AND_1|12
.print DEVP B_AND_1|13
.print DEVP B_AND_1|14
.print DEVP B_AND_1|15
.print DEVP BD1|1
.print DEVP BD1|2
.print DEVP BD1|3
.print DEVP BD1|4
.print DEVP BD3|1
.print DEVP BD3|2
.print DEVP B_XOR|1
.print DEVP B_XOR|2
.print DEVP B_XOR|3
.print DEVP B_XOR|4
.print DEVP B_XOR|5
.print DEVP B_XOR|6
.print DEVP B_XOR|7
.print DEVP B_XOR|8
.print DEVP B_XOR|9
.print DEVP B_XOR|10
.print DEVP B_XOR|11
.print DEVP BJTLOUT|1|1
.print DEVP BJTLOUT|2|1
