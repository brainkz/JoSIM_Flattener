*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM TCLOCK=6e-11
.PARAM OS=3e-12
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 17000E-12
R_S0 S0 0  1
R_S1 S1 0  1
R_S2 S2 0  1
R_S3 S3 0  1
R_S4 S4 0  1
IA0|A 0 A0_TX  PWL(0 0 7.38e-11 0 7.68e-11 0.0007 7.98e-11 0 1.938e-10 0 1.968e-10 0.0007 1.998e-10 0 3.138e-10 0 3.168e-10 0.0007 3.198e-10 0 4.338e-10 0 4.368e-10 0.0007 4.398e-10 0 5.538e-10 0 5.568e-10 0.0007 5.598e-10 0 6.738e-10 0 6.768e-10 0.0007 6.798e-10 0 7.938e-10 0 7.968e-10 0.0007 7.998e-10 0 9.138e-10 0 9.168e-10 0.0007 9.198e-10 0 1.0338e-09 0 1.0368e-09 0.0007 1.0398e-09 0 1.1538e-09 0 1.1568e-09 0.0007 1.1598e-09 0 1.2738e-09 0 1.2768e-09 0.0007 1.2798e-09 0 1.3938e-09 0 1.3968e-09 0.0007 1.3998e-09 0 1.5138e-09 0 1.5168e-09 0.0007 1.5198e-09 0 1.6338e-09 0 1.6368e-09 0.0007 1.6398e-09 0 1.7538e-09 0 1.7568e-09 0.0007 1.7598e-09 0 1.8738e-09 0 1.8768e-09 0.0007 1.8798e-09 0 1.9938e-09 0 1.9968e-09 0.0007 1.9998e-09 0 2.1138e-09 0 2.1168e-09 0.0007 2.1198e-09 0 2.2338e-09 0 2.2368e-09 0.0007 2.2398e-09 0 2.3538e-09 0 2.3568e-09 0.0007 2.3598e-09 0 2.4738e-09 0 2.4768e-09 0.0007 2.4798e-09 0 2.5938e-09 0 2.5968e-09 0.0007 2.5998e-09 0 2.7138e-09 0 2.7168e-09 0.0007 2.7198e-09 0 2.8338e-09 0 2.8368e-09 0.0007 2.8398e-09 0 2.9538e-09 0 2.9568e-09 0.0007 2.9598e-09 0 3.0738e-09 0 3.0768e-09 0.0007 3.0798e-09 0 3.1938e-09 0 3.1968e-09 0.0007 3.1998e-09 0 3.3138e-09 0 3.3168e-09 0.0007 3.3198e-09 0 3.4338e-09 0 3.4368e-09 0.0007 3.4398e-09 0 3.5538e-09 0 3.5568e-09 0.0007 3.5598e-09 0 3.6738e-09 0 3.6768e-09 0.0007 3.6798e-09 0 3.7938e-09 0 3.7968e-09 0.0007 3.7998e-09 0 3.9138e-09 0 3.9168e-09 0.0007 3.9198e-09 0 4.0338e-09 0 4.0368e-09 0.0007 4.0398e-09 0 4.1538e-09 0 4.1568e-09 0.0007 4.1598e-09 0 4.2738e-09 0 4.2768e-09 0.0007 4.2798e-09 0 4.3938e-09 0 4.3968e-09 0.0007 4.3998e-09 0 4.5138e-09 0 4.5168e-09 0.0007 4.5198e-09 0 4.6338e-09 0 4.6368e-09 0.0007 4.6398e-09 0 4.7538e-09 0 4.7568e-09 0.0007 4.7598e-09 0 4.8738e-09 0 4.8768e-09 0.0007 4.8798e-09 0 4.9938e-09 0 4.9968e-09 0.0007 4.9998e-09 0 5.1138e-09 0 5.1168e-09 0.0007 5.1198e-09 0 5.2338e-09 0 5.2368e-09 0.0007 5.2398e-09 0 5.3538e-09 0 5.3568e-09 0.0007 5.3598e-09 0 5.4738e-09 0 5.4768e-09 0.0007 5.4798e-09 0 5.5938e-09 0 5.5968e-09 0.0007 5.5998e-09 0 5.7138e-09 0 5.7168e-09 0.0007 5.7198e-09 0 5.8338e-09 0 5.8368e-09 0.0007 5.8398e-09 0 5.9538e-09 0 5.9568e-09 0.0007 5.9598e-09 0 6.0738e-09 0 6.0768e-09 0.0007 6.0798e-09 0 6.1938e-09 0 6.1968e-09 0.0007 6.1998e-09 0 6.3138e-09 0 6.3168e-09 0.0007 6.3198e-09 0 6.4338e-09 0 6.4368e-09 0.0007 6.4398e-09 0 6.5538e-09 0 6.5568e-09 0.0007 6.5598e-09 0 6.6738e-09 0 6.6768e-09 0.0007 6.6798e-09 0 6.7938e-09 0 6.7968e-09 0.0007 6.7998e-09 0 6.9138e-09 0 6.9168e-09 0.0007 6.9198e-09 0 7.0338e-09 0 7.0368e-09 0.0007 7.0398e-09 0 7.1538e-09 0 7.1568e-09 0.0007 7.1598e-09 0 7.2738e-09 0 7.2768e-09 0.0007 7.2798e-09 0 7.3938e-09 0 7.3968e-09 0.0007 7.3998e-09 0 7.5138e-09 0 7.5168e-09 0.0007 7.5198e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 7.7538e-09 0 7.7568e-09 0.0007 7.7598e-09 0 7.8738e-09 0 7.8768e-09 0.0007 7.8798e-09 0 7.9938e-09 0 7.9968e-09 0.0007 7.9998e-09 0 8.1138e-09 0 8.1168e-09 0.0007 8.1198e-09 0 8.2338e-09 0 8.2368e-09 0.0007 8.2398e-09 0 8.3538e-09 0 8.3568e-09 0.0007 8.3598e-09 0 8.4738e-09 0 8.4768e-09 0.0007 8.4798e-09 0 8.5938e-09 0 8.5968e-09 0.0007 8.5998e-09 0 8.7138e-09 0 8.7168e-09 0.0007 8.7198e-09 0 8.8338e-09 0 8.8368e-09 0.0007 8.8398e-09 0 8.9538e-09 0 8.9568e-09 0.0007 8.9598e-09 0 9.0738e-09 0 9.0768e-09 0.0007 9.0798e-09 0 9.1938e-09 0 9.1968e-09 0.0007 9.1998e-09 0 9.3138e-09 0 9.3168e-09 0.0007 9.3198e-09 0 9.4338e-09 0 9.4368e-09 0.0007 9.4398e-09 0 9.5538e-09 0 9.5568e-09 0.0007 9.5598e-09 0 9.6738e-09 0 9.6768e-09 0.0007 9.6798e-09 0 9.7938e-09 0 9.7968e-09 0.0007 9.7998e-09 0 9.9138e-09 0 9.9168e-09 0.0007 9.9198e-09 0 1.00338e-08 0 1.00368e-08 0.0007 1.00398e-08 0 1.01538e-08 0 1.01568e-08 0.0007 1.01598e-08 0 1.02738e-08 0 1.02768e-08 0.0007 1.02798e-08 0 1.03938e-08 0 1.03968e-08 0.0007 1.03998e-08 0 1.05138e-08 0 1.05168e-08 0.0007 1.05198e-08 0 1.06338e-08 0 1.06368e-08 0.0007 1.06398e-08 0 1.07538e-08 0 1.07568e-08 0.0007 1.07598e-08 0 1.08738e-08 0 1.08768e-08 0.0007 1.08798e-08 0 1.09938e-08 0 1.09968e-08 0.0007 1.09998e-08 0 1.11138e-08 0 1.11168e-08 0.0007 1.11198e-08 0 1.12338e-08 0 1.12368e-08 0.0007 1.12398e-08 0 1.13538e-08 0 1.13568e-08 0.0007 1.13598e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.15938e-08 0 1.15968e-08 0.0007 1.15998e-08 0 1.17138e-08 0 1.17168e-08 0.0007 1.17198e-08 0 1.18338e-08 0 1.18368e-08 0.0007 1.18398e-08 0 1.19538e-08 0 1.19568e-08 0.0007 1.19598e-08 0 1.20738e-08 0 1.20768e-08 0.0007 1.20798e-08 0 1.21938e-08 0 1.21968e-08 0.0007 1.21998e-08 0 1.23138e-08 0 1.23168e-08 0.0007 1.23198e-08 0 1.24338e-08 0 1.24368e-08 0.0007 1.24398e-08 0 1.25538e-08 0 1.25568e-08 0.0007 1.25598e-08 0 1.26738e-08 0 1.26768e-08 0.0007 1.26798e-08 0 1.27938e-08 0 1.27968e-08 0.0007 1.27998e-08 0 1.29138e-08 0 1.29168e-08 0.0007 1.29198e-08 0 1.30338e-08 0 1.30368e-08 0.0007 1.30398e-08 0 1.31538e-08 0 1.31568e-08 0.0007 1.31598e-08 0 1.32738e-08 0 1.32768e-08 0.0007 1.32798e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.35138e-08 0 1.35168e-08 0.0007 1.35198e-08 0 1.36338e-08 0 1.36368e-08 0.0007 1.36398e-08 0 1.37538e-08 0 1.37568e-08 0.0007 1.37598e-08 0 1.38738e-08 0 1.38768e-08 0.0007 1.38798e-08 0 1.39938e-08 0 1.39968e-08 0.0007 1.39998e-08 0 1.41138e-08 0 1.41168e-08 0.0007 1.41198e-08 0 1.42338e-08 0 1.42368e-08 0.0007 1.42398e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.44738e-08 0 1.44768e-08 0.0007 1.44798e-08 0 1.45938e-08 0 1.45968e-08 0.0007 1.45998e-08 0 1.47138e-08 0 1.47168e-08 0.0007 1.47198e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.49538e-08 0 1.49568e-08 0.0007 1.49598e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IB0|B 0 B0_TX  PWL(0 0 1.338e-10 0 1.368e-10 0.0007 1.398e-10 0 1.938e-10 0 1.968e-10 0.0007 1.998e-10 0 3.738e-10 0 3.768e-10 0.0007 3.798e-10 0 4.338e-10 0 4.368e-10 0.0007 4.398e-10 0 6.138e-10 0 6.168e-10 0.0007 6.198e-10 0 6.738e-10 0 6.768e-10 0.0007 6.798e-10 0 8.538e-10 0 8.568e-10 0.0007 8.598e-10 0 9.138e-10 0 9.168e-10 0.0007 9.198e-10 0 1.0938e-09 0 1.0968e-09 0.0007 1.0998e-09 0 1.1538e-09 0 1.1568e-09 0.0007 1.1598e-09 0 1.3338e-09 0 1.3368e-09 0.0007 1.3398e-09 0 1.3938e-09 0 1.3968e-09 0.0007 1.3998e-09 0 1.5738e-09 0 1.5768e-09 0.0007 1.5798e-09 0 1.6338e-09 0 1.6368e-09 0.0007 1.6398e-09 0 1.8138e-09 0 1.8168e-09 0.0007 1.8198e-09 0 1.8738e-09 0 1.8768e-09 0.0007 1.8798e-09 0 2.0538e-09 0 2.0568e-09 0.0007 2.0598e-09 0 2.1138e-09 0 2.1168e-09 0.0007 2.1198e-09 0 2.2938e-09 0 2.2968e-09 0.0007 2.2998e-09 0 2.3538e-09 0 2.3568e-09 0.0007 2.3598e-09 0 2.5338e-09 0 2.5368e-09 0.0007 2.5398e-09 0 2.5938e-09 0 2.5968e-09 0.0007 2.5998e-09 0 2.7738e-09 0 2.7768e-09 0.0007 2.7798e-09 0 2.8338e-09 0 2.8368e-09 0.0007 2.8398e-09 0 3.0138e-09 0 3.0168e-09 0.0007 3.0198e-09 0 3.0738e-09 0 3.0768e-09 0.0007 3.0798e-09 0 3.2538e-09 0 3.2568e-09 0.0007 3.2598e-09 0 3.3138e-09 0 3.3168e-09 0.0007 3.3198e-09 0 3.4938e-09 0 3.4968e-09 0.0007 3.4998e-09 0 3.5538e-09 0 3.5568e-09 0.0007 3.5598e-09 0 3.7338e-09 0 3.7368e-09 0.0007 3.7398e-09 0 3.7938e-09 0 3.7968e-09 0.0007 3.7998e-09 0 3.9738e-09 0 3.9768e-09 0.0007 3.9798e-09 0 4.0338e-09 0 4.0368e-09 0.0007 4.0398e-09 0 4.2138e-09 0 4.2168e-09 0.0007 4.2198e-09 0 4.2738e-09 0 4.2768e-09 0.0007 4.2798e-09 0 4.4538e-09 0 4.4568e-09 0.0007 4.4598e-09 0 4.5138e-09 0 4.5168e-09 0.0007 4.5198e-09 0 4.6938e-09 0 4.6968e-09 0.0007 4.6998e-09 0 4.7538e-09 0 4.7568e-09 0.0007 4.7598e-09 0 4.9338e-09 0 4.9368e-09 0.0007 4.9398e-09 0 4.9938e-09 0 4.9968e-09 0.0007 4.9998e-09 0 5.1738e-09 0 5.1768e-09 0.0007 5.1798e-09 0 5.2338e-09 0 5.2368e-09 0.0007 5.2398e-09 0 5.4138e-09 0 5.4168e-09 0.0007 5.4198e-09 0 5.4738e-09 0 5.4768e-09 0.0007 5.4798e-09 0 5.6538e-09 0 5.6568e-09 0.0007 5.6598e-09 0 5.7138e-09 0 5.7168e-09 0.0007 5.7198e-09 0 5.8938e-09 0 5.8968e-09 0.0007 5.8998e-09 0 5.9538e-09 0 5.9568e-09 0.0007 5.9598e-09 0 6.1338e-09 0 6.1368e-09 0.0007 6.1398e-09 0 6.1938e-09 0 6.1968e-09 0.0007 6.1998e-09 0 6.3738e-09 0 6.3768e-09 0.0007 6.3798e-09 0 6.4338e-09 0 6.4368e-09 0.0007 6.4398e-09 0 6.6138e-09 0 6.6168e-09 0.0007 6.6198e-09 0 6.6738e-09 0 6.6768e-09 0.0007 6.6798e-09 0 6.8538e-09 0 6.8568e-09 0.0007 6.8598e-09 0 6.9138e-09 0 6.9168e-09 0.0007 6.9198e-09 0 7.0938e-09 0 7.0968e-09 0.0007 7.0998e-09 0 7.1538e-09 0 7.1568e-09 0.0007 7.1598e-09 0 7.3338e-09 0 7.3368e-09 0.0007 7.3398e-09 0 7.3938e-09 0 7.3968e-09 0.0007 7.3998e-09 0 7.5738e-09 0 7.5768e-09 0.0007 7.5798e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 7.8138e-09 0 7.8168e-09 0.0007 7.8198e-09 0 7.8738e-09 0 7.8768e-09 0.0007 7.8798e-09 0 8.0538e-09 0 8.0568e-09 0.0007 8.0598e-09 0 8.1138e-09 0 8.1168e-09 0.0007 8.1198e-09 0 8.2938e-09 0 8.2968e-09 0.0007 8.2998e-09 0 8.3538e-09 0 8.3568e-09 0.0007 8.3598e-09 0 8.5338e-09 0 8.5368e-09 0.0007 8.5398e-09 0 8.5938e-09 0 8.5968e-09 0.0007 8.5998e-09 0 8.7738e-09 0 8.7768e-09 0.0007 8.7798e-09 0 8.8338e-09 0 8.8368e-09 0.0007 8.8398e-09 0 9.0138e-09 0 9.0168e-09 0.0007 9.0198e-09 0 9.0738e-09 0 9.0768e-09 0.0007 9.0798e-09 0 9.2538e-09 0 9.2568e-09 0.0007 9.2598e-09 0 9.3138e-09 0 9.3168e-09 0.0007 9.3198e-09 0 9.4938e-09 0 9.4968e-09 0.0007 9.4998e-09 0 9.5538e-09 0 9.5568e-09 0.0007 9.5598e-09 0 9.7338e-09 0 9.7368e-09 0.0007 9.7398e-09 0 9.7938e-09 0 9.7968e-09 0.0007 9.7998e-09 0 9.9738e-09 0 9.9768e-09 0.0007 9.9798e-09 0 1.00338e-08 0 1.00368e-08 0.0007 1.00398e-08 0 1.02138e-08 0 1.02168e-08 0.0007 1.02198e-08 0 1.02738e-08 0 1.02768e-08 0.0007 1.02798e-08 0 1.04538e-08 0 1.04568e-08 0.0007 1.04598e-08 0 1.05138e-08 0 1.05168e-08 0.0007 1.05198e-08 0 1.06938e-08 0 1.06968e-08 0.0007 1.06998e-08 0 1.07538e-08 0 1.07568e-08 0.0007 1.07598e-08 0 1.09338e-08 0 1.09368e-08 0.0007 1.09398e-08 0 1.09938e-08 0 1.09968e-08 0.0007 1.09998e-08 0 1.11738e-08 0 1.11768e-08 0.0007 1.11798e-08 0 1.12338e-08 0 1.12368e-08 0.0007 1.12398e-08 0 1.14138e-08 0 1.14168e-08 0.0007 1.14198e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.16538e-08 0 1.16568e-08 0.0007 1.16598e-08 0 1.17138e-08 0 1.17168e-08 0.0007 1.17198e-08 0 1.18938e-08 0 1.18968e-08 0.0007 1.18998e-08 0 1.19538e-08 0 1.19568e-08 0.0007 1.19598e-08 0 1.21338e-08 0 1.21368e-08 0.0007 1.21398e-08 0 1.21938e-08 0 1.21968e-08 0.0007 1.21998e-08 0 1.23738e-08 0 1.23768e-08 0.0007 1.23798e-08 0 1.24338e-08 0 1.24368e-08 0.0007 1.24398e-08 0 1.26138e-08 0 1.26168e-08 0.0007 1.26198e-08 0 1.26738e-08 0 1.26768e-08 0.0007 1.26798e-08 0 1.28538e-08 0 1.28568e-08 0.0007 1.28598e-08 0 1.29138e-08 0 1.29168e-08 0.0007 1.29198e-08 0 1.30938e-08 0 1.30968e-08 0.0007 1.30998e-08 0 1.31538e-08 0 1.31568e-08 0.0007 1.31598e-08 0 1.33338e-08 0 1.33368e-08 0.0007 1.33398e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.35738e-08 0 1.35768e-08 0.0007 1.35798e-08 0 1.36338e-08 0 1.36368e-08 0.0007 1.36398e-08 0 1.38138e-08 0 1.38168e-08 0.0007 1.38198e-08 0 1.38738e-08 0 1.38768e-08 0.0007 1.38798e-08 0 1.40538e-08 0 1.40568e-08 0.0007 1.40598e-08 0 1.41138e-08 0 1.41168e-08 0.0007 1.41198e-08 0 1.42938e-08 0 1.42968e-08 0.0007 1.42998e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.45338e-08 0 1.45368e-08 0.0007 1.45398e-08 0 1.45938e-08 0 1.45968e-08 0.0007 1.45998e-08 0 1.47738e-08 0 1.47768e-08 0.0007 1.47798e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.50138e-08 0 1.50168e-08 0.0007 1.50198e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IA1|C 0 A1_TX  PWL(0 0 2.538e-10 0 2.568e-10 0.0007 2.598e-10 0 3.138e-10 0 3.168e-10 0.0007 3.198e-10 0 3.738e-10 0 3.768e-10 0.0007 3.798e-10 0 4.338e-10 0 4.368e-10 0.0007 4.398e-10 0 7.338e-10 0 7.368e-10 0.0007 7.398e-10 0 7.938e-10 0 7.968e-10 0.0007 7.998e-10 0 8.538e-10 0 8.568e-10 0.0007 8.598e-10 0 9.138e-10 0 9.168e-10 0.0007 9.198e-10 0 1.2138e-09 0 1.2168e-09 0.0007 1.2198e-09 0 1.2738e-09 0 1.2768e-09 0.0007 1.2798e-09 0 1.3338e-09 0 1.3368e-09 0.0007 1.3398e-09 0 1.3938e-09 0 1.3968e-09 0.0007 1.3998e-09 0 1.6938e-09 0 1.6968e-09 0.0007 1.6998e-09 0 1.7538e-09 0 1.7568e-09 0.0007 1.7598e-09 0 1.8138e-09 0 1.8168e-09 0.0007 1.8198e-09 0 1.8738e-09 0 1.8768e-09 0.0007 1.8798e-09 0 2.1738e-09 0 2.1768e-09 0.0007 2.1798e-09 0 2.2338e-09 0 2.2368e-09 0.0007 2.2398e-09 0 2.2938e-09 0 2.2968e-09 0.0007 2.2998e-09 0 2.3538e-09 0 2.3568e-09 0.0007 2.3598e-09 0 2.6538e-09 0 2.6568e-09 0.0007 2.6598e-09 0 2.7138e-09 0 2.7168e-09 0.0007 2.7198e-09 0 2.7738e-09 0 2.7768e-09 0.0007 2.7798e-09 0 2.8338e-09 0 2.8368e-09 0.0007 2.8398e-09 0 3.1338e-09 0 3.1368e-09 0.0007 3.1398e-09 0 3.1938e-09 0 3.1968e-09 0.0007 3.1998e-09 0 3.2538e-09 0 3.2568e-09 0.0007 3.2598e-09 0 3.3138e-09 0 3.3168e-09 0.0007 3.3198e-09 0 3.6138e-09 0 3.6168e-09 0.0007 3.6198e-09 0 3.6738e-09 0 3.6768e-09 0.0007 3.6798e-09 0 3.7338e-09 0 3.7368e-09 0.0007 3.7398e-09 0 3.7938e-09 0 3.7968e-09 0.0007 3.7998e-09 0 4.0938e-09 0 4.0968e-09 0.0007 4.0998e-09 0 4.1538e-09 0 4.1568e-09 0.0007 4.1598e-09 0 4.2138e-09 0 4.2168e-09 0.0007 4.2198e-09 0 4.2738e-09 0 4.2768e-09 0.0007 4.2798e-09 0 4.5738e-09 0 4.5768e-09 0.0007 4.5798e-09 0 4.6338e-09 0 4.6368e-09 0.0007 4.6398e-09 0 4.6938e-09 0 4.6968e-09 0.0007 4.6998e-09 0 4.7538e-09 0 4.7568e-09 0.0007 4.7598e-09 0 5.0538e-09 0 5.0568e-09 0.0007 5.0598e-09 0 5.1138e-09 0 5.1168e-09 0.0007 5.1198e-09 0 5.1738e-09 0 5.1768e-09 0.0007 5.1798e-09 0 5.2338e-09 0 5.2368e-09 0.0007 5.2398e-09 0 5.5338e-09 0 5.5368e-09 0.0007 5.5398e-09 0 5.5938e-09 0 5.5968e-09 0.0007 5.5998e-09 0 5.6538e-09 0 5.6568e-09 0.0007 5.6598e-09 0 5.7138e-09 0 5.7168e-09 0.0007 5.7198e-09 0 6.0138e-09 0 6.0168e-09 0.0007 6.0198e-09 0 6.0738e-09 0 6.0768e-09 0.0007 6.0798e-09 0 6.1338e-09 0 6.1368e-09 0.0007 6.1398e-09 0 6.1938e-09 0 6.1968e-09 0.0007 6.1998e-09 0 6.4938e-09 0 6.4968e-09 0.0007 6.4998e-09 0 6.5538e-09 0 6.5568e-09 0.0007 6.5598e-09 0 6.6138e-09 0 6.6168e-09 0.0007 6.6198e-09 0 6.6738e-09 0 6.6768e-09 0.0007 6.6798e-09 0 6.9738e-09 0 6.9768e-09 0.0007 6.9798e-09 0 7.0338e-09 0 7.0368e-09 0.0007 7.0398e-09 0 7.0938e-09 0 7.0968e-09 0.0007 7.0998e-09 0 7.1538e-09 0 7.1568e-09 0.0007 7.1598e-09 0 7.4538e-09 0 7.4568e-09 0.0007 7.4598e-09 0 7.5138e-09 0 7.5168e-09 0.0007 7.5198e-09 0 7.5738e-09 0 7.5768e-09 0.0007 7.5798e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 7.9338e-09 0 7.9368e-09 0.0007 7.9398e-09 0 7.9938e-09 0 7.9968e-09 0.0007 7.9998e-09 0 8.0538e-09 0 8.0568e-09 0.0007 8.0598e-09 0 8.1138e-09 0 8.1168e-09 0.0007 8.1198e-09 0 8.4138e-09 0 8.4168e-09 0.0007 8.4198e-09 0 8.4738e-09 0 8.4768e-09 0.0007 8.4798e-09 0 8.5338e-09 0 8.5368e-09 0.0007 8.5398e-09 0 8.5938e-09 0 8.5968e-09 0.0007 8.5998e-09 0 8.8938e-09 0 8.8968e-09 0.0007 8.8998e-09 0 8.9538e-09 0 8.9568e-09 0.0007 8.9598e-09 0 9.0138e-09 0 9.0168e-09 0.0007 9.0198e-09 0 9.0738e-09 0 9.0768e-09 0.0007 9.0798e-09 0 9.3738e-09 0 9.3768e-09 0.0007 9.3798e-09 0 9.4338e-09 0 9.4368e-09 0.0007 9.4398e-09 0 9.4938e-09 0 9.4968e-09 0.0007 9.4998e-09 0 9.5538e-09 0 9.5568e-09 0.0007 9.5598e-09 0 9.8538e-09 0 9.8568e-09 0.0007 9.8598e-09 0 9.9138e-09 0 9.9168e-09 0.0007 9.9198e-09 0 9.9738e-09 0 9.9768e-09 0.0007 9.9798e-09 0 1.00338e-08 0 1.00368e-08 0.0007 1.00398e-08 0 1.03338e-08 0 1.03368e-08 0.0007 1.03398e-08 0 1.03938e-08 0 1.03968e-08 0.0007 1.03998e-08 0 1.04538e-08 0 1.04568e-08 0.0007 1.04598e-08 0 1.05138e-08 0 1.05168e-08 0.0007 1.05198e-08 0 1.08138e-08 0 1.08168e-08 0.0007 1.08198e-08 0 1.08738e-08 0 1.08768e-08 0.0007 1.08798e-08 0 1.09338e-08 0 1.09368e-08 0.0007 1.09398e-08 0 1.09938e-08 0 1.09968e-08 0.0007 1.09998e-08 0 1.12938e-08 0 1.12968e-08 0.0007 1.12998e-08 0 1.13538e-08 0 1.13568e-08 0.0007 1.13598e-08 0 1.14138e-08 0 1.14168e-08 0.0007 1.14198e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.17738e-08 0 1.17768e-08 0.0007 1.17798e-08 0 1.18338e-08 0 1.18368e-08 0.0007 1.18398e-08 0 1.18938e-08 0 1.18968e-08 0.0007 1.18998e-08 0 1.19538e-08 0 1.19568e-08 0.0007 1.19598e-08 0 1.22538e-08 0 1.22568e-08 0.0007 1.22598e-08 0 1.23138e-08 0 1.23168e-08 0.0007 1.23198e-08 0 1.23738e-08 0 1.23768e-08 0.0007 1.23798e-08 0 1.24338e-08 0 1.24368e-08 0.0007 1.24398e-08 0 1.27338e-08 0 1.27368e-08 0.0007 1.27398e-08 0 1.27938e-08 0 1.27968e-08 0.0007 1.27998e-08 0 1.28538e-08 0 1.28568e-08 0.0007 1.28598e-08 0 1.29138e-08 0 1.29168e-08 0.0007 1.29198e-08 0 1.32138e-08 0 1.32168e-08 0.0007 1.32198e-08 0 1.32738e-08 0 1.32768e-08 0.0007 1.32798e-08 0 1.33338e-08 0 1.33368e-08 0.0007 1.33398e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.36938e-08 0 1.36968e-08 0.0007 1.36998e-08 0 1.37538e-08 0 1.37568e-08 0.0007 1.37598e-08 0 1.38138e-08 0 1.38168e-08 0.0007 1.38198e-08 0 1.38738e-08 0 1.38768e-08 0.0007 1.38798e-08 0 1.41738e-08 0 1.41768e-08 0.0007 1.41798e-08 0 1.42338e-08 0 1.42368e-08 0.0007 1.42398e-08 0 1.42938e-08 0 1.42968e-08 0.0007 1.42998e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.46538e-08 0 1.46568e-08 0.0007 1.46598e-08 0 1.47138e-08 0 1.47168e-08 0.0007 1.47198e-08 0 1.47738e-08 0 1.47768e-08 0.0007 1.47798e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.51338e-08 0 1.51368e-08 0.0007 1.51398e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IB1|D 0 B1_TX  PWL(0 0 4.938e-10 0 4.968e-10 0.0007 4.998e-10 0 5.538e-10 0 5.568e-10 0.0007 5.598e-10 0 6.138e-10 0 6.168e-10 0.0007 6.198e-10 0 6.738e-10 0 6.768e-10 0.0007 6.798e-10 0 7.338e-10 0 7.368e-10 0.0007 7.398e-10 0 7.938e-10 0 7.968e-10 0.0007 7.998e-10 0 8.538e-10 0 8.568e-10 0.0007 8.598e-10 0 9.138e-10 0 9.168e-10 0.0007 9.198e-10 0 1.4538e-09 0 1.4568e-09 0.0007 1.4598e-09 0 1.5138e-09 0 1.5168e-09 0.0007 1.5198e-09 0 1.5738e-09 0 1.5768e-09 0.0007 1.5798e-09 0 1.6338e-09 0 1.6368e-09 0.0007 1.6398e-09 0 1.6938e-09 0 1.6968e-09 0.0007 1.6998e-09 0 1.7538e-09 0 1.7568e-09 0.0007 1.7598e-09 0 1.8138e-09 0 1.8168e-09 0.0007 1.8198e-09 0 1.8738e-09 0 1.8768e-09 0.0007 1.8798e-09 0 2.4138e-09 0 2.4168e-09 0.0007 2.4198e-09 0 2.4738e-09 0 2.4768e-09 0.0007 2.4798e-09 0 2.5338e-09 0 2.5368e-09 0.0007 2.5398e-09 0 2.5938e-09 0 2.5968e-09 0.0007 2.5998e-09 0 2.6538e-09 0 2.6568e-09 0.0007 2.6598e-09 0 2.7138e-09 0 2.7168e-09 0.0007 2.7198e-09 0 2.7738e-09 0 2.7768e-09 0.0007 2.7798e-09 0 2.8338e-09 0 2.8368e-09 0.0007 2.8398e-09 0 3.3738e-09 0 3.3768e-09 0.0007 3.3798e-09 0 3.4338e-09 0 3.4368e-09 0.0007 3.4398e-09 0 3.4938e-09 0 3.4968e-09 0.0007 3.4998e-09 0 3.5538e-09 0 3.5568e-09 0.0007 3.5598e-09 0 3.6138e-09 0 3.6168e-09 0.0007 3.6198e-09 0 3.6738e-09 0 3.6768e-09 0.0007 3.6798e-09 0 3.7338e-09 0 3.7368e-09 0.0007 3.7398e-09 0 3.7938e-09 0 3.7968e-09 0.0007 3.7998e-09 0 4.3338e-09 0 4.3368e-09 0.0007 4.3398e-09 0 4.3938e-09 0 4.3968e-09 0.0007 4.3998e-09 0 4.4538e-09 0 4.4568e-09 0.0007 4.4598e-09 0 4.5138e-09 0 4.5168e-09 0.0007 4.5198e-09 0 4.5738e-09 0 4.5768e-09 0.0007 4.5798e-09 0 4.6338e-09 0 4.6368e-09 0.0007 4.6398e-09 0 4.6938e-09 0 4.6968e-09 0.0007 4.6998e-09 0 4.7538e-09 0 4.7568e-09 0.0007 4.7598e-09 0 5.2938e-09 0 5.2968e-09 0.0007 5.2998e-09 0 5.3538e-09 0 5.3568e-09 0.0007 5.3598e-09 0 5.4138e-09 0 5.4168e-09 0.0007 5.4198e-09 0 5.4738e-09 0 5.4768e-09 0.0007 5.4798e-09 0 5.5338e-09 0 5.5368e-09 0.0007 5.5398e-09 0 5.5938e-09 0 5.5968e-09 0.0007 5.5998e-09 0 5.6538e-09 0 5.6568e-09 0.0007 5.6598e-09 0 5.7138e-09 0 5.7168e-09 0.0007 5.7198e-09 0 6.2538e-09 0 6.2568e-09 0.0007 6.2598e-09 0 6.3138e-09 0 6.3168e-09 0.0007 6.3198e-09 0 6.3738e-09 0 6.3768e-09 0.0007 6.3798e-09 0 6.4338e-09 0 6.4368e-09 0.0007 6.4398e-09 0 6.4938e-09 0 6.4968e-09 0.0007 6.4998e-09 0 6.5538e-09 0 6.5568e-09 0.0007 6.5598e-09 0 6.6138e-09 0 6.6168e-09 0.0007 6.6198e-09 0 6.6738e-09 0 6.6768e-09 0.0007 6.6798e-09 0 7.2138e-09 0 7.2168e-09 0.0007 7.2198e-09 0 7.2738e-09 0 7.2768e-09 0.0007 7.2798e-09 0 7.3338e-09 0 7.3368e-09 0.0007 7.3398e-09 0 7.3938e-09 0 7.3968e-09 0.0007 7.3998e-09 0 7.4538e-09 0 7.4568e-09 0.0007 7.4598e-09 0 7.5138e-09 0 7.5168e-09 0.0007 7.5198e-09 0 7.5738e-09 0 7.5768e-09 0.0007 7.5798e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 8.1738e-09 0 8.1768e-09 0.0007 8.1798e-09 0 8.2338e-09 0 8.2368e-09 0.0007 8.2398e-09 0 8.2938e-09 0 8.2968e-09 0.0007 8.2998e-09 0 8.3538e-09 0 8.3568e-09 0.0007 8.3598e-09 0 8.4138e-09 0 8.4168e-09 0.0007 8.4198e-09 0 8.4738e-09 0 8.4768e-09 0.0007 8.4798e-09 0 8.5338e-09 0 8.5368e-09 0.0007 8.5398e-09 0 8.5938e-09 0 8.5968e-09 0.0007 8.5998e-09 0 9.1338e-09 0 9.1368e-09 0.0007 9.1398e-09 0 9.1938e-09 0 9.1968e-09 0.0007 9.1998e-09 0 9.2538e-09 0 9.2568e-09 0.0007 9.2598e-09 0 9.3138e-09 0 9.3168e-09 0.0007 9.3198e-09 0 9.3738e-09 0 9.3768e-09 0.0007 9.3798e-09 0 9.4338e-09 0 9.4368e-09 0.0007 9.4398e-09 0 9.4938e-09 0 9.4968e-09 0.0007 9.4998e-09 0 9.5538e-09 0 9.5568e-09 0.0007 9.5598e-09 0 1.00938e-08 0 1.00968e-08 0.0007 1.00998e-08 0 1.01538e-08 0 1.01568e-08 0.0007 1.01598e-08 0 1.02138e-08 0 1.02168e-08 0.0007 1.02198e-08 0 1.02738e-08 0 1.02768e-08 0.0007 1.02798e-08 0 1.03338e-08 0 1.03368e-08 0.0007 1.03398e-08 0 1.03938e-08 0 1.03968e-08 0.0007 1.03998e-08 0 1.04538e-08 0 1.04568e-08 0.0007 1.04598e-08 0 1.05138e-08 0 1.05168e-08 0.0007 1.05198e-08 0 1.10538e-08 0 1.10568e-08 0.0007 1.10598e-08 0 1.11138e-08 0 1.11168e-08 0.0007 1.11198e-08 0 1.11738e-08 0 1.11768e-08 0.0007 1.11798e-08 0 1.12338e-08 0 1.12368e-08 0.0007 1.12398e-08 0 1.12938e-08 0 1.12968e-08 0.0007 1.12998e-08 0 1.13538e-08 0 1.13568e-08 0.0007 1.13598e-08 0 1.14138e-08 0 1.14168e-08 0.0007 1.14198e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.20138e-08 0 1.20168e-08 0.0007 1.20198e-08 0 1.20738e-08 0 1.20768e-08 0.0007 1.20798e-08 0 1.21338e-08 0 1.21368e-08 0.0007 1.21398e-08 0 1.21938e-08 0 1.21968e-08 0.0007 1.21998e-08 0 1.22538e-08 0 1.22568e-08 0.0007 1.22598e-08 0 1.23138e-08 0 1.23168e-08 0.0007 1.23198e-08 0 1.23738e-08 0 1.23768e-08 0.0007 1.23798e-08 0 1.24338e-08 0 1.24368e-08 0.0007 1.24398e-08 0 1.29738e-08 0 1.29768e-08 0.0007 1.29798e-08 0 1.30338e-08 0 1.30368e-08 0.0007 1.30398e-08 0 1.30938e-08 0 1.30968e-08 0.0007 1.30998e-08 0 1.31538e-08 0 1.31568e-08 0.0007 1.31598e-08 0 1.32138e-08 0 1.32168e-08 0.0007 1.32198e-08 0 1.32738e-08 0 1.32768e-08 0.0007 1.32798e-08 0 1.33338e-08 0 1.33368e-08 0.0007 1.33398e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.39338e-08 0 1.39368e-08 0.0007 1.39398e-08 0 1.39938e-08 0 1.39968e-08 0.0007 1.39998e-08 0 1.40538e-08 0 1.40568e-08 0.0007 1.40598e-08 0 1.41138e-08 0 1.41168e-08 0.0007 1.41198e-08 0 1.41738e-08 0 1.41768e-08 0.0007 1.41798e-08 0 1.42338e-08 0 1.42368e-08 0.0007 1.42398e-08 0 1.42938e-08 0 1.42968e-08 0.0007 1.42998e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.48938e-08 0 1.48968e-08 0.0007 1.48998e-08 0 1.49538e-08 0 1.49568e-08 0.0007 1.49598e-08 0 1.50138e-08 0 1.50168e-08 0.0007 1.50198e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.51338e-08 0 1.51368e-08 0.0007 1.51398e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IA2|E 0 A2_TX  PWL(0 0 9.738e-10 0 9.768e-10 0.0007 9.798e-10 0 1.0338e-09 0 1.0368e-09 0.0007 1.0398e-09 0 1.0938e-09 0 1.0968e-09 0.0007 1.0998e-09 0 1.1538e-09 0 1.1568e-09 0.0007 1.1598e-09 0 1.2138e-09 0 1.2168e-09 0.0007 1.2198e-09 0 1.2738e-09 0 1.2768e-09 0.0007 1.2798e-09 0 1.3338e-09 0 1.3368e-09 0.0007 1.3398e-09 0 1.3938e-09 0 1.3968e-09 0.0007 1.3998e-09 0 1.4538e-09 0 1.4568e-09 0.0007 1.4598e-09 0 1.5138e-09 0 1.5168e-09 0.0007 1.5198e-09 0 1.5738e-09 0 1.5768e-09 0.0007 1.5798e-09 0 1.6338e-09 0 1.6368e-09 0.0007 1.6398e-09 0 1.6938e-09 0 1.6968e-09 0.0007 1.6998e-09 0 1.7538e-09 0 1.7568e-09 0.0007 1.7598e-09 0 1.8138e-09 0 1.8168e-09 0.0007 1.8198e-09 0 1.8738e-09 0 1.8768e-09 0.0007 1.8798e-09 0 2.8938e-09 0 2.8968e-09 0.0007 2.8998e-09 0 2.9538e-09 0 2.9568e-09 0.0007 2.9598e-09 0 3.0138e-09 0 3.0168e-09 0.0007 3.0198e-09 0 3.0738e-09 0 3.0768e-09 0.0007 3.0798e-09 0 3.1338e-09 0 3.1368e-09 0.0007 3.1398e-09 0 3.1938e-09 0 3.1968e-09 0.0007 3.1998e-09 0 3.2538e-09 0 3.2568e-09 0.0007 3.2598e-09 0 3.3138e-09 0 3.3168e-09 0.0007 3.3198e-09 0 3.3738e-09 0 3.3768e-09 0.0007 3.3798e-09 0 3.4338e-09 0 3.4368e-09 0.0007 3.4398e-09 0 3.4938e-09 0 3.4968e-09 0.0007 3.4998e-09 0 3.5538e-09 0 3.5568e-09 0.0007 3.5598e-09 0 3.6138e-09 0 3.6168e-09 0.0007 3.6198e-09 0 3.6738e-09 0 3.6768e-09 0.0007 3.6798e-09 0 3.7338e-09 0 3.7368e-09 0.0007 3.7398e-09 0 3.7938e-09 0 3.7968e-09 0.0007 3.7998e-09 0 4.8138e-09 0 4.8168e-09 0.0007 4.8198e-09 0 4.8738e-09 0 4.8768e-09 0.0007 4.8798e-09 0 4.9338e-09 0 4.9368e-09 0.0007 4.9398e-09 0 4.9938e-09 0 4.9968e-09 0.0007 4.9998e-09 0 5.0538e-09 0 5.0568e-09 0.0007 5.0598e-09 0 5.1138e-09 0 5.1168e-09 0.0007 5.1198e-09 0 5.1738e-09 0 5.1768e-09 0.0007 5.1798e-09 0 5.2338e-09 0 5.2368e-09 0.0007 5.2398e-09 0 5.2938e-09 0 5.2968e-09 0.0007 5.2998e-09 0 5.3538e-09 0 5.3568e-09 0.0007 5.3598e-09 0 5.4138e-09 0 5.4168e-09 0.0007 5.4198e-09 0 5.4738e-09 0 5.4768e-09 0.0007 5.4798e-09 0 5.5338e-09 0 5.5368e-09 0.0007 5.5398e-09 0 5.5938e-09 0 5.5968e-09 0.0007 5.5998e-09 0 5.6538e-09 0 5.6568e-09 0.0007 5.6598e-09 0 5.7138e-09 0 5.7168e-09 0.0007 5.7198e-09 0 6.7338e-09 0 6.7368e-09 0.0007 6.7398e-09 0 6.7938e-09 0 6.7968e-09 0.0007 6.7998e-09 0 6.8538e-09 0 6.8568e-09 0.0007 6.8598e-09 0 6.9138e-09 0 6.9168e-09 0.0007 6.9198e-09 0 6.9738e-09 0 6.9768e-09 0.0007 6.9798e-09 0 7.0338e-09 0 7.0368e-09 0.0007 7.0398e-09 0 7.0938e-09 0 7.0968e-09 0.0007 7.0998e-09 0 7.1538e-09 0 7.1568e-09 0.0007 7.1598e-09 0 7.2138e-09 0 7.2168e-09 0.0007 7.2198e-09 0 7.2738e-09 0 7.2768e-09 0.0007 7.2798e-09 0 7.3338e-09 0 7.3368e-09 0.0007 7.3398e-09 0 7.3938e-09 0 7.3968e-09 0.0007 7.3998e-09 0 7.4538e-09 0 7.4568e-09 0.0007 7.4598e-09 0 7.5138e-09 0 7.5168e-09 0.0007 7.5198e-09 0 7.5738e-09 0 7.5768e-09 0.0007 7.5798e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 8.6538e-09 0 8.6568e-09 0.0007 8.6598e-09 0 8.7138e-09 0 8.7168e-09 0.0007 8.7198e-09 0 8.7738e-09 0 8.7768e-09 0.0007 8.7798e-09 0 8.8338e-09 0 8.8368e-09 0.0007 8.8398e-09 0 8.8938e-09 0 8.8968e-09 0.0007 8.8998e-09 0 8.9538e-09 0 8.9568e-09 0.0007 8.9598e-09 0 9.0138e-09 0 9.0168e-09 0.0007 9.0198e-09 0 9.0738e-09 0 9.0768e-09 0.0007 9.0798e-09 0 9.1338e-09 0 9.1368e-09 0.0007 9.1398e-09 0 9.1938e-09 0 9.1968e-09 0.0007 9.1998e-09 0 9.2538e-09 0 9.2568e-09 0.0007 9.2598e-09 0 9.3138e-09 0 9.3168e-09 0.0007 9.3198e-09 0 9.3738e-09 0 9.3768e-09 0.0007 9.3798e-09 0 9.4338e-09 0 9.4368e-09 0.0007 9.4398e-09 0 9.4938e-09 0 9.4968e-09 0.0007 9.4998e-09 0 9.5538e-09 0 9.5568e-09 0.0007 9.5598e-09 0 1.05738e-08 0 1.05768e-08 0.0007 1.05798e-08 0 1.06338e-08 0 1.06368e-08 0.0007 1.06398e-08 0 1.06938e-08 0 1.06968e-08 0.0007 1.06998e-08 0 1.07538e-08 0 1.07568e-08 0.0007 1.07598e-08 0 1.08138e-08 0 1.08168e-08 0.0007 1.08198e-08 0 1.08738e-08 0 1.08768e-08 0.0007 1.08798e-08 0 1.09338e-08 0 1.09368e-08 0.0007 1.09398e-08 0 1.09938e-08 0 1.09968e-08 0.0007 1.09998e-08 0 1.10538e-08 0 1.10568e-08 0.0007 1.10598e-08 0 1.11138e-08 0 1.11168e-08 0.0007 1.11198e-08 0 1.11738e-08 0 1.11768e-08 0.0007 1.11798e-08 0 1.12338e-08 0 1.12368e-08 0.0007 1.12398e-08 0 1.12938e-08 0 1.12968e-08 0.0007 1.12998e-08 0 1.13538e-08 0 1.13568e-08 0.0007 1.13598e-08 0 1.14138e-08 0 1.14168e-08 0.0007 1.14198e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.24938e-08 0 1.24968e-08 0.0007 1.24998e-08 0 1.25538e-08 0 1.25568e-08 0.0007 1.25598e-08 0 1.26138e-08 0 1.26168e-08 0.0007 1.26198e-08 0 1.26738e-08 0 1.26768e-08 0.0007 1.26798e-08 0 1.27338e-08 0 1.27368e-08 0.0007 1.27398e-08 0 1.27938e-08 0 1.27968e-08 0.0007 1.27998e-08 0 1.28538e-08 0 1.28568e-08 0.0007 1.28598e-08 0 1.29138e-08 0 1.29168e-08 0.0007 1.29198e-08 0 1.29738e-08 0 1.29768e-08 0.0007 1.29798e-08 0 1.30338e-08 0 1.30368e-08 0.0007 1.30398e-08 0 1.30938e-08 0 1.30968e-08 0.0007 1.30998e-08 0 1.31538e-08 0 1.31568e-08 0.0007 1.31598e-08 0 1.32138e-08 0 1.32168e-08 0.0007 1.32198e-08 0 1.32738e-08 0 1.32768e-08 0.0007 1.32798e-08 0 1.33338e-08 0 1.33368e-08 0.0007 1.33398e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.44138e-08 0 1.44168e-08 0.0007 1.44198e-08 0 1.44738e-08 0 1.44768e-08 0.0007 1.44798e-08 0 1.45338e-08 0 1.45368e-08 0.0007 1.45398e-08 0 1.45938e-08 0 1.45968e-08 0.0007 1.45998e-08 0 1.46538e-08 0 1.46568e-08 0.0007 1.46598e-08 0 1.47138e-08 0 1.47168e-08 0.0007 1.47198e-08 0 1.47738e-08 0 1.47768e-08 0.0007 1.47798e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.48938e-08 0 1.48968e-08 0.0007 1.48998e-08 0 1.49538e-08 0 1.49568e-08 0.0007 1.49598e-08 0 1.50138e-08 0 1.50168e-08 0.0007 1.50198e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.51338e-08 0 1.51368e-08 0.0007 1.51398e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IB2|F 0 B2_TX  PWL(0 0 1.9338e-09 0 1.9368e-09 0.0007 1.9398e-09 0 1.9938e-09 0 1.9968e-09 0.0007 1.9998e-09 0 2.0538e-09 0 2.0568e-09 0.0007 2.0598e-09 0 2.1138e-09 0 2.1168e-09 0.0007 2.1198e-09 0 2.1738e-09 0 2.1768e-09 0.0007 2.1798e-09 0 2.2338e-09 0 2.2368e-09 0.0007 2.2398e-09 0 2.2938e-09 0 2.2968e-09 0.0007 2.2998e-09 0 2.3538e-09 0 2.3568e-09 0.0007 2.3598e-09 0 2.4138e-09 0 2.4168e-09 0.0007 2.4198e-09 0 2.4738e-09 0 2.4768e-09 0.0007 2.4798e-09 0 2.5338e-09 0 2.5368e-09 0.0007 2.5398e-09 0 2.5938e-09 0 2.5968e-09 0.0007 2.5998e-09 0 2.6538e-09 0 2.6568e-09 0.0007 2.6598e-09 0 2.7138e-09 0 2.7168e-09 0.0007 2.7198e-09 0 2.7738e-09 0 2.7768e-09 0.0007 2.7798e-09 0 2.8338e-09 0 2.8368e-09 0.0007 2.8398e-09 0 2.8938e-09 0 2.8968e-09 0.0007 2.8998e-09 0 2.9538e-09 0 2.9568e-09 0.0007 2.9598e-09 0 3.0138e-09 0 3.0168e-09 0.0007 3.0198e-09 0 3.0738e-09 0 3.0768e-09 0.0007 3.0798e-09 0 3.1338e-09 0 3.1368e-09 0.0007 3.1398e-09 0 3.1938e-09 0 3.1968e-09 0.0007 3.1998e-09 0 3.2538e-09 0 3.2568e-09 0.0007 3.2598e-09 0 3.3138e-09 0 3.3168e-09 0.0007 3.3198e-09 0 3.3738e-09 0 3.3768e-09 0.0007 3.3798e-09 0 3.4338e-09 0 3.4368e-09 0.0007 3.4398e-09 0 3.4938e-09 0 3.4968e-09 0.0007 3.4998e-09 0 3.5538e-09 0 3.5568e-09 0.0007 3.5598e-09 0 3.6138e-09 0 3.6168e-09 0.0007 3.6198e-09 0 3.6738e-09 0 3.6768e-09 0.0007 3.6798e-09 0 3.7338e-09 0 3.7368e-09 0.0007 3.7398e-09 0 3.7938e-09 0 3.7968e-09 0.0007 3.7998e-09 0 5.7738e-09 0 5.7768e-09 0.0007 5.7798e-09 0 5.8338e-09 0 5.8368e-09 0.0007 5.8398e-09 0 5.8938e-09 0 5.8968e-09 0.0007 5.8998e-09 0 5.9538e-09 0 5.9568e-09 0.0007 5.9598e-09 0 6.0138e-09 0 6.0168e-09 0.0007 6.0198e-09 0 6.0738e-09 0 6.0768e-09 0.0007 6.0798e-09 0 6.1338e-09 0 6.1368e-09 0.0007 6.1398e-09 0 6.1938e-09 0 6.1968e-09 0.0007 6.1998e-09 0 6.2538e-09 0 6.2568e-09 0.0007 6.2598e-09 0 6.3138e-09 0 6.3168e-09 0.0007 6.3198e-09 0 6.3738e-09 0 6.3768e-09 0.0007 6.3798e-09 0 6.4338e-09 0 6.4368e-09 0.0007 6.4398e-09 0 6.4938e-09 0 6.4968e-09 0.0007 6.4998e-09 0 6.5538e-09 0 6.5568e-09 0.0007 6.5598e-09 0 6.6138e-09 0 6.6168e-09 0.0007 6.6198e-09 0 6.6738e-09 0 6.6768e-09 0.0007 6.6798e-09 0 6.7338e-09 0 6.7368e-09 0.0007 6.7398e-09 0 6.7938e-09 0 6.7968e-09 0.0007 6.7998e-09 0 6.8538e-09 0 6.8568e-09 0.0007 6.8598e-09 0 6.9138e-09 0 6.9168e-09 0.0007 6.9198e-09 0 6.9738e-09 0 6.9768e-09 0.0007 6.9798e-09 0 7.0338e-09 0 7.0368e-09 0.0007 7.0398e-09 0 7.0938e-09 0 7.0968e-09 0.0007 7.0998e-09 0 7.1538e-09 0 7.1568e-09 0.0007 7.1598e-09 0 7.2138e-09 0 7.2168e-09 0.0007 7.2198e-09 0 7.2738e-09 0 7.2768e-09 0.0007 7.2798e-09 0 7.3338e-09 0 7.3368e-09 0.0007 7.3398e-09 0 7.3938e-09 0 7.3968e-09 0.0007 7.3998e-09 0 7.4538e-09 0 7.4568e-09 0.0007 7.4598e-09 0 7.5138e-09 0 7.5168e-09 0.0007 7.5198e-09 0 7.5738e-09 0 7.5768e-09 0.0007 7.5798e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 9.6138e-09 0 9.6168e-09 0.0007 9.6198e-09 0 9.6738e-09 0 9.6768e-09 0.0007 9.6798e-09 0 9.7338e-09 0 9.7368e-09 0.0007 9.7398e-09 0 9.7938e-09 0 9.7968e-09 0.0007 9.7998e-09 0 9.8538e-09 0 9.8568e-09 0.0007 9.8598e-09 0 9.9138e-09 0 9.9168e-09 0.0007 9.9198e-09 0 9.9738e-09 0 9.9768e-09 0.0007 9.9798e-09 0 1.00338e-08 0 1.00368e-08 0.0007 1.00398e-08 0 1.00938e-08 0 1.00968e-08 0.0007 1.00998e-08 0 1.01538e-08 0 1.01568e-08 0.0007 1.01598e-08 0 1.02138e-08 0 1.02168e-08 0.0007 1.02198e-08 0 1.02738e-08 0 1.02768e-08 0.0007 1.02798e-08 0 1.03338e-08 0 1.03368e-08 0.0007 1.03398e-08 0 1.03938e-08 0 1.03968e-08 0.0007 1.03998e-08 0 1.04538e-08 0 1.04568e-08 0.0007 1.04598e-08 0 1.05138e-08 0 1.05168e-08 0.0007 1.05198e-08 0 1.05738e-08 0 1.05768e-08 0.0007 1.05798e-08 0 1.06338e-08 0 1.06368e-08 0.0007 1.06398e-08 0 1.06938e-08 0 1.06968e-08 0.0007 1.06998e-08 0 1.07538e-08 0 1.07568e-08 0.0007 1.07598e-08 0 1.08138e-08 0 1.08168e-08 0.0007 1.08198e-08 0 1.08738e-08 0 1.08768e-08 0.0007 1.08798e-08 0 1.09338e-08 0 1.09368e-08 0.0007 1.09398e-08 0 1.09938e-08 0 1.09968e-08 0.0007 1.09998e-08 0 1.10538e-08 0 1.10568e-08 0.0007 1.10598e-08 0 1.11138e-08 0 1.11168e-08 0.0007 1.11198e-08 0 1.11738e-08 0 1.11768e-08 0.0007 1.11798e-08 0 1.12338e-08 0 1.12368e-08 0.0007 1.12398e-08 0 1.12938e-08 0 1.12968e-08 0.0007 1.12998e-08 0 1.13538e-08 0 1.13568e-08 0.0007 1.13598e-08 0 1.14138e-08 0 1.14168e-08 0.0007 1.14198e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.34538e-08 0 1.34568e-08 0.0007 1.34598e-08 0 1.35138e-08 0 1.35168e-08 0.0007 1.35198e-08 0 1.35738e-08 0 1.35768e-08 0.0007 1.35798e-08 0 1.36338e-08 0 1.36368e-08 0.0007 1.36398e-08 0 1.36938e-08 0 1.36968e-08 0.0007 1.36998e-08 0 1.37538e-08 0 1.37568e-08 0.0007 1.37598e-08 0 1.38138e-08 0 1.38168e-08 0.0007 1.38198e-08 0 1.38738e-08 0 1.38768e-08 0.0007 1.38798e-08 0 1.39338e-08 0 1.39368e-08 0.0007 1.39398e-08 0 1.39938e-08 0 1.39968e-08 0.0007 1.39998e-08 0 1.40538e-08 0 1.40568e-08 0.0007 1.40598e-08 0 1.41138e-08 0 1.41168e-08 0.0007 1.41198e-08 0 1.41738e-08 0 1.41768e-08 0.0007 1.41798e-08 0 1.42338e-08 0 1.42368e-08 0.0007 1.42398e-08 0 1.42938e-08 0 1.42968e-08 0.0007 1.42998e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.44138e-08 0 1.44168e-08 0.0007 1.44198e-08 0 1.44738e-08 0 1.44768e-08 0.0007 1.44798e-08 0 1.45338e-08 0 1.45368e-08 0.0007 1.45398e-08 0 1.45938e-08 0 1.45968e-08 0.0007 1.45998e-08 0 1.46538e-08 0 1.46568e-08 0.0007 1.46598e-08 0 1.47138e-08 0 1.47168e-08 0.0007 1.47198e-08 0 1.47738e-08 0 1.47768e-08 0.0007 1.47798e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.48938e-08 0 1.48968e-08 0.0007 1.48998e-08 0 1.49538e-08 0 1.49568e-08 0.0007 1.49598e-08 0 1.50138e-08 0 1.50168e-08 0.0007 1.50198e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.51338e-08 0 1.51368e-08 0.0007 1.51398e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IA3|G 0 A3_TX  PWL(0 0 3.8538e-09 0 3.8568e-09 0.0007 3.8598e-09 0 3.9138e-09 0 3.9168e-09 0.0007 3.9198e-09 0 3.9738e-09 0 3.9768e-09 0.0007 3.9798e-09 0 4.0338e-09 0 4.0368e-09 0.0007 4.0398e-09 0 4.0938e-09 0 4.0968e-09 0.0007 4.0998e-09 0 4.1538e-09 0 4.1568e-09 0.0007 4.1598e-09 0 4.2138e-09 0 4.2168e-09 0.0007 4.2198e-09 0 4.2738e-09 0 4.2768e-09 0.0007 4.2798e-09 0 4.3338e-09 0 4.3368e-09 0.0007 4.3398e-09 0 4.3938e-09 0 4.3968e-09 0.0007 4.3998e-09 0 4.4538e-09 0 4.4568e-09 0.0007 4.4598e-09 0 4.5138e-09 0 4.5168e-09 0.0007 4.5198e-09 0 4.5738e-09 0 4.5768e-09 0.0007 4.5798e-09 0 4.6338e-09 0 4.6368e-09 0.0007 4.6398e-09 0 4.6938e-09 0 4.6968e-09 0.0007 4.6998e-09 0 4.7538e-09 0 4.7568e-09 0.0007 4.7598e-09 0 4.8138e-09 0 4.8168e-09 0.0007 4.8198e-09 0 4.8738e-09 0 4.8768e-09 0.0007 4.8798e-09 0 4.9338e-09 0 4.9368e-09 0.0007 4.9398e-09 0 4.9938e-09 0 4.9968e-09 0.0007 4.9998e-09 0 5.0538e-09 0 5.0568e-09 0.0007 5.0598e-09 0 5.1138e-09 0 5.1168e-09 0.0007 5.1198e-09 0 5.1738e-09 0 5.1768e-09 0.0007 5.1798e-09 0 5.2338e-09 0 5.2368e-09 0.0007 5.2398e-09 0 5.2938e-09 0 5.2968e-09 0.0007 5.2998e-09 0 5.3538e-09 0 5.3568e-09 0.0007 5.3598e-09 0 5.4138e-09 0 5.4168e-09 0.0007 5.4198e-09 0 5.4738e-09 0 5.4768e-09 0.0007 5.4798e-09 0 5.5338e-09 0 5.5368e-09 0.0007 5.5398e-09 0 5.5938e-09 0 5.5968e-09 0.0007 5.5998e-09 0 5.6538e-09 0 5.6568e-09 0.0007 5.6598e-09 0 5.7138e-09 0 5.7168e-09 0.0007 5.7198e-09 0 5.7738e-09 0 5.7768e-09 0.0007 5.7798e-09 0 5.8338e-09 0 5.8368e-09 0.0007 5.8398e-09 0 5.8938e-09 0 5.8968e-09 0.0007 5.8998e-09 0 5.9538e-09 0 5.9568e-09 0.0007 5.9598e-09 0 6.0138e-09 0 6.0168e-09 0.0007 6.0198e-09 0 6.0738e-09 0 6.0768e-09 0.0007 6.0798e-09 0 6.1338e-09 0 6.1368e-09 0.0007 6.1398e-09 0 6.1938e-09 0 6.1968e-09 0.0007 6.1998e-09 0 6.2538e-09 0 6.2568e-09 0.0007 6.2598e-09 0 6.3138e-09 0 6.3168e-09 0.0007 6.3198e-09 0 6.3738e-09 0 6.3768e-09 0.0007 6.3798e-09 0 6.4338e-09 0 6.4368e-09 0.0007 6.4398e-09 0 6.4938e-09 0 6.4968e-09 0.0007 6.4998e-09 0 6.5538e-09 0 6.5568e-09 0.0007 6.5598e-09 0 6.6138e-09 0 6.6168e-09 0.0007 6.6198e-09 0 6.6738e-09 0 6.6768e-09 0.0007 6.6798e-09 0 6.7338e-09 0 6.7368e-09 0.0007 6.7398e-09 0 6.7938e-09 0 6.7968e-09 0.0007 6.7998e-09 0 6.8538e-09 0 6.8568e-09 0.0007 6.8598e-09 0 6.9138e-09 0 6.9168e-09 0.0007 6.9198e-09 0 6.9738e-09 0 6.9768e-09 0.0007 6.9798e-09 0 7.0338e-09 0 7.0368e-09 0.0007 7.0398e-09 0 7.0938e-09 0 7.0968e-09 0.0007 7.0998e-09 0 7.1538e-09 0 7.1568e-09 0.0007 7.1598e-09 0 7.2138e-09 0 7.2168e-09 0.0007 7.2198e-09 0 7.2738e-09 0 7.2768e-09 0.0007 7.2798e-09 0 7.3338e-09 0 7.3368e-09 0.0007 7.3398e-09 0 7.3938e-09 0 7.3968e-09 0.0007 7.3998e-09 0 7.4538e-09 0 7.4568e-09 0.0007 7.4598e-09 0 7.5138e-09 0 7.5168e-09 0.0007 7.5198e-09 0 7.5738e-09 0 7.5768e-09 0.0007 7.5798e-09 0 7.6338e-09 0 7.6368e-09 0.0007 7.6398e-09 0 1.15338e-08 0 1.15368e-08 0.0007 1.15398e-08 0 1.15938e-08 0 1.15968e-08 0.0007 1.15998e-08 0 1.16538e-08 0 1.16568e-08 0.0007 1.16598e-08 0 1.17138e-08 0 1.17168e-08 0.0007 1.17198e-08 0 1.17738e-08 0 1.17768e-08 0.0007 1.17798e-08 0 1.18338e-08 0 1.18368e-08 0.0007 1.18398e-08 0 1.18938e-08 0 1.18968e-08 0.0007 1.18998e-08 0 1.19538e-08 0 1.19568e-08 0.0007 1.19598e-08 0 1.20138e-08 0 1.20168e-08 0.0007 1.20198e-08 0 1.20738e-08 0 1.20768e-08 0.0007 1.20798e-08 0 1.21338e-08 0 1.21368e-08 0.0007 1.21398e-08 0 1.21938e-08 0 1.21968e-08 0.0007 1.21998e-08 0 1.22538e-08 0 1.22568e-08 0.0007 1.22598e-08 0 1.23138e-08 0 1.23168e-08 0.0007 1.23198e-08 0 1.23738e-08 0 1.23768e-08 0.0007 1.23798e-08 0 1.24338e-08 0 1.24368e-08 0.0007 1.24398e-08 0 1.24938e-08 0 1.24968e-08 0.0007 1.24998e-08 0 1.25538e-08 0 1.25568e-08 0.0007 1.25598e-08 0 1.26138e-08 0 1.26168e-08 0.0007 1.26198e-08 0 1.26738e-08 0 1.26768e-08 0.0007 1.26798e-08 0 1.27338e-08 0 1.27368e-08 0.0007 1.27398e-08 0 1.27938e-08 0 1.27968e-08 0.0007 1.27998e-08 0 1.28538e-08 0 1.28568e-08 0.0007 1.28598e-08 0 1.29138e-08 0 1.29168e-08 0.0007 1.29198e-08 0 1.29738e-08 0 1.29768e-08 0.0007 1.29798e-08 0 1.30338e-08 0 1.30368e-08 0.0007 1.30398e-08 0 1.30938e-08 0 1.30968e-08 0.0007 1.30998e-08 0 1.31538e-08 0 1.31568e-08 0.0007 1.31598e-08 0 1.32138e-08 0 1.32168e-08 0.0007 1.32198e-08 0 1.32738e-08 0 1.32768e-08 0.0007 1.32798e-08 0 1.33338e-08 0 1.33368e-08 0.0007 1.33398e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.34538e-08 0 1.34568e-08 0.0007 1.34598e-08 0 1.35138e-08 0 1.35168e-08 0.0007 1.35198e-08 0 1.35738e-08 0 1.35768e-08 0.0007 1.35798e-08 0 1.36338e-08 0 1.36368e-08 0.0007 1.36398e-08 0 1.36938e-08 0 1.36968e-08 0.0007 1.36998e-08 0 1.37538e-08 0 1.37568e-08 0.0007 1.37598e-08 0 1.38138e-08 0 1.38168e-08 0.0007 1.38198e-08 0 1.38738e-08 0 1.38768e-08 0.0007 1.38798e-08 0 1.39338e-08 0 1.39368e-08 0.0007 1.39398e-08 0 1.39938e-08 0 1.39968e-08 0.0007 1.39998e-08 0 1.40538e-08 0 1.40568e-08 0.0007 1.40598e-08 0 1.41138e-08 0 1.41168e-08 0.0007 1.41198e-08 0 1.41738e-08 0 1.41768e-08 0.0007 1.41798e-08 0 1.42338e-08 0 1.42368e-08 0.0007 1.42398e-08 0 1.42938e-08 0 1.42968e-08 0.0007 1.42998e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.44138e-08 0 1.44168e-08 0.0007 1.44198e-08 0 1.44738e-08 0 1.44768e-08 0.0007 1.44798e-08 0 1.45338e-08 0 1.45368e-08 0.0007 1.45398e-08 0 1.45938e-08 0 1.45968e-08 0.0007 1.45998e-08 0 1.46538e-08 0 1.46568e-08 0.0007 1.46598e-08 0 1.47138e-08 0 1.47168e-08 0.0007 1.47198e-08 0 1.47738e-08 0 1.47768e-08 0.0007 1.47798e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.48938e-08 0 1.48968e-08 0.0007 1.48998e-08 0 1.49538e-08 0 1.49568e-08 0.0007 1.49598e-08 0 1.50138e-08 0 1.50168e-08 0.0007 1.50198e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.51338e-08 0 1.51368e-08 0.0007 1.51398e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IB3|H 0 B3_TX  PWL(0 0 7.6938e-09 0 7.6968e-09 0.0007 7.6998e-09 0 7.7538e-09 0 7.7568e-09 0.0007 7.7598e-09 0 7.8138e-09 0 7.8168e-09 0.0007 7.8198e-09 0 7.8738e-09 0 7.8768e-09 0.0007 7.8798e-09 0 7.9338e-09 0 7.9368e-09 0.0007 7.9398e-09 0 7.9938e-09 0 7.9968e-09 0.0007 7.9998e-09 0 8.0538e-09 0 8.0568e-09 0.0007 8.0598e-09 0 8.1138e-09 0 8.1168e-09 0.0007 8.1198e-09 0 8.1738e-09 0 8.1768e-09 0.0007 8.1798e-09 0 8.2338e-09 0 8.2368e-09 0.0007 8.2398e-09 0 8.2938e-09 0 8.2968e-09 0.0007 8.2998e-09 0 8.3538e-09 0 8.3568e-09 0.0007 8.3598e-09 0 8.4138e-09 0 8.4168e-09 0.0007 8.4198e-09 0 8.4738e-09 0 8.4768e-09 0.0007 8.4798e-09 0 8.5338e-09 0 8.5368e-09 0.0007 8.5398e-09 0 8.5938e-09 0 8.5968e-09 0.0007 8.5998e-09 0 8.6538e-09 0 8.6568e-09 0.0007 8.6598e-09 0 8.7138e-09 0 8.7168e-09 0.0007 8.7198e-09 0 8.7738e-09 0 8.7768e-09 0.0007 8.7798e-09 0 8.8338e-09 0 8.8368e-09 0.0007 8.8398e-09 0 8.8938e-09 0 8.8968e-09 0.0007 8.8998e-09 0 8.9538e-09 0 8.9568e-09 0.0007 8.9598e-09 0 9.0138e-09 0 9.0168e-09 0.0007 9.0198e-09 0 9.0738e-09 0 9.0768e-09 0.0007 9.0798e-09 0 9.1338e-09 0 9.1368e-09 0.0007 9.1398e-09 0 9.1938e-09 0 9.1968e-09 0.0007 9.1998e-09 0 9.2538e-09 0 9.2568e-09 0.0007 9.2598e-09 0 9.3138e-09 0 9.3168e-09 0.0007 9.3198e-09 0 9.3738e-09 0 9.3768e-09 0.0007 9.3798e-09 0 9.4338e-09 0 9.4368e-09 0.0007 9.4398e-09 0 9.4938e-09 0 9.4968e-09 0.0007 9.4998e-09 0 9.5538e-09 0 9.5568e-09 0.0007 9.5598e-09 0 9.6138e-09 0 9.6168e-09 0.0007 9.6198e-09 0 9.6738e-09 0 9.6768e-09 0.0007 9.6798e-09 0 9.7338e-09 0 9.7368e-09 0.0007 9.7398e-09 0 9.7938e-09 0 9.7968e-09 0.0007 9.7998e-09 0 9.8538e-09 0 9.8568e-09 0.0007 9.8598e-09 0 9.9138e-09 0 9.9168e-09 0.0007 9.9198e-09 0 9.9738e-09 0 9.9768e-09 0.0007 9.9798e-09 0 1.00338e-08 0 1.00368e-08 0.0007 1.00398e-08 0 1.00938e-08 0 1.00968e-08 0.0007 1.00998e-08 0 1.01538e-08 0 1.01568e-08 0.0007 1.01598e-08 0 1.02138e-08 0 1.02168e-08 0.0007 1.02198e-08 0 1.02738e-08 0 1.02768e-08 0.0007 1.02798e-08 0 1.03338e-08 0 1.03368e-08 0.0007 1.03398e-08 0 1.03938e-08 0 1.03968e-08 0.0007 1.03998e-08 0 1.04538e-08 0 1.04568e-08 0.0007 1.04598e-08 0 1.05138e-08 0 1.05168e-08 0.0007 1.05198e-08 0 1.05738e-08 0 1.05768e-08 0.0007 1.05798e-08 0 1.06338e-08 0 1.06368e-08 0.0007 1.06398e-08 0 1.06938e-08 0 1.06968e-08 0.0007 1.06998e-08 0 1.07538e-08 0 1.07568e-08 0.0007 1.07598e-08 0 1.08138e-08 0 1.08168e-08 0.0007 1.08198e-08 0 1.08738e-08 0 1.08768e-08 0.0007 1.08798e-08 0 1.09338e-08 0 1.09368e-08 0.0007 1.09398e-08 0 1.09938e-08 0 1.09968e-08 0.0007 1.09998e-08 0 1.10538e-08 0 1.10568e-08 0.0007 1.10598e-08 0 1.11138e-08 0 1.11168e-08 0.0007 1.11198e-08 0 1.11738e-08 0 1.11768e-08 0.0007 1.11798e-08 0 1.12338e-08 0 1.12368e-08 0.0007 1.12398e-08 0 1.12938e-08 0 1.12968e-08 0.0007 1.12998e-08 0 1.13538e-08 0 1.13568e-08 0.0007 1.13598e-08 0 1.14138e-08 0 1.14168e-08 0.0007 1.14198e-08 0 1.14738e-08 0 1.14768e-08 0.0007 1.14798e-08 0 1.15338e-08 0 1.15368e-08 0.0007 1.15398e-08 0 1.15938e-08 0 1.15968e-08 0.0007 1.15998e-08 0 1.16538e-08 0 1.16568e-08 0.0007 1.16598e-08 0 1.17138e-08 0 1.17168e-08 0.0007 1.17198e-08 0 1.17738e-08 0 1.17768e-08 0.0007 1.17798e-08 0 1.18338e-08 0 1.18368e-08 0.0007 1.18398e-08 0 1.18938e-08 0 1.18968e-08 0.0007 1.18998e-08 0 1.19538e-08 0 1.19568e-08 0.0007 1.19598e-08 0 1.20138e-08 0 1.20168e-08 0.0007 1.20198e-08 0 1.20738e-08 0 1.20768e-08 0.0007 1.20798e-08 0 1.21338e-08 0 1.21368e-08 0.0007 1.21398e-08 0 1.21938e-08 0 1.21968e-08 0.0007 1.21998e-08 0 1.22538e-08 0 1.22568e-08 0.0007 1.22598e-08 0 1.23138e-08 0 1.23168e-08 0.0007 1.23198e-08 0 1.23738e-08 0 1.23768e-08 0.0007 1.23798e-08 0 1.24338e-08 0 1.24368e-08 0.0007 1.24398e-08 0 1.24938e-08 0 1.24968e-08 0.0007 1.24998e-08 0 1.25538e-08 0 1.25568e-08 0.0007 1.25598e-08 0 1.26138e-08 0 1.26168e-08 0.0007 1.26198e-08 0 1.26738e-08 0 1.26768e-08 0.0007 1.26798e-08 0 1.27338e-08 0 1.27368e-08 0.0007 1.27398e-08 0 1.27938e-08 0 1.27968e-08 0.0007 1.27998e-08 0 1.28538e-08 0 1.28568e-08 0.0007 1.28598e-08 0 1.29138e-08 0 1.29168e-08 0.0007 1.29198e-08 0 1.29738e-08 0 1.29768e-08 0.0007 1.29798e-08 0 1.30338e-08 0 1.30368e-08 0.0007 1.30398e-08 0 1.30938e-08 0 1.30968e-08 0.0007 1.30998e-08 0 1.31538e-08 0 1.31568e-08 0.0007 1.31598e-08 0 1.32138e-08 0 1.32168e-08 0.0007 1.32198e-08 0 1.32738e-08 0 1.32768e-08 0.0007 1.32798e-08 0 1.33338e-08 0 1.33368e-08 0.0007 1.33398e-08 0 1.33938e-08 0 1.33968e-08 0.0007 1.33998e-08 0 1.34538e-08 0 1.34568e-08 0.0007 1.34598e-08 0 1.35138e-08 0 1.35168e-08 0.0007 1.35198e-08 0 1.35738e-08 0 1.35768e-08 0.0007 1.35798e-08 0 1.36338e-08 0 1.36368e-08 0.0007 1.36398e-08 0 1.36938e-08 0 1.36968e-08 0.0007 1.36998e-08 0 1.37538e-08 0 1.37568e-08 0.0007 1.37598e-08 0 1.38138e-08 0 1.38168e-08 0.0007 1.38198e-08 0 1.38738e-08 0 1.38768e-08 0.0007 1.38798e-08 0 1.39338e-08 0 1.39368e-08 0.0007 1.39398e-08 0 1.39938e-08 0 1.39968e-08 0.0007 1.39998e-08 0 1.40538e-08 0 1.40568e-08 0.0007 1.40598e-08 0 1.41138e-08 0 1.41168e-08 0.0007 1.41198e-08 0 1.41738e-08 0 1.41768e-08 0.0007 1.41798e-08 0 1.42338e-08 0 1.42368e-08 0.0007 1.42398e-08 0 1.42938e-08 0 1.42968e-08 0.0007 1.42998e-08 0 1.43538e-08 0 1.43568e-08 0.0007 1.43598e-08 0 1.44138e-08 0 1.44168e-08 0.0007 1.44198e-08 0 1.44738e-08 0 1.44768e-08 0.0007 1.44798e-08 0 1.45338e-08 0 1.45368e-08 0.0007 1.45398e-08 0 1.45938e-08 0 1.45968e-08 0.0007 1.45998e-08 0 1.46538e-08 0 1.46568e-08 0.0007 1.46598e-08 0 1.47138e-08 0 1.47168e-08 0.0007 1.47198e-08 0 1.47738e-08 0 1.47768e-08 0.0007 1.47798e-08 0 1.48338e-08 0 1.48368e-08 0.0007 1.48398e-08 0 1.48938e-08 0 1.48968e-08 0.0007 1.48998e-08 0 1.49538e-08 0 1.49568e-08 0.0007 1.49598e-08 0 1.50138e-08 0 1.50168e-08 0.0007 1.50198e-08 0 1.50738e-08 0 1.50768e-08 0.0007 1.50798e-08 0 1.51338e-08 0 1.51368e-08 0.0007 1.51398e-08 0 1.51938e-08 0 1.51968e-08 0.0007 1.51998e-08 0 1.52538e-08 0 1.52568e-08 0.0007 1.52598e-08 0 1.53138e-08 0 1.53168e-08 0.0007 1.53198e-08 0)
IT00|T 0 T00  PWL(0 0 9e-12 0 1.2e-11 0.0021 1.5e-11 0 6.9e-11 0 7.2e-11 0.0021 7.5e-11 0 1.29e-10 0 1.32e-10 0.0021 1.35e-10 0 1.89e-10 0 1.92e-10 0.0021 1.95e-10 0 2.49e-10 0 2.52e-10 0.0021 2.55e-10 0 3.09e-10 0 3.12e-10 0.0021 3.15e-10 0 3.69e-10 0 3.72e-10 0.0021 3.75e-10 0 4.29e-10 0 4.32e-10 0.0021 4.35e-10 0 4.89e-10 0 4.92e-10 0.0021 4.95e-10 0 5.49e-10 0 5.52e-10 0.0021 5.55e-10 0 6.09e-10 0 6.12e-10 0.0021 6.15e-10 0 6.69e-10 0 6.72e-10 0.0021 6.75e-10 0 7.29e-10 0 7.32e-10 0.0021 7.35e-10 0 7.89e-10 0 7.92e-10 0.0021 7.95e-10 0 8.49e-10 0 8.52e-10 0.0021 8.55e-10 0 9.09e-10 0 9.12e-10 0.0021 9.15e-10 0 9.69e-10 0 9.72e-10 0.0021 9.75e-10 0 1.029e-09 0 1.032e-09 0.0021 1.035e-09 0 1.089e-09 0 1.092e-09 0.0021 1.095e-09 0 1.149e-09 0 1.152e-09 0.0021 1.155e-09 0 1.209e-09 0 1.212e-09 0.0021 1.215e-09 0 1.269e-09 0 1.272e-09 0.0021 1.275e-09 0 1.329e-09 0 1.332e-09 0.0021 1.335e-09 0 1.389e-09 0 1.392e-09 0.0021 1.395e-09 0 1.449e-09 0 1.452e-09 0.0021 1.455e-09 0 1.509e-09 0 1.512e-09 0.0021 1.515e-09 0 1.569e-09 0 1.572e-09 0.0021 1.575e-09 0 1.629e-09 0 1.632e-09 0.0021 1.635e-09 0 1.689e-09 0 1.692e-09 0.0021 1.695e-09 0 1.749e-09 0 1.752e-09 0.0021 1.755e-09 0 1.809e-09 0 1.812e-09 0.0021 1.815e-09 0 1.869e-09 0 1.872e-09 0.0021 1.875e-09 0 1.929e-09 0 1.932e-09 0.0021 1.935e-09 0 1.989e-09 0 1.992e-09 0.0021 1.995e-09 0 2.049e-09 0 2.052e-09 0.0021 2.055e-09 0 2.109e-09 0 2.112e-09 0.0021 2.115e-09 0 2.169e-09 0 2.172e-09 0.0021 2.175e-09 0 2.229e-09 0 2.232e-09 0.0021 2.235e-09 0 2.289e-09 0 2.292e-09 0.0021 2.295e-09 0 2.349e-09 0 2.352e-09 0.0021 2.355e-09 0 2.409e-09 0 2.412e-09 0.0021 2.415e-09 0 2.469e-09 0 2.472e-09 0.0021 2.475e-09 0 2.529e-09 0 2.532e-09 0.0021 2.535e-09 0 2.589e-09 0 2.592e-09 0.0021 2.595e-09 0 2.649e-09 0 2.652e-09 0.0021 2.655e-09 0 2.709e-09 0 2.712e-09 0.0021 2.715e-09 0 2.769e-09 0 2.772e-09 0.0021 2.775e-09 0 2.829e-09 0 2.832e-09 0.0021 2.835e-09 0 2.889e-09 0 2.892e-09 0.0021 2.895e-09 0 2.949e-09 0 2.952e-09 0.0021 2.955e-09 0 3.009e-09 0 3.012e-09 0.0021 3.015e-09 0 3.069e-09 0 3.072e-09 0.0021 3.075e-09 0 3.129e-09 0 3.132e-09 0.0021 3.135e-09 0 3.189e-09 0 3.192e-09 0.0021 3.195e-09 0 3.249e-09 0 3.252e-09 0.0021 3.255e-09 0 3.309e-09 0 3.312e-09 0.0021 3.315e-09 0 3.369e-09 0 3.372e-09 0.0021 3.375e-09 0 3.429e-09 0 3.432e-09 0.0021 3.435e-09 0 3.489e-09 0 3.492e-09 0.0021 3.495e-09 0 3.549e-09 0 3.552e-09 0.0021 3.555e-09 0 3.609e-09 0 3.612e-09 0.0021 3.615e-09 0 3.669e-09 0 3.672e-09 0.0021 3.675e-09 0 3.729e-09 0 3.732e-09 0.0021 3.735e-09 0 3.789e-09 0 3.792e-09 0.0021 3.795e-09 0 3.849e-09 0 3.852e-09 0.0021 3.855e-09 0 3.909e-09 0 3.912e-09 0.0021 3.915e-09 0 3.969e-09 0 3.972e-09 0.0021 3.975e-09 0 4.029e-09 0 4.032e-09 0.0021 4.035e-09 0 4.089e-09 0 4.092e-09 0.0021 4.095e-09 0 4.149e-09 0 4.152e-09 0.0021 4.155e-09 0 4.209e-09 0 4.212e-09 0.0021 4.215e-09 0 4.269e-09 0 4.272e-09 0.0021 4.275e-09 0 4.329e-09 0 4.332e-09 0.0021 4.335e-09 0 4.389e-09 0 4.392e-09 0.0021 4.395e-09 0 4.449e-09 0 4.452e-09 0.0021 4.455e-09 0 4.509e-09 0 4.512e-09 0.0021 4.515e-09 0 4.569e-09 0 4.572e-09 0.0021 4.575e-09 0 4.629e-09 0 4.632e-09 0.0021 4.635e-09 0 4.689e-09 0 4.692e-09 0.0021 4.695e-09 0 4.749e-09 0 4.752e-09 0.0021 4.755e-09 0 4.809e-09 0 4.812e-09 0.0021 4.815e-09 0 4.869e-09 0 4.872e-09 0.0021 4.875e-09 0 4.929e-09 0 4.932e-09 0.0021 4.935e-09 0 4.989e-09 0 4.992e-09 0.0021 4.995e-09 0 5.049e-09 0 5.052e-09 0.0021 5.055e-09 0 5.109e-09 0 5.112e-09 0.0021 5.115e-09 0 5.169e-09 0 5.172e-09 0.0021 5.175e-09 0 5.229e-09 0 5.232e-09 0.0021 5.235e-09 0 5.289e-09 0 5.292e-09 0.0021 5.295e-09 0 5.349e-09 0 5.352e-09 0.0021 5.355e-09 0 5.409e-09 0 5.412e-09 0.0021 5.415e-09 0 5.469e-09 0 5.472e-09 0.0021 5.475e-09 0 5.529e-09 0 5.532e-09 0.0021 5.535e-09 0 5.589e-09 0 5.592e-09 0.0021 5.595e-09 0 5.649e-09 0 5.652e-09 0.0021 5.655e-09 0 5.709e-09 0 5.712e-09 0.0021 5.715e-09 0 5.769e-09 0 5.772e-09 0.0021 5.775e-09 0 5.829e-09 0 5.832e-09 0.0021 5.835e-09 0 5.889e-09 0 5.892e-09 0.0021 5.895e-09 0 5.949e-09 0 5.952e-09 0.0021 5.955e-09 0 6.009e-09 0 6.012e-09 0.0021 6.015e-09 0 6.069e-09 0 6.072e-09 0.0021 6.075e-09 0 6.129e-09 0 6.132e-09 0.0021 6.135e-09 0 6.189e-09 0 6.192e-09 0.0021 6.195e-09 0 6.249e-09 0 6.252e-09 0.0021 6.255e-09 0 6.309e-09 0 6.312e-09 0.0021 6.315e-09 0 6.369e-09 0 6.372e-09 0.0021 6.375e-09 0 6.429e-09 0 6.432e-09 0.0021 6.435e-09 0 6.489e-09 0 6.492e-09 0.0021 6.495e-09 0 6.549e-09 0 6.552e-09 0.0021 6.555e-09 0 6.609e-09 0 6.612e-09 0.0021 6.615e-09 0 6.669e-09 0 6.672e-09 0.0021 6.675e-09 0 6.729e-09 0 6.732e-09 0.0021 6.735e-09 0 6.789e-09 0 6.792e-09 0.0021 6.795e-09 0 6.849e-09 0 6.852e-09 0.0021 6.855e-09 0 6.909e-09 0 6.912e-09 0.0021 6.915e-09 0 6.969e-09 0 6.972e-09 0.0021 6.975e-09 0 7.029e-09 0 7.032e-09 0.0021 7.035e-09 0 7.089e-09 0 7.092e-09 0.0021 7.095e-09 0 7.149e-09 0 7.152e-09 0.0021 7.155e-09 0 7.209e-09 0 7.212e-09 0.0021 7.215e-09 0 7.269e-09 0 7.272e-09 0.0021 7.275e-09 0 7.329e-09 0 7.332e-09 0.0021 7.335e-09 0 7.389e-09 0 7.392e-09 0.0021 7.395e-09 0 7.449e-09 0 7.452e-09 0.0021 7.455e-09 0 7.509e-09 0 7.512e-09 0.0021 7.515e-09 0 7.569e-09 0 7.572e-09 0.0021 7.575e-09 0 7.629e-09 0 7.632e-09 0.0021 7.635e-09 0 7.689e-09 0 7.692e-09 0.0021 7.695e-09 0 7.749e-09 0 7.752e-09 0.0021 7.755e-09 0 7.809e-09 0 7.812e-09 0.0021 7.815e-09 0 7.869e-09 0 7.872e-09 0.0021 7.875e-09 0 7.929e-09 0 7.932e-09 0.0021 7.935e-09 0 7.989e-09 0 7.992e-09 0.0021 7.995e-09 0 8.049e-09 0 8.052e-09 0.0021 8.055e-09 0 8.109e-09 0 8.112e-09 0.0021 8.115e-09 0 8.169e-09 0 8.172e-09 0.0021 8.175e-09 0 8.229e-09 0 8.232e-09 0.0021 8.235e-09 0 8.289e-09 0 8.292e-09 0.0021 8.295e-09 0 8.349e-09 0 8.352e-09 0.0021 8.355e-09 0 8.409e-09 0 8.412e-09 0.0021 8.415e-09 0 8.469e-09 0 8.472e-09 0.0021 8.475e-09 0 8.529e-09 0 8.532e-09 0.0021 8.535e-09 0 8.589e-09 0 8.592e-09 0.0021 8.595e-09 0 8.649e-09 0 8.652e-09 0.0021 8.655e-09 0 8.709e-09 0 8.712e-09 0.0021 8.715e-09 0 8.769e-09 0 8.772e-09 0.0021 8.775e-09 0 8.829e-09 0 8.832e-09 0.0021 8.835e-09 0 8.889e-09 0 8.892e-09 0.0021 8.895e-09 0 8.949e-09 0 8.952e-09 0.0021 8.955e-09 0 9.009e-09 0 9.012e-09 0.0021 9.015e-09 0 9.069e-09 0 9.072e-09 0.0021 9.075e-09 0 9.129e-09 0 9.132e-09 0.0021 9.135e-09 0 9.189e-09 0 9.192e-09 0.0021 9.195e-09 0 9.249e-09 0 9.252e-09 0.0021 9.255e-09 0 9.309e-09 0 9.312e-09 0.0021 9.315e-09 0 9.369e-09 0 9.372e-09 0.0021 9.375e-09 0 9.429e-09 0 9.432e-09 0.0021 9.435e-09 0 9.489e-09 0 9.492e-09 0.0021 9.495e-09 0 9.549e-09 0 9.552e-09 0.0021 9.555e-09 0 9.609e-09 0 9.612e-09 0.0021 9.615e-09 0 9.669e-09 0 9.672e-09 0.0021 9.675e-09 0 9.729e-09 0 9.732e-09 0.0021 9.735e-09 0 9.789e-09 0 9.792e-09 0.0021 9.795e-09 0 9.849e-09 0 9.852e-09 0.0021 9.855e-09 0 9.909e-09 0 9.912e-09 0.0021 9.915e-09 0 9.969e-09 0 9.972e-09 0.0021 9.975e-09 0 1.0029e-08 0 1.0032e-08 0.0021 1.0035e-08 0 1.0089e-08 0 1.0092e-08 0.0021 1.0095e-08 0 1.0149e-08 0 1.0152e-08 0.0021 1.0155e-08 0 1.0209e-08 0 1.0212e-08 0.0021 1.0215e-08 0 1.0269e-08 0 1.0272e-08 0.0021 1.0275e-08 0 1.0329e-08 0 1.0332e-08 0.0021 1.0335e-08 0 1.0389e-08 0 1.0392e-08 0.0021 1.0395e-08 0 1.0449e-08 0 1.0452e-08 0.0021 1.0455e-08 0 1.0509e-08 0 1.0512e-08 0.0021 1.0515e-08 0 1.0569e-08 0 1.0572e-08 0.0021 1.0575e-08 0 1.0629e-08 0 1.0632e-08 0.0021 1.0635e-08 0 1.0689e-08 0 1.0692e-08 0.0021 1.0695e-08 0 1.0749e-08 0 1.0752e-08 0.0021 1.0755e-08 0 1.0809e-08 0 1.0812e-08 0.0021 1.0815e-08 0 1.0869e-08 0 1.0872e-08 0.0021 1.0875e-08 0 1.0929e-08 0 1.0932e-08 0.0021 1.0935e-08 0 1.0989e-08 0 1.0992e-08 0.0021 1.0995e-08 0 1.1049e-08 0 1.1052e-08 0.0021 1.1055e-08 0 1.1109e-08 0 1.1112e-08 0.0021 1.1115e-08 0 1.1169e-08 0 1.1172e-08 0.0021 1.1175e-08 0 1.1229e-08 0 1.1232e-08 0.0021 1.1235e-08 0 1.1289e-08 0 1.1292e-08 0.0021 1.1295e-08 0 1.1349e-08 0 1.1352e-08 0.0021 1.1355e-08 0 1.1409e-08 0 1.1412e-08 0.0021 1.1415e-08 0 1.1469e-08 0 1.1472e-08 0.0021 1.1475e-08 0 1.1529e-08 0 1.1532e-08 0.0021 1.1535e-08 0 1.1589e-08 0 1.1592e-08 0.0021 1.1595e-08 0 1.1649e-08 0 1.1652e-08 0.0021 1.1655e-08 0 1.1709e-08 0 1.1712e-08 0.0021 1.1715e-08 0 1.1769e-08 0 1.1772e-08 0.0021 1.1775e-08 0 1.1829e-08 0 1.1832e-08 0.0021 1.1835e-08 0 1.1889e-08 0 1.1892e-08 0.0021 1.1895e-08 0 1.1949e-08 0 1.1952e-08 0.0021 1.1955e-08 0 1.2009e-08 0 1.2012e-08 0.0021 1.2015e-08 0 1.2069e-08 0 1.2072e-08 0.0021 1.2075e-08 0 1.2129e-08 0 1.2132e-08 0.0021 1.2135e-08 0 1.2189e-08 0 1.2192e-08 0.0021 1.2195e-08 0 1.2249e-08 0 1.2252e-08 0.0021 1.2255e-08 0 1.2309e-08 0 1.2312e-08 0.0021 1.2315e-08 0 1.2369e-08 0 1.2372e-08 0.0021 1.2375e-08 0 1.2429e-08 0 1.2432e-08 0.0021 1.2435e-08 0 1.2489e-08 0 1.2492e-08 0.0021 1.2495e-08 0 1.2549e-08 0 1.2552e-08 0.0021 1.2555e-08 0 1.2609e-08 0 1.2612e-08 0.0021 1.2615e-08 0 1.2669e-08 0 1.2672e-08 0.0021 1.2675e-08 0 1.2729e-08 0 1.2732e-08 0.0021 1.2735e-08 0 1.2789e-08 0 1.2792e-08 0.0021 1.2795e-08 0 1.2849e-08 0 1.2852e-08 0.0021 1.2855e-08 0 1.2909e-08 0 1.2912e-08 0.0021 1.2915e-08 0 1.2969e-08 0 1.2972e-08 0.0021 1.2975e-08 0 1.3029e-08 0 1.3032e-08 0.0021 1.3035e-08 0 1.3089e-08 0 1.3092e-08 0.0021 1.3095e-08 0 1.3149e-08 0 1.3152e-08 0.0021 1.3155e-08 0 1.3209e-08 0 1.3212e-08 0.0021 1.3215e-08 0 1.3269e-08 0 1.3272e-08 0.0021 1.3275e-08 0 1.3329e-08 0 1.3332e-08 0.0021 1.3335e-08 0 1.3389e-08 0 1.3392e-08 0.0021 1.3395e-08 0 1.3449e-08 0 1.3452e-08 0.0021 1.3455e-08 0 1.3509e-08 0 1.3512e-08 0.0021 1.3515e-08 0 1.3569e-08 0 1.3572e-08 0.0021 1.3575e-08 0 1.3629e-08 0 1.3632e-08 0.0021 1.3635e-08 0 1.3689e-08 0 1.3692e-08 0.0021 1.3695e-08 0 1.3749e-08 0 1.3752e-08 0.0021 1.3755e-08 0 1.3809e-08 0 1.3812e-08 0.0021 1.3815e-08 0 1.3869e-08 0 1.3872e-08 0.0021 1.3875e-08 0 1.3929e-08 0 1.3932e-08 0.0021 1.3935e-08 0 1.3989e-08 0 1.3992e-08 0.0021 1.3995e-08 0 1.4049e-08 0 1.4052e-08 0.0021 1.4055e-08 0 1.4109e-08 0 1.4112e-08 0.0021 1.4115e-08 0 1.4169e-08 0 1.4172e-08 0.0021 1.4175e-08 0 1.4229e-08 0 1.4232e-08 0.0021 1.4235e-08 0 1.4289e-08 0 1.4292e-08 0.0021 1.4295e-08 0 1.4349e-08 0 1.4352e-08 0.0021 1.4355e-08 0 1.4409e-08 0 1.4412e-08 0.0021 1.4415e-08 0 1.4469e-08 0 1.4472e-08 0.0021 1.4475e-08 0 1.4529e-08 0 1.4532e-08 0.0021 1.4535e-08 0 1.4589e-08 0 1.4592e-08 0.0021 1.4595e-08 0 1.4649e-08 0 1.4652e-08 0.0021 1.4655e-08 0 1.4709e-08 0 1.4712e-08 0.0021 1.4715e-08 0 1.4769e-08 0 1.4772e-08 0.0021 1.4775e-08 0 1.4829e-08 0 1.4832e-08 0.0021 1.4835e-08 0 1.4889e-08 0 1.4892e-08 0.0021 1.4895e-08 0 1.4949e-08 0 1.4952e-08 0.0021 1.4955e-08 0 1.5009e-08 0 1.5012e-08 0.0021 1.5015e-08 0 1.5069e-08 0 1.5072e-08 0.0021 1.5075e-08 0 1.5129e-08 0 1.5132e-08 0.0021 1.5135e-08 0 1.5189e-08 0 1.5192e-08 0.0021 1.5195e-08 0 1.5249e-08 0 1.5252e-08 0.0021 1.5255e-08 0 1.5309e-08 0 1.5312e-08 0.0021 1.5315e-08 0 1.5369e-08 0 1.5372e-08 0.0021 1.5375e-08 0 1.5429e-08 0 1.5432e-08 0.0021 1.5435e-08 0 1.5489e-08 0 1.5492e-08 0.0021 1.5495e-08 0 1.5549e-08 0 1.5552e-08 0.0021 1.5555e-08 0 1.5609e-08 0 1.5612e-08 0.0021 1.5615e-08 0 1.5669e-08 0 1.5672e-08 0.0021 1.5675e-08 0 1.5729e-08 0 1.5732e-08 0.0021 1.5735e-08 0 1.5789e-08 0 1.5792e-08 0.0021 1.5795e-08 0 1.5849e-08 0 1.5852e-08 0.0021 1.5855e-08 0 1.5909e-08 0 1.5912e-08 0.0021 1.5915e-08 0 1.5969e-08 0 1.5972e-08 0.0021 1.5975e-08 0 1.6029e-08 0 1.6032e-08 0.0021 1.6035e-08 0 1.6089e-08 0 1.6092e-08 0.0021 1.6095e-08 0 1.6149e-08 0 1.6152e-08 0.0021 1.6155e-08 0 1.6209e-08 0 1.6212e-08 0.0021 1.6215e-08 0 1.6269e-08 0 1.6272e-08 0.0021 1.6275e-08 0 1.6329e-08 0 1.6332e-08 0.0021 1.6335e-08 0 1.6389e-08 0 1.6392e-08 0.0021 1.6395e-08 0 1.6449e-08 0 1.6452e-08 0.0021 1.6455e-08 0 1.6509e-08 0 1.6512e-08 0.0021 1.6515e-08 0 1.6569e-08 0 1.6572e-08 0.0021 1.6575e-08 0 1.6629e-08 0 1.6632e-08 0.0021 1.6635e-08 0 1.6689e-08 0 1.6692e-08 0.0021 1.6695e-08 0 1.6749e-08 0 1.6752e-08 0.0021 1.6755e-08 0 1.6809e-08 0 1.6812e-08 0.0021 1.6815e-08 0 1.6869e-08 0 1.6872e-08 0.0021 1.6875e-08 0 1.6929e-08 0 1.6932e-08 0.0021 1.6935e-08 0 1.6989e-08 0 1.6992e-08 0.0021 1.6995e-08 0 1.7049e-08 0 1.7052e-08 0.0021 1.7055e-08 0 1.7109e-08 0 1.7112e-08 0.0021 1.7115e-08 0 1.7169e-08 0 1.7172e-08 0.0021 1.7175e-08 0 1.7229e-08 0 1.7232e-08 0.0021 1.7235e-08 0 1.7289e-08 0 1.7292e-08 0.0021 1.7295e-08 0 1.7349e-08 0 1.7352e-08 0.0021 1.7355e-08 0 1.7409e-08 0 1.7412e-08 0.0021 1.7415e-08 0 1.7469e-08 0 1.7472e-08 0.0021 1.7475e-08 0 1.7529e-08 0 1.7532e-08 0.0021 1.7535e-08 0 1.7589e-08 0 1.7592e-08 0.0021 1.7595e-08 0 1.7649e-08 0 1.7652e-08 0.0021 1.7655e-08 0 1.7709e-08 0 1.7712e-08 0.0021 1.7715e-08 0 1.7769e-08 0 1.7772e-08 0.0021 1.7775e-08 0 1.7829e-08 0 1.7832e-08 0.0021 1.7835e-08 0 1.7889e-08 0 1.7892e-08 0.0021 1.7895e-08 0 1.7949e-08 0 1.7952e-08 0.0021 1.7955e-08 0 1.8009e-08 0 1.8012e-08 0.0021 1.8015e-08 0 1.8069e-08 0 1.8072e-08 0.0021 1.8075e-08 0 1.8129e-08 0 1.8132e-08 0.0021 1.8135e-08 0 1.8189e-08 0 1.8192e-08 0.0021 1.8195e-08 0 1.8249e-08 0 1.8252e-08 0.0021 1.8255e-08 0 1.8309e-08 0 1.8312e-08 0.0021 1.8315e-08 0 1.8369e-08 0 1.8372e-08 0.0021 1.8375e-08 0 1.8429e-08 0 1.8432e-08 0.0021 1.8435e-08 0 1.8489e-08 0 1.8492e-08 0.0021 1.8495e-08 0 1.8549e-08 0 1.8552e-08 0.0021 1.8555e-08 0 1.8609e-08 0 1.8612e-08 0.0021 1.8615e-08 0 1.8669e-08 0 1.8672e-08 0.0021 1.8675e-08 0 1.8729e-08 0 1.8732e-08 0.0021 1.8735e-08 0 1.8789e-08 0 1.8792e-08 0.0021 1.8795e-08 0 1.8849e-08 0 1.8852e-08 0.0021 1.8855e-08 0 1.8909e-08 0 1.8912e-08 0.0021 1.8915e-08 0 1.8969e-08 0 1.8972e-08 0.0021 1.8975e-08 0 1.9029e-08 0 1.9032e-08 0.0021 1.9035e-08 0 1.9089e-08 0 1.9092e-08 0.0021 1.9095e-08 0 1.9149e-08 0 1.9152e-08 0.0021 1.9155e-08 0 1.9209e-08 0 1.9212e-08 0.0021 1.9215e-08 0 1.9269e-08 0 1.9272e-08 0.0021 1.9275e-08 0 1.9329e-08 0 1.9332e-08 0.0021 1.9335e-08 0 1.9389e-08 0 1.9392e-08 0.0021 1.9395e-08 0 1.9449e-08 0 1.9452e-08 0.0021 1.9455e-08 0 1.9509e-08 0 1.9512e-08 0.0021 1.9515e-08 0 1.9569e-08 0 1.9572e-08 0.0021 1.9575e-08 0 1.9629e-08 0 1.9632e-08 0.0021 1.9635e-08 0 1.9689e-08 0 1.9692e-08 0.0021 1.9695e-08 0 1.9749e-08 0 1.9752e-08 0.0021 1.9755e-08 0 1.9809e-08 0 1.9812e-08 0.0021 1.9815e-08 0 1.9869e-08 0 1.9872e-08 0.0021 1.9875e-08 0 1.9929e-08 0 1.9932e-08 0.0021 1.9935e-08 0 1.9989e-08 0 1.9992e-08 0.0021 1.9995e-08 0 2.0049e-08 0 2.0052e-08 0.0021 2.0055e-08 0 2.0109e-08 0 2.0112e-08 0.0021 2.0115e-08 0 2.0169e-08 0 2.0172e-08 0.0021 2.0175e-08 0 2.0229e-08 0 2.0232e-08 0.0021 2.0235e-08 0 2.0289e-08 0 2.0292e-08 0.0021 2.0295e-08 0 2.0349e-08 0 2.0352e-08 0.0021 2.0355e-08 0 2.0409e-08 0 2.0412e-08 0.0021 2.0415e-08 0 2.0469e-08 0 2.0472e-08 0.0021 2.0475e-08 0 2.0529e-08 0 2.0532e-08 0.0021 2.0535e-08 0 2.0589e-08 0 2.0592e-08 0.0021 2.0595e-08 0 2.0649e-08 0 2.0652e-08 0.0021 2.0655e-08 0 2.0709e-08 0 2.0712e-08 0.0021 2.0715e-08 0 2.0769e-08 0 2.0772e-08 0.0021 2.0775e-08 0 2.0829e-08 0 2.0832e-08 0.0021 2.0835e-08 0 2.0889e-08 0 2.0892e-08 0.0021 2.0895e-08 0 2.0949e-08 0 2.0952e-08 0.0021 2.0955e-08 0 2.1009e-08 0 2.1012e-08 0.0021 2.1015e-08 0 2.1069e-08 0 2.1072e-08 0.0021 2.1075e-08 0 2.1129e-08 0 2.1132e-08 0.0021 2.1135e-08 0 2.1189e-08 0 2.1192e-08 0.0021 2.1195e-08 0 2.1249e-08 0 2.1252e-08 0.0021 2.1255e-08 0 2.1309e-08 0 2.1312e-08 0.0021 2.1315e-08 0 2.1369e-08 0 2.1372e-08 0.0021 2.1375e-08 0 2.1429e-08 0 2.1432e-08 0.0021 2.1435e-08 0 2.1489e-08 0 2.1492e-08 0.0021 2.1495e-08 0 2.1549e-08 0 2.1552e-08 0.0021 2.1555e-08 0 2.1609e-08 0 2.1612e-08 0.0021 2.1615e-08 0 2.1669e-08 0 2.1672e-08 0.0021 2.1675e-08 0 2.1729e-08 0 2.1732e-08 0.0021 2.1735e-08 0 2.1789e-08 0 2.1792e-08 0.0021 2.1795e-08 0 2.1849e-08 0 2.1852e-08 0.0021 2.1855e-08 0 2.1909e-08 0 2.1912e-08 0.0021 2.1915e-08 0 2.1969e-08 0 2.1972e-08 0.0021 2.1975e-08 0 2.2029e-08 0 2.2032e-08 0.0021 2.2035e-08 0 2.2089e-08 0 2.2092e-08 0.0021 2.2095e-08 0 2.2149e-08 0 2.2152e-08 0.0021 2.2155e-08 0 2.2209e-08 0 2.2212e-08 0.0021 2.2215e-08 0 2.2269e-08 0 2.2272e-08 0.0021 2.2275e-08 0 2.2329e-08 0 2.2332e-08 0.0021 2.2335e-08 0 2.2389e-08 0 2.2392e-08 0.0021 2.2395e-08 0 2.2449e-08 0 2.2452e-08 0.0021 2.2455e-08 0 2.2509e-08 0 2.2512e-08 0.0021 2.2515e-08 0 2.2569e-08 0 2.2572e-08 0.0021 2.2575e-08 0 2.2629e-08 0 2.2632e-08 0.0021 2.2635e-08 0 2.2689e-08 0 2.2692e-08 0.0021 2.2695e-08 0 2.2749e-08 0 2.2752e-08 0.0021 2.2755e-08 0 2.2809e-08 0 2.2812e-08 0.0021 2.2815e-08 0 2.2869e-08 0 2.2872e-08 0.0021 2.2875e-08 0 2.2929e-08 0 2.2932e-08 0.0021 2.2935e-08 0 2.2989e-08 0 2.2992e-08 0.0021 2.2995e-08 0 2.3049e-08 0 2.3052e-08 0.0021 2.3055e-08 0 2.3109e-08 0 2.3112e-08 0.0021 2.3115e-08 0 2.3169e-08 0 2.3172e-08 0.0021 2.3175e-08 0 2.3229e-08 0 2.3232e-08 0.0021 2.3235e-08 0 2.3289e-08 0 2.3292e-08 0.0021 2.3295e-08 0 2.3349e-08 0 2.3352e-08 0.0021 2.3355e-08 0 2.3409e-08 0 2.3412e-08 0.0021 2.3415e-08 0 2.3469e-08 0 2.3472e-08 0.0021 2.3475e-08 0 2.3529e-08 0 2.3532e-08 0.0021 2.3535e-08 0 2.3589e-08 0 2.3592e-08 0.0021 2.3595e-08 0 2.3649e-08 0 2.3652e-08 0.0021 2.3655e-08 0 2.3709e-08 0 2.3712e-08 0.0021 2.3715e-08 0 2.3769e-08 0 2.3772e-08 0.0021 2.3775e-08 0 2.3829e-08 0 2.3832e-08 0.0021 2.3835e-08 0 2.3889e-08 0 2.3892e-08 0.0021 2.3895e-08 0)
IT01|T 0 T01  PWL(0 0 9e-12 0 1.2e-11 0.0021 1.5e-11 0 6.9e-11 0 7.2e-11 0.0021 7.5e-11 0 1.29e-10 0 1.32e-10 0.0021 1.35e-10 0 1.89e-10 0 1.92e-10 0.0021 1.95e-10 0 2.49e-10 0 2.52e-10 0.0021 2.55e-10 0 3.09e-10 0 3.12e-10 0.0021 3.15e-10 0 3.69e-10 0 3.72e-10 0.0021 3.75e-10 0 4.29e-10 0 4.32e-10 0.0021 4.35e-10 0 4.89e-10 0 4.92e-10 0.0021 4.95e-10 0 5.49e-10 0 5.52e-10 0.0021 5.55e-10 0 6.09e-10 0 6.12e-10 0.0021 6.15e-10 0 6.69e-10 0 6.72e-10 0.0021 6.75e-10 0 7.29e-10 0 7.32e-10 0.0021 7.35e-10 0 7.89e-10 0 7.92e-10 0.0021 7.95e-10 0 8.49e-10 0 8.52e-10 0.0021 8.55e-10 0 9.09e-10 0 9.12e-10 0.0021 9.15e-10 0 9.69e-10 0 9.72e-10 0.0021 9.75e-10 0 1.029e-09 0 1.032e-09 0.0021 1.035e-09 0 1.089e-09 0 1.092e-09 0.0021 1.095e-09 0 1.149e-09 0 1.152e-09 0.0021 1.155e-09 0 1.209e-09 0 1.212e-09 0.0021 1.215e-09 0 1.269e-09 0 1.272e-09 0.0021 1.275e-09 0 1.329e-09 0 1.332e-09 0.0021 1.335e-09 0 1.389e-09 0 1.392e-09 0.0021 1.395e-09 0 1.449e-09 0 1.452e-09 0.0021 1.455e-09 0 1.509e-09 0 1.512e-09 0.0021 1.515e-09 0 1.569e-09 0 1.572e-09 0.0021 1.575e-09 0 1.629e-09 0 1.632e-09 0.0021 1.635e-09 0 1.689e-09 0 1.692e-09 0.0021 1.695e-09 0 1.749e-09 0 1.752e-09 0.0021 1.755e-09 0 1.809e-09 0 1.812e-09 0.0021 1.815e-09 0 1.869e-09 0 1.872e-09 0.0021 1.875e-09 0 1.929e-09 0 1.932e-09 0.0021 1.935e-09 0 1.989e-09 0 1.992e-09 0.0021 1.995e-09 0 2.049e-09 0 2.052e-09 0.0021 2.055e-09 0 2.109e-09 0 2.112e-09 0.0021 2.115e-09 0 2.169e-09 0 2.172e-09 0.0021 2.175e-09 0 2.229e-09 0 2.232e-09 0.0021 2.235e-09 0 2.289e-09 0 2.292e-09 0.0021 2.295e-09 0 2.349e-09 0 2.352e-09 0.0021 2.355e-09 0 2.409e-09 0 2.412e-09 0.0021 2.415e-09 0 2.469e-09 0 2.472e-09 0.0021 2.475e-09 0 2.529e-09 0 2.532e-09 0.0021 2.535e-09 0 2.589e-09 0 2.592e-09 0.0021 2.595e-09 0 2.649e-09 0 2.652e-09 0.0021 2.655e-09 0 2.709e-09 0 2.712e-09 0.0021 2.715e-09 0 2.769e-09 0 2.772e-09 0.0021 2.775e-09 0 2.829e-09 0 2.832e-09 0.0021 2.835e-09 0 2.889e-09 0 2.892e-09 0.0021 2.895e-09 0 2.949e-09 0 2.952e-09 0.0021 2.955e-09 0 3.009e-09 0 3.012e-09 0.0021 3.015e-09 0 3.069e-09 0 3.072e-09 0.0021 3.075e-09 0 3.129e-09 0 3.132e-09 0.0021 3.135e-09 0 3.189e-09 0 3.192e-09 0.0021 3.195e-09 0 3.249e-09 0 3.252e-09 0.0021 3.255e-09 0 3.309e-09 0 3.312e-09 0.0021 3.315e-09 0 3.369e-09 0 3.372e-09 0.0021 3.375e-09 0 3.429e-09 0 3.432e-09 0.0021 3.435e-09 0 3.489e-09 0 3.492e-09 0.0021 3.495e-09 0 3.549e-09 0 3.552e-09 0.0021 3.555e-09 0 3.609e-09 0 3.612e-09 0.0021 3.615e-09 0 3.669e-09 0 3.672e-09 0.0021 3.675e-09 0 3.729e-09 0 3.732e-09 0.0021 3.735e-09 0 3.789e-09 0 3.792e-09 0.0021 3.795e-09 0 3.849e-09 0 3.852e-09 0.0021 3.855e-09 0 3.909e-09 0 3.912e-09 0.0021 3.915e-09 0 3.969e-09 0 3.972e-09 0.0021 3.975e-09 0 4.029e-09 0 4.032e-09 0.0021 4.035e-09 0 4.089e-09 0 4.092e-09 0.0021 4.095e-09 0 4.149e-09 0 4.152e-09 0.0021 4.155e-09 0 4.209e-09 0 4.212e-09 0.0021 4.215e-09 0 4.269e-09 0 4.272e-09 0.0021 4.275e-09 0 4.329e-09 0 4.332e-09 0.0021 4.335e-09 0 4.389e-09 0 4.392e-09 0.0021 4.395e-09 0 4.449e-09 0 4.452e-09 0.0021 4.455e-09 0 4.509e-09 0 4.512e-09 0.0021 4.515e-09 0 4.569e-09 0 4.572e-09 0.0021 4.575e-09 0 4.629e-09 0 4.632e-09 0.0021 4.635e-09 0 4.689e-09 0 4.692e-09 0.0021 4.695e-09 0 4.749e-09 0 4.752e-09 0.0021 4.755e-09 0 4.809e-09 0 4.812e-09 0.0021 4.815e-09 0 4.869e-09 0 4.872e-09 0.0021 4.875e-09 0 4.929e-09 0 4.932e-09 0.0021 4.935e-09 0 4.989e-09 0 4.992e-09 0.0021 4.995e-09 0 5.049e-09 0 5.052e-09 0.0021 5.055e-09 0 5.109e-09 0 5.112e-09 0.0021 5.115e-09 0 5.169e-09 0 5.172e-09 0.0021 5.175e-09 0 5.229e-09 0 5.232e-09 0.0021 5.235e-09 0 5.289e-09 0 5.292e-09 0.0021 5.295e-09 0 5.349e-09 0 5.352e-09 0.0021 5.355e-09 0 5.409e-09 0 5.412e-09 0.0021 5.415e-09 0 5.469e-09 0 5.472e-09 0.0021 5.475e-09 0 5.529e-09 0 5.532e-09 0.0021 5.535e-09 0 5.589e-09 0 5.592e-09 0.0021 5.595e-09 0 5.649e-09 0 5.652e-09 0.0021 5.655e-09 0 5.709e-09 0 5.712e-09 0.0021 5.715e-09 0 5.769e-09 0 5.772e-09 0.0021 5.775e-09 0 5.829e-09 0 5.832e-09 0.0021 5.835e-09 0 5.889e-09 0 5.892e-09 0.0021 5.895e-09 0 5.949e-09 0 5.952e-09 0.0021 5.955e-09 0 6.009e-09 0 6.012e-09 0.0021 6.015e-09 0 6.069e-09 0 6.072e-09 0.0021 6.075e-09 0 6.129e-09 0 6.132e-09 0.0021 6.135e-09 0 6.189e-09 0 6.192e-09 0.0021 6.195e-09 0 6.249e-09 0 6.252e-09 0.0021 6.255e-09 0 6.309e-09 0 6.312e-09 0.0021 6.315e-09 0 6.369e-09 0 6.372e-09 0.0021 6.375e-09 0 6.429e-09 0 6.432e-09 0.0021 6.435e-09 0 6.489e-09 0 6.492e-09 0.0021 6.495e-09 0 6.549e-09 0 6.552e-09 0.0021 6.555e-09 0 6.609e-09 0 6.612e-09 0.0021 6.615e-09 0 6.669e-09 0 6.672e-09 0.0021 6.675e-09 0 6.729e-09 0 6.732e-09 0.0021 6.735e-09 0 6.789e-09 0 6.792e-09 0.0021 6.795e-09 0 6.849e-09 0 6.852e-09 0.0021 6.855e-09 0 6.909e-09 0 6.912e-09 0.0021 6.915e-09 0 6.969e-09 0 6.972e-09 0.0021 6.975e-09 0 7.029e-09 0 7.032e-09 0.0021 7.035e-09 0 7.089e-09 0 7.092e-09 0.0021 7.095e-09 0 7.149e-09 0 7.152e-09 0.0021 7.155e-09 0 7.209e-09 0 7.212e-09 0.0021 7.215e-09 0 7.269e-09 0 7.272e-09 0.0021 7.275e-09 0 7.329e-09 0 7.332e-09 0.0021 7.335e-09 0 7.389e-09 0 7.392e-09 0.0021 7.395e-09 0 7.449e-09 0 7.452e-09 0.0021 7.455e-09 0 7.509e-09 0 7.512e-09 0.0021 7.515e-09 0 7.569e-09 0 7.572e-09 0.0021 7.575e-09 0 7.629e-09 0 7.632e-09 0.0021 7.635e-09 0 7.689e-09 0 7.692e-09 0.0021 7.695e-09 0 7.749e-09 0 7.752e-09 0.0021 7.755e-09 0 7.809e-09 0 7.812e-09 0.0021 7.815e-09 0 7.869e-09 0 7.872e-09 0.0021 7.875e-09 0 7.929e-09 0 7.932e-09 0.0021 7.935e-09 0 7.989e-09 0 7.992e-09 0.0021 7.995e-09 0 8.049e-09 0 8.052e-09 0.0021 8.055e-09 0 8.109e-09 0 8.112e-09 0.0021 8.115e-09 0 8.169e-09 0 8.172e-09 0.0021 8.175e-09 0 8.229e-09 0 8.232e-09 0.0021 8.235e-09 0 8.289e-09 0 8.292e-09 0.0021 8.295e-09 0 8.349e-09 0 8.352e-09 0.0021 8.355e-09 0 8.409e-09 0 8.412e-09 0.0021 8.415e-09 0 8.469e-09 0 8.472e-09 0.0021 8.475e-09 0 8.529e-09 0 8.532e-09 0.0021 8.535e-09 0 8.589e-09 0 8.592e-09 0.0021 8.595e-09 0 8.649e-09 0 8.652e-09 0.0021 8.655e-09 0 8.709e-09 0 8.712e-09 0.0021 8.715e-09 0 8.769e-09 0 8.772e-09 0.0021 8.775e-09 0 8.829e-09 0 8.832e-09 0.0021 8.835e-09 0 8.889e-09 0 8.892e-09 0.0021 8.895e-09 0 8.949e-09 0 8.952e-09 0.0021 8.955e-09 0 9.009e-09 0 9.012e-09 0.0021 9.015e-09 0 9.069e-09 0 9.072e-09 0.0021 9.075e-09 0 9.129e-09 0 9.132e-09 0.0021 9.135e-09 0 9.189e-09 0 9.192e-09 0.0021 9.195e-09 0 9.249e-09 0 9.252e-09 0.0021 9.255e-09 0 9.309e-09 0 9.312e-09 0.0021 9.315e-09 0 9.369e-09 0 9.372e-09 0.0021 9.375e-09 0 9.429e-09 0 9.432e-09 0.0021 9.435e-09 0 9.489e-09 0 9.492e-09 0.0021 9.495e-09 0 9.549e-09 0 9.552e-09 0.0021 9.555e-09 0 9.609e-09 0 9.612e-09 0.0021 9.615e-09 0 9.669e-09 0 9.672e-09 0.0021 9.675e-09 0 9.729e-09 0 9.732e-09 0.0021 9.735e-09 0 9.789e-09 0 9.792e-09 0.0021 9.795e-09 0 9.849e-09 0 9.852e-09 0.0021 9.855e-09 0 9.909e-09 0 9.912e-09 0.0021 9.915e-09 0 9.969e-09 0 9.972e-09 0.0021 9.975e-09 0 1.0029e-08 0 1.0032e-08 0.0021 1.0035e-08 0 1.0089e-08 0 1.0092e-08 0.0021 1.0095e-08 0 1.0149e-08 0 1.0152e-08 0.0021 1.0155e-08 0 1.0209e-08 0 1.0212e-08 0.0021 1.0215e-08 0 1.0269e-08 0 1.0272e-08 0.0021 1.0275e-08 0 1.0329e-08 0 1.0332e-08 0.0021 1.0335e-08 0 1.0389e-08 0 1.0392e-08 0.0021 1.0395e-08 0 1.0449e-08 0 1.0452e-08 0.0021 1.0455e-08 0 1.0509e-08 0 1.0512e-08 0.0021 1.0515e-08 0 1.0569e-08 0 1.0572e-08 0.0021 1.0575e-08 0 1.0629e-08 0 1.0632e-08 0.0021 1.0635e-08 0 1.0689e-08 0 1.0692e-08 0.0021 1.0695e-08 0 1.0749e-08 0 1.0752e-08 0.0021 1.0755e-08 0 1.0809e-08 0 1.0812e-08 0.0021 1.0815e-08 0 1.0869e-08 0 1.0872e-08 0.0021 1.0875e-08 0 1.0929e-08 0 1.0932e-08 0.0021 1.0935e-08 0 1.0989e-08 0 1.0992e-08 0.0021 1.0995e-08 0 1.1049e-08 0 1.1052e-08 0.0021 1.1055e-08 0 1.1109e-08 0 1.1112e-08 0.0021 1.1115e-08 0 1.1169e-08 0 1.1172e-08 0.0021 1.1175e-08 0 1.1229e-08 0 1.1232e-08 0.0021 1.1235e-08 0 1.1289e-08 0 1.1292e-08 0.0021 1.1295e-08 0 1.1349e-08 0 1.1352e-08 0.0021 1.1355e-08 0 1.1409e-08 0 1.1412e-08 0.0021 1.1415e-08 0 1.1469e-08 0 1.1472e-08 0.0021 1.1475e-08 0 1.1529e-08 0 1.1532e-08 0.0021 1.1535e-08 0 1.1589e-08 0 1.1592e-08 0.0021 1.1595e-08 0 1.1649e-08 0 1.1652e-08 0.0021 1.1655e-08 0 1.1709e-08 0 1.1712e-08 0.0021 1.1715e-08 0 1.1769e-08 0 1.1772e-08 0.0021 1.1775e-08 0 1.1829e-08 0 1.1832e-08 0.0021 1.1835e-08 0 1.1889e-08 0 1.1892e-08 0.0021 1.1895e-08 0 1.1949e-08 0 1.1952e-08 0.0021 1.1955e-08 0 1.2009e-08 0 1.2012e-08 0.0021 1.2015e-08 0 1.2069e-08 0 1.2072e-08 0.0021 1.2075e-08 0 1.2129e-08 0 1.2132e-08 0.0021 1.2135e-08 0 1.2189e-08 0 1.2192e-08 0.0021 1.2195e-08 0 1.2249e-08 0 1.2252e-08 0.0021 1.2255e-08 0 1.2309e-08 0 1.2312e-08 0.0021 1.2315e-08 0 1.2369e-08 0 1.2372e-08 0.0021 1.2375e-08 0 1.2429e-08 0 1.2432e-08 0.0021 1.2435e-08 0 1.2489e-08 0 1.2492e-08 0.0021 1.2495e-08 0 1.2549e-08 0 1.2552e-08 0.0021 1.2555e-08 0 1.2609e-08 0 1.2612e-08 0.0021 1.2615e-08 0 1.2669e-08 0 1.2672e-08 0.0021 1.2675e-08 0 1.2729e-08 0 1.2732e-08 0.0021 1.2735e-08 0 1.2789e-08 0 1.2792e-08 0.0021 1.2795e-08 0 1.2849e-08 0 1.2852e-08 0.0021 1.2855e-08 0 1.2909e-08 0 1.2912e-08 0.0021 1.2915e-08 0 1.2969e-08 0 1.2972e-08 0.0021 1.2975e-08 0 1.3029e-08 0 1.3032e-08 0.0021 1.3035e-08 0 1.3089e-08 0 1.3092e-08 0.0021 1.3095e-08 0 1.3149e-08 0 1.3152e-08 0.0021 1.3155e-08 0 1.3209e-08 0 1.3212e-08 0.0021 1.3215e-08 0 1.3269e-08 0 1.3272e-08 0.0021 1.3275e-08 0 1.3329e-08 0 1.3332e-08 0.0021 1.3335e-08 0 1.3389e-08 0 1.3392e-08 0.0021 1.3395e-08 0 1.3449e-08 0 1.3452e-08 0.0021 1.3455e-08 0 1.3509e-08 0 1.3512e-08 0.0021 1.3515e-08 0 1.3569e-08 0 1.3572e-08 0.0021 1.3575e-08 0 1.3629e-08 0 1.3632e-08 0.0021 1.3635e-08 0 1.3689e-08 0 1.3692e-08 0.0021 1.3695e-08 0 1.3749e-08 0 1.3752e-08 0.0021 1.3755e-08 0 1.3809e-08 0 1.3812e-08 0.0021 1.3815e-08 0 1.3869e-08 0 1.3872e-08 0.0021 1.3875e-08 0 1.3929e-08 0 1.3932e-08 0.0021 1.3935e-08 0 1.3989e-08 0 1.3992e-08 0.0021 1.3995e-08 0 1.4049e-08 0 1.4052e-08 0.0021 1.4055e-08 0 1.4109e-08 0 1.4112e-08 0.0021 1.4115e-08 0 1.4169e-08 0 1.4172e-08 0.0021 1.4175e-08 0 1.4229e-08 0 1.4232e-08 0.0021 1.4235e-08 0 1.4289e-08 0 1.4292e-08 0.0021 1.4295e-08 0 1.4349e-08 0 1.4352e-08 0.0021 1.4355e-08 0 1.4409e-08 0 1.4412e-08 0.0021 1.4415e-08 0 1.4469e-08 0 1.4472e-08 0.0021 1.4475e-08 0 1.4529e-08 0 1.4532e-08 0.0021 1.4535e-08 0 1.4589e-08 0 1.4592e-08 0.0021 1.4595e-08 0 1.4649e-08 0 1.4652e-08 0.0021 1.4655e-08 0 1.4709e-08 0 1.4712e-08 0.0021 1.4715e-08 0 1.4769e-08 0 1.4772e-08 0.0021 1.4775e-08 0 1.4829e-08 0 1.4832e-08 0.0021 1.4835e-08 0 1.4889e-08 0 1.4892e-08 0.0021 1.4895e-08 0 1.4949e-08 0 1.4952e-08 0.0021 1.4955e-08 0 1.5009e-08 0 1.5012e-08 0.0021 1.5015e-08 0 1.5069e-08 0 1.5072e-08 0.0021 1.5075e-08 0 1.5129e-08 0 1.5132e-08 0.0021 1.5135e-08 0 1.5189e-08 0 1.5192e-08 0.0021 1.5195e-08 0 1.5249e-08 0 1.5252e-08 0.0021 1.5255e-08 0 1.5309e-08 0 1.5312e-08 0.0021 1.5315e-08 0 1.5369e-08 0 1.5372e-08 0.0021 1.5375e-08 0 1.5429e-08 0 1.5432e-08 0.0021 1.5435e-08 0 1.5489e-08 0 1.5492e-08 0.0021 1.5495e-08 0 1.5549e-08 0 1.5552e-08 0.0021 1.5555e-08 0 1.5609e-08 0 1.5612e-08 0.0021 1.5615e-08 0 1.5669e-08 0 1.5672e-08 0.0021 1.5675e-08 0 1.5729e-08 0 1.5732e-08 0.0021 1.5735e-08 0 1.5789e-08 0 1.5792e-08 0.0021 1.5795e-08 0 1.5849e-08 0 1.5852e-08 0.0021 1.5855e-08 0 1.5909e-08 0 1.5912e-08 0.0021 1.5915e-08 0 1.5969e-08 0 1.5972e-08 0.0021 1.5975e-08 0 1.6029e-08 0 1.6032e-08 0.0021 1.6035e-08 0 1.6089e-08 0 1.6092e-08 0.0021 1.6095e-08 0 1.6149e-08 0 1.6152e-08 0.0021 1.6155e-08 0 1.6209e-08 0 1.6212e-08 0.0021 1.6215e-08 0 1.6269e-08 0 1.6272e-08 0.0021 1.6275e-08 0 1.6329e-08 0 1.6332e-08 0.0021 1.6335e-08 0 1.6389e-08 0 1.6392e-08 0.0021 1.6395e-08 0 1.6449e-08 0 1.6452e-08 0.0021 1.6455e-08 0 1.6509e-08 0 1.6512e-08 0.0021 1.6515e-08 0 1.6569e-08 0 1.6572e-08 0.0021 1.6575e-08 0 1.6629e-08 0 1.6632e-08 0.0021 1.6635e-08 0 1.6689e-08 0 1.6692e-08 0.0021 1.6695e-08 0 1.6749e-08 0 1.6752e-08 0.0021 1.6755e-08 0 1.6809e-08 0 1.6812e-08 0.0021 1.6815e-08 0 1.6869e-08 0 1.6872e-08 0.0021 1.6875e-08 0 1.6929e-08 0 1.6932e-08 0.0021 1.6935e-08 0 1.6989e-08 0 1.6992e-08 0.0021 1.6995e-08 0 1.7049e-08 0 1.7052e-08 0.0021 1.7055e-08 0 1.7109e-08 0 1.7112e-08 0.0021 1.7115e-08 0 1.7169e-08 0 1.7172e-08 0.0021 1.7175e-08 0 1.7229e-08 0 1.7232e-08 0.0021 1.7235e-08 0 1.7289e-08 0 1.7292e-08 0.0021 1.7295e-08 0 1.7349e-08 0 1.7352e-08 0.0021 1.7355e-08 0 1.7409e-08 0 1.7412e-08 0.0021 1.7415e-08 0 1.7469e-08 0 1.7472e-08 0.0021 1.7475e-08 0 1.7529e-08 0 1.7532e-08 0.0021 1.7535e-08 0 1.7589e-08 0 1.7592e-08 0.0021 1.7595e-08 0 1.7649e-08 0 1.7652e-08 0.0021 1.7655e-08 0 1.7709e-08 0 1.7712e-08 0.0021 1.7715e-08 0 1.7769e-08 0 1.7772e-08 0.0021 1.7775e-08 0 1.7829e-08 0 1.7832e-08 0.0021 1.7835e-08 0 1.7889e-08 0 1.7892e-08 0.0021 1.7895e-08 0 1.7949e-08 0 1.7952e-08 0.0021 1.7955e-08 0 1.8009e-08 0 1.8012e-08 0.0021 1.8015e-08 0 1.8069e-08 0 1.8072e-08 0.0021 1.8075e-08 0 1.8129e-08 0 1.8132e-08 0.0021 1.8135e-08 0 1.8189e-08 0 1.8192e-08 0.0021 1.8195e-08 0 1.8249e-08 0 1.8252e-08 0.0021 1.8255e-08 0 1.8309e-08 0 1.8312e-08 0.0021 1.8315e-08 0 1.8369e-08 0 1.8372e-08 0.0021 1.8375e-08 0 1.8429e-08 0 1.8432e-08 0.0021 1.8435e-08 0 1.8489e-08 0 1.8492e-08 0.0021 1.8495e-08 0 1.8549e-08 0 1.8552e-08 0.0021 1.8555e-08 0 1.8609e-08 0 1.8612e-08 0.0021 1.8615e-08 0 1.8669e-08 0 1.8672e-08 0.0021 1.8675e-08 0 1.8729e-08 0 1.8732e-08 0.0021 1.8735e-08 0 1.8789e-08 0 1.8792e-08 0.0021 1.8795e-08 0 1.8849e-08 0 1.8852e-08 0.0021 1.8855e-08 0 1.8909e-08 0 1.8912e-08 0.0021 1.8915e-08 0 1.8969e-08 0 1.8972e-08 0.0021 1.8975e-08 0 1.9029e-08 0 1.9032e-08 0.0021 1.9035e-08 0 1.9089e-08 0 1.9092e-08 0.0021 1.9095e-08 0 1.9149e-08 0 1.9152e-08 0.0021 1.9155e-08 0 1.9209e-08 0 1.9212e-08 0.0021 1.9215e-08 0 1.9269e-08 0 1.9272e-08 0.0021 1.9275e-08 0 1.9329e-08 0 1.9332e-08 0.0021 1.9335e-08 0 1.9389e-08 0 1.9392e-08 0.0021 1.9395e-08 0 1.9449e-08 0 1.9452e-08 0.0021 1.9455e-08 0 1.9509e-08 0 1.9512e-08 0.0021 1.9515e-08 0 1.9569e-08 0 1.9572e-08 0.0021 1.9575e-08 0 1.9629e-08 0 1.9632e-08 0.0021 1.9635e-08 0 1.9689e-08 0 1.9692e-08 0.0021 1.9695e-08 0 1.9749e-08 0 1.9752e-08 0.0021 1.9755e-08 0 1.9809e-08 0 1.9812e-08 0.0021 1.9815e-08 0 1.9869e-08 0 1.9872e-08 0.0021 1.9875e-08 0 1.9929e-08 0 1.9932e-08 0.0021 1.9935e-08 0 1.9989e-08 0 1.9992e-08 0.0021 1.9995e-08 0 2.0049e-08 0 2.0052e-08 0.0021 2.0055e-08 0 2.0109e-08 0 2.0112e-08 0.0021 2.0115e-08 0 2.0169e-08 0 2.0172e-08 0.0021 2.0175e-08 0 2.0229e-08 0 2.0232e-08 0.0021 2.0235e-08 0 2.0289e-08 0 2.0292e-08 0.0021 2.0295e-08 0 2.0349e-08 0 2.0352e-08 0.0021 2.0355e-08 0 2.0409e-08 0 2.0412e-08 0.0021 2.0415e-08 0 2.0469e-08 0 2.0472e-08 0.0021 2.0475e-08 0 2.0529e-08 0 2.0532e-08 0.0021 2.0535e-08 0 2.0589e-08 0 2.0592e-08 0.0021 2.0595e-08 0 2.0649e-08 0 2.0652e-08 0.0021 2.0655e-08 0 2.0709e-08 0 2.0712e-08 0.0021 2.0715e-08 0 2.0769e-08 0 2.0772e-08 0.0021 2.0775e-08 0 2.0829e-08 0 2.0832e-08 0.0021 2.0835e-08 0 2.0889e-08 0 2.0892e-08 0.0021 2.0895e-08 0 2.0949e-08 0 2.0952e-08 0.0021 2.0955e-08 0 2.1009e-08 0 2.1012e-08 0.0021 2.1015e-08 0 2.1069e-08 0 2.1072e-08 0.0021 2.1075e-08 0 2.1129e-08 0 2.1132e-08 0.0021 2.1135e-08 0 2.1189e-08 0 2.1192e-08 0.0021 2.1195e-08 0 2.1249e-08 0 2.1252e-08 0.0021 2.1255e-08 0 2.1309e-08 0 2.1312e-08 0.0021 2.1315e-08 0 2.1369e-08 0 2.1372e-08 0.0021 2.1375e-08 0 2.1429e-08 0 2.1432e-08 0.0021 2.1435e-08 0 2.1489e-08 0 2.1492e-08 0.0021 2.1495e-08 0 2.1549e-08 0 2.1552e-08 0.0021 2.1555e-08 0 2.1609e-08 0 2.1612e-08 0.0021 2.1615e-08 0 2.1669e-08 0 2.1672e-08 0.0021 2.1675e-08 0 2.1729e-08 0 2.1732e-08 0.0021 2.1735e-08 0 2.1789e-08 0 2.1792e-08 0.0021 2.1795e-08 0 2.1849e-08 0 2.1852e-08 0.0021 2.1855e-08 0 2.1909e-08 0 2.1912e-08 0.0021 2.1915e-08 0 2.1969e-08 0 2.1972e-08 0.0021 2.1975e-08 0 2.2029e-08 0 2.2032e-08 0.0021 2.2035e-08 0 2.2089e-08 0 2.2092e-08 0.0021 2.2095e-08 0 2.2149e-08 0 2.2152e-08 0.0021 2.2155e-08 0 2.2209e-08 0 2.2212e-08 0.0021 2.2215e-08 0 2.2269e-08 0 2.2272e-08 0.0021 2.2275e-08 0 2.2329e-08 0 2.2332e-08 0.0021 2.2335e-08 0 2.2389e-08 0 2.2392e-08 0.0021 2.2395e-08 0 2.2449e-08 0 2.2452e-08 0.0021 2.2455e-08 0 2.2509e-08 0 2.2512e-08 0.0021 2.2515e-08 0 2.2569e-08 0 2.2572e-08 0.0021 2.2575e-08 0 2.2629e-08 0 2.2632e-08 0.0021 2.2635e-08 0 2.2689e-08 0 2.2692e-08 0.0021 2.2695e-08 0 2.2749e-08 0 2.2752e-08 0.0021 2.2755e-08 0 2.2809e-08 0 2.2812e-08 0.0021 2.2815e-08 0 2.2869e-08 0 2.2872e-08 0.0021 2.2875e-08 0 2.2929e-08 0 2.2932e-08 0.0021 2.2935e-08 0 2.2989e-08 0 2.2992e-08 0.0021 2.2995e-08 0 2.3049e-08 0 2.3052e-08 0.0021 2.3055e-08 0 2.3109e-08 0 2.3112e-08 0.0021 2.3115e-08 0 2.3169e-08 0 2.3172e-08 0.0021 2.3175e-08 0 2.3229e-08 0 2.3232e-08 0.0021 2.3235e-08 0 2.3289e-08 0 2.3292e-08 0.0021 2.3295e-08 0 2.3349e-08 0 2.3352e-08 0.0021 2.3355e-08 0 2.3409e-08 0 2.3412e-08 0.0021 2.3415e-08 0 2.3469e-08 0 2.3472e-08 0.0021 2.3475e-08 0 2.3529e-08 0 2.3532e-08 0.0021 2.3535e-08 0 2.3589e-08 0 2.3592e-08 0.0021 2.3595e-08 0 2.3649e-08 0 2.3652e-08 0.0021 2.3655e-08 0 2.3709e-08 0 2.3712e-08 0.0021 2.3715e-08 0 2.3769e-08 0 2.3772e-08 0.0021 2.3775e-08 0 2.3829e-08 0 2.3832e-08 0.0021 2.3835e-08 0 2.3889e-08 0 2.3892e-08 0.0021 2.3895e-08 0)
IT02|T 0 T02  PWL(0 0 9e-12 0 1.2e-11 0.0021 1.5e-11 0 6.9e-11 0 7.2e-11 0.0021 7.5e-11 0 1.29e-10 0 1.32e-10 0.0021 1.35e-10 0 1.89e-10 0 1.92e-10 0.0021 1.95e-10 0 2.49e-10 0 2.52e-10 0.0021 2.55e-10 0 3.09e-10 0 3.12e-10 0.0021 3.15e-10 0 3.69e-10 0 3.72e-10 0.0021 3.75e-10 0 4.29e-10 0 4.32e-10 0.0021 4.35e-10 0 4.89e-10 0 4.92e-10 0.0021 4.95e-10 0 5.49e-10 0 5.52e-10 0.0021 5.55e-10 0 6.09e-10 0 6.12e-10 0.0021 6.15e-10 0 6.69e-10 0 6.72e-10 0.0021 6.75e-10 0 7.29e-10 0 7.32e-10 0.0021 7.35e-10 0 7.89e-10 0 7.92e-10 0.0021 7.95e-10 0 8.49e-10 0 8.52e-10 0.0021 8.55e-10 0 9.09e-10 0 9.12e-10 0.0021 9.15e-10 0 9.69e-10 0 9.72e-10 0.0021 9.75e-10 0 1.029e-09 0 1.032e-09 0.0021 1.035e-09 0 1.089e-09 0 1.092e-09 0.0021 1.095e-09 0 1.149e-09 0 1.152e-09 0.0021 1.155e-09 0 1.209e-09 0 1.212e-09 0.0021 1.215e-09 0 1.269e-09 0 1.272e-09 0.0021 1.275e-09 0 1.329e-09 0 1.332e-09 0.0021 1.335e-09 0 1.389e-09 0 1.392e-09 0.0021 1.395e-09 0 1.449e-09 0 1.452e-09 0.0021 1.455e-09 0 1.509e-09 0 1.512e-09 0.0021 1.515e-09 0 1.569e-09 0 1.572e-09 0.0021 1.575e-09 0 1.629e-09 0 1.632e-09 0.0021 1.635e-09 0 1.689e-09 0 1.692e-09 0.0021 1.695e-09 0 1.749e-09 0 1.752e-09 0.0021 1.755e-09 0 1.809e-09 0 1.812e-09 0.0021 1.815e-09 0 1.869e-09 0 1.872e-09 0.0021 1.875e-09 0 1.929e-09 0 1.932e-09 0.0021 1.935e-09 0 1.989e-09 0 1.992e-09 0.0021 1.995e-09 0 2.049e-09 0 2.052e-09 0.0021 2.055e-09 0 2.109e-09 0 2.112e-09 0.0021 2.115e-09 0 2.169e-09 0 2.172e-09 0.0021 2.175e-09 0 2.229e-09 0 2.232e-09 0.0021 2.235e-09 0 2.289e-09 0 2.292e-09 0.0021 2.295e-09 0 2.349e-09 0 2.352e-09 0.0021 2.355e-09 0 2.409e-09 0 2.412e-09 0.0021 2.415e-09 0 2.469e-09 0 2.472e-09 0.0021 2.475e-09 0 2.529e-09 0 2.532e-09 0.0021 2.535e-09 0 2.589e-09 0 2.592e-09 0.0021 2.595e-09 0 2.649e-09 0 2.652e-09 0.0021 2.655e-09 0 2.709e-09 0 2.712e-09 0.0021 2.715e-09 0 2.769e-09 0 2.772e-09 0.0021 2.775e-09 0 2.829e-09 0 2.832e-09 0.0021 2.835e-09 0 2.889e-09 0 2.892e-09 0.0021 2.895e-09 0 2.949e-09 0 2.952e-09 0.0021 2.955e-09 0 3.009e-09 0 3.012e-09 0.0021 3.015e-09 0 3.069e-09 0 3.072e-09 0.0021 3.075e-09 0 3.129e-09 0 3.132e-09 0.0021 3.135e-09 0 3.189e-09 0 3.192e-09 0.0021 3.195e-09 0 3.249e-09 0 3.252e-09 0.0021 3.255e-09 0 3.309e-09 0 3.312e-09 0.0021 3.315e-09 0 3.369e-09 0 3.372e-09 0.0021 3.375e-09 0 3.429e-09 0 3.432e-09 0.0021 3.435e-09 0 3.489e-09 0 3.492e-09 0.0021 3.495e-09 0 3.549e-09 0 3.552e-09 0.0021 3.555e-09 0 3.609e-09 0 3.612e-09 0.0021 3.615e-09 0 3.669e-09 0 3.672e-09 0.0021 3.675e-09 0 3.729e-09 0 3.732e-09 0.0021 3.735e-09 0 3.789e-09 0 3.792e-09 0.0021 3.795e-09 0 3.849e-09 0 3.852e-09 0.0021 3.855e-09 0 3.909e-09 0 3.912e-09 0.0021 3.915e-09 0 3.969e-09 0 3.972e-09 0.0021 3.975e-09 0 4.029e-09 0 4.032e-09 0.0021 4.035e-09 0 4.089e-09 0 4.092e-09 0.0021 4.095e-09 0 4.149e-09 0 4.152e-09 0.0021 4.155e-09 0 4.209e-09 0 4.212e-09 0.0021 4.215e-09 0 4.269e-09 0 4.272e-09 0.0021 4.275e-09 0 4.329e-09 0 4.332e-09 0.0021 4.335e-09 0 4.389e-09 0 4.392e-09 0.0021 4.395e-09 0 4.449e-09 0 4.452e-09 0.0021 4.455e-09 0 4.509e-09 0 4.512e-09 0.0021 4.515e-09 0 4.569e-09 0 4.572e-09 0.0021 4.575e-09 0 4.629e-09 0 4.632e-09 0.0021 4.635e-09 0 4.689e-09 0 4.692e-09 0.0021 4.695e-09 0 4.749e-09 0 4.752e-09 0.0021 4.755e-09 0 4.809e-09 0 4.812e-09 0.0021 4.815e-09 0 4.869e-09 0 4.872e-09 0.0021 4.875e-09 0 4.929e-09 0 4.932e-09 0.0021 4.935e-09 0 4.989e-09 0 4.992e-09 0.0021 4.995e-09 0 5.049e-09 0 5.052e-09 0.0021 5.055e-09 0 5.109e-09 0 5.112e-09 0.0021 5.115e-09 0 5.169e-09 0 5.172e-09 0.0021 5.175e-09 0 5.229e-09 0 5.232e-09 0.0021 5.235e-09 0 5.289e-09 0 5.292e-09 0.0021 5.295e-09 0 5.349e-09 0 5.352e-09 0.0021 5.355e-09 0 5.409e-09 0 5.412e-09 0.0021 5.415e-09 0 5.469e-09 0 5.472e-09 0.0021 5.475e-09 0 5.529e-09 0 5.532e-09 0.0021 5.535e-09 0 5.589e-09 0 5.592e-09 0.0021 5.595e-09 0 5.649e-09 0 5.652e-09 0.0021 5.655e-09 0 5.709e-09 0 5.712e-09 0.0021 5.715e-09 0 5.769e-09 0 5.772e-09 0.0021 5.775e-09 0 5.829e-09 0 5.832e-09 0.0021 5.835e-09 0 5.889e-09 0 5.892e-09 0.0021 5.895e-09 0 5.949e-09 0 5.952e-09 0.0021 5.955e-09 0 6.009e-09 0 6.012e-09 0.0021 6.015e-09 0 6.069e-09 0 6.072e-09 0.0021 6.075e-09 0 6.129e-09 0 6.132e-09 0.0021 6.135e-09 0 6.189e-09 0 6.192e-09 0.0021 6.195e-09 0 6.249e-09 0 6.252e-09 0.0021 6.255e-09 0 6.309e-09 0 6.312e-09 0.0021 6.315e-09 0 6.369e-09 0 6.372e-09 0.0021 6.375e-09 0 6.429e-09 0 6.432e-09 0.0021 6.435e-09 0 6.489e-09 0 6.492e-09 0.0021 6.495e-09 0 6.549e-09 0 6.552e-09 0.0021 6.555e-09 0 6.609e-09 0 6.612e-09 0.0021 6.615e-09 0 6.669e-09 0 6.672e-09 0.0021 6.675e-09 0 6.729e-09 0 6.732e-09 0.0021 6.735e-09 0 6.789e-09 0 6.792e-09 0.0021 6.795e-09 0 6.849e-09 0 6.852e-09 0.0021 6.855e-09 0 6.909e-09 0 6.912e-09 0.0021 6.915e-09 0 6.969e-09 0 6.972e-09 0.0021 6.975e-09 0 7.029e-09 0 7.032e-09 0.0021 7.035e-09 0 7.089e-09 0 7.092e-09 0.0021 7.095e-09 0 7.149e-09 0 7.152e-09 0.0021 7.155e-09 0 7.209e-09 0 7.212e-09 0.0021 7.215e-09 0 7.269e-09 0 7.272e-09 0.0021 7.275e-09 0 7.329e-09 0 7.332e-09 0.0021 7.335e-09 0 7.389e-09 0 7.392e-09 0.0021 7.395e-09 0 7.449e-09 0 7.452e-09 0.0021 7.455e-09 0 7.509e-09 0 7.512e-09 0.0021 7.515e-09 0 7.569e-09 0 7.572e-09 0.0021 7.575e-09 0 7.629e-09 0 7.632e-09 0.0021 7.635e-09 0 7.689e-09 0 7.692e-09 0.0021 7.695e-09 0 7.749e-09 0 7.752e-09 0.0021 7.755e-09 0 7.809e-09 0 7.812e-09 0.0021 7.815e-09 0 7.869e-09 0 7.872e-09 0.0021 7.875e-09 0 7.929e-09 0 7.932e-09 0.0021 7.935e-09 0 7.989e-09 0 7.992e-09 0.0021 7.995e-09 0 8.049e-09 0 8.052e-09 0.0021 8.055e-09 0 8.109e-09 0 8.112e-09 0.0021 8.115e-09 0 8.169e-09 0 8.172e-09 0.0021 8.175e-09 0 8.229e-09 0 8.232e-09 0.0021 8.235e-09 0 8.289e-09 0 8.292e-09 0.0021 8.295e-09 0 8.349e-09 0 8.352e-09 0.0021 8.355e-09 0 8.409e-09 0 8.412e-09 0.0021 8.415e-09 0 8.469e-09 0 8.472e-09 0.0021 8.475e-09 0 8.529e-09 0 8.532e-09 0.0021 8.535e-09 0 8.589e-09 0 8.592e-09 0.0021 8.595e-09 0 8.649e-09 0 8.652e-09 0.0021 8.655e-09 0 8.709e-09 0 8.712e-09 0.0021 8.715e-09 0 8.769e-09 0 8.772e-09 0.0021 8.775e-09 0 8.829e-09 0 8.832e-09 0.0021 8.835e-09 0 8.889e-09 0 8.892e-09 0.0021 8.895e-09 0 8.949e-09 0 8.952e-09 0.0021 8.955e-09 0 9.009e-09 0 9.012e-09 0.0021 9.015e-09 0 9.069e-09 0 9.072e-09 0.0021 9.075e-09 0 9.129e-09 0 9.132e-09 0.0021 9.135e-09 0 9.189e-09 0 9.192e-09 0.0021 9.195e-09 0 9.249e-09 0 9.252e-09 0.0021 9.255e-09 0 9.309e-09 0 9.312e-09 0.0021 9.315e-09 0 9.369e-09 0 9.372e-09 0.0021 9.375e-09 0 9.429e-09 0 9.432e-09 0.0021 9.435e-09 0 9.489e-09 0 9.492e-09 0.0021 9.495e-09 0 9.549e-09 0 9.552e-09 0.0021 9.555e-09 0 9.609e-09 0 9.612e-09 0.0021 9.615e-09 0 9.669e-09 0 9.672e-09 0.0021 9.675e-09 0 9.729e-09 0 9.732e-09 0.0021 9.735e-09 0 9.789e-09 0 9.792e-09 0.0021 9.795e-09 0 9.849e-09 0 9.852e-09 0.0021 9.855e-09 0 9.909e-09 0 9.912e-09 0.0021 9.915e-09 0 9.969e-09 0 9.972e-09 0.0021 9.975e-09 0 1.0029e-08 0 1.0032e-08 0.0021 1.0035e-08 0 1.0089e-08 0 1.0092e-08 0.0021 1.0095e-08 0 1.0149e-08 0 1.0152e-08 0.0021 1.0155e-08 0 1.0209e-08 0 1.0212e-08 0.0021 1.0215e-08 0 1.0269e-08 0 1.0272e-08 0.0021 1.0275e-08 0 1.0329e-08 0 1.0332e-08 0.0021 1.0335e-08 0 1.0389e-08 0 1.0392e-08 0.0021 1.0395e-08 0 1.0449e-08 0 1.0452e-08 0.0021 1.0455e-08 0 1.0509e-08 0 1.0512e-08 0.0021 1.0515e-08 0 1.0569e-08 0 1.0572e-08 0.0021 1.0575e-08 0 1.0629e-08 0 1.0632e-08 0.0021 1.0635e-08 0 1.0689e-08 0 1.0692e-08 0.0021 1.0695e-08 0 1.0749e-08 0 1.0752e-08 0.0021 1.0755e-08 0 1.0809e-08 0 1.0812e-08 0.0021 1.0815e-08 0 1.0869e-08 0 1.0872e-08 0.0021 1.0875e-08 0 1.0929e-08 0 1.0932e-08 0.0021 1.0935e-08 0 1.0989e-08 0 1.0992e-08 0.0021 1.0995e-08 0 1.1049e-08 0 1.1052e-08 0.0021 1.1055e-08 0 1.1109e-08 0 1.1112e-08 0.0021 1.1115e-08 0 1.1169e-08 0 1.1172e-08 0.0021 1.1175e-08 0 1.1229e-08 0 1.1232e-08 0.0021 1.1235e-08 0 1.1289e-08 0 1.1292e-08 0.0021 1.1295e-08 0 1.1349e-08 0 1.1352e-08 0.0021 1.1355e-08 0 1.1409e-08 0 1.1412e-08 0.0021 1.1415e-08 0 1.1469e-08 0 1.1472e-08 0.0021 1.1475e-08 0 1.1529e-08 0 1.1532e-08 0.0021 1.1535e-08 0 1.1589e-08 0 1.1592e-08 0.0021 1.1595e-08 0 1.1649e-08 0 1.1652e-08 0.0021 1.1655e-08 0 1.1709e-08 0 1.1712e-08 0.0021 1.1715e-08 0 1.1769e-08 0 1.1772e-08 0.0021 1.1775e-08 0 1.1829e-08 0 1.1832e-08 0.0021 1.1835e-08 0 1.1889e-08 0 1.1892e-08 0.0021 1.1895e-08 0 1.1949e-08 0 1.1952e-08 0.0021 1.1955e-08 0 1.2009e-08 0 1.2012e-08 0.0021 1.2015e-08 0 1.2069e-08 0 1.2072e-08 0.0021 1.2075e-08 0 1.2129e-08 0 1.2132e-08 0.0021 1.2135e-08 0 1.2189e-08 0 1.2192e-08 0.0021 1.2195e-08 0 1.2249e-08 0 1.2252e-08 0.0021 1.2255e-08 0 1.2309e-08 0 1.2312e-08 0.0021 1.2315e-08 0 1.2369e-08 0 1.2372e-08 0.0021 1.2375e-08 0 1.2429e-08 0 1.2432e-08 0.0021 1.2435e-08 0 1.2489e-08 0 1.2492e-08 0.0021 1.2495e-08 0 1.2549e-08 0 1.2552e-08 0.0021 1.2555e-08 0 1.2609e-08 0 1.2612e-08 0.0021 1.2615e-08 0 1.2669e-08 0 1.2672e-08 0.0021 1.2675e-08 0 1.2729e-08 0 1.2732e-08 0.0021 1.2735e-08 0 1.2789e-08 0 1.2792e-08 0.0021 1.2795e-08 0 1.2849e-08 0 1.2852e-08 0.0021 1.2855e-08 0 1.2909e-08 0 1.2912e-08 0.0021 1.2915e-08 0 1.2969e-08 0 1.2972e-08 0.0021 1.2975e-08 0 1.3029e-08 0 1.3032e-08 0.0021 1.3035e-08 0 1.3089e-08 0 1.3092e-08 0.0021 1.3095e-08 0 1.3149e-08 0 1.3152e-08 0.0021 1.3155e-08 0 1.3209e-08 0 1.3212e-08 0.0021 1.3215e-08 0 1.3269e-08 0 1.3272e-08 0.0021 1.3275e-08 0 1.3329e-08 0 1.3332e-08 0.0021 1.3335e-08 0 1.3389e-08 0 1.3392e-08 0.0021 1.3395e-08 0 1.3449e-08 0 1.3452e-08 0.0021 1.3455e-08 0 1.3509e-08 0 1.3512e-08 0.0021 1.3515e-08 0 1.3569e-08 0 1.3572e-08 0.0021 1.3575e-08 0 1.3629e-08 0 1.3632e-08 0.0021 1.3635e-08 0 1.3689e-08 0 1.3692e-08 0.0021 1.3695e-08 0 1.3749e-08 0 1.3752e-08 0.0021 1.3755e-08 0 1.3809e-08 0 1.3812e-08 0.0021 1.3815e-08 0 1.3869e-08 0 1.3872e-08 0.0021 1.3875e-08 0 1.3929e-08 0 1.3932e-08 0.0021 1.3935e-08 0 1.3989e-08 0 1.3992e-08 0.0021 1.3995e-08 0 1.4049e-08 0 1.4052e-08 0.0021 1.4055e-08 0 1.4109e-08 0 1.4112e-08 0.0021 1.4115e-08 0 1.4169e-08 0 1.4172e-08 0.0021 1.4175e-08 0 1.4229e-08 0 1.4232e-08 0.0021 1.4235e-08 0 1.4289e-08 0 1.4292e-08 0.0021 1.4295e-08 0 1.4349e-08 0 1.4352e-08 0.0021 1.4355e-08 0 1.4409e-08 0 1.4412e-08 0.0021 1.4415e-08 0 1.4469e-08 0 1.4472e-08 0.0021 1.4475e-08 0 1.4529e-08 0 1.4532e-08 0.0021 1.4535e-08 0 1.4589e-08 0 1.4592e-08 0.0021 1.4595e-08 0 1.4649e-08 0 1.4652e-08 0.0021 1.4655e-08 0 1.4709e-08 0 1.4712e-08 0.0021 1.4715e-08 0 1.4769e-08 0 1.4772e-08 0.0021 1.4775e-08 0 1.4829e-08 0 1.4832e-08 0.0021 1.4835e-08 0 1.4889e-08 0 1.4892e-08 0.0021 1.4895e-08 0 1.4949e-08 0 1.4952e-08 0.0021 1.4955e-08 0 1.5009e-08 0 1.5012e-08 0.0021 1.5015e-08 0 1.5069e-08 0 1.5072e-08 0.0021 1.5075e-08 0 1.5129e-08 0 1.5132e-08 0.0021 1.5135e-08 0 1.5189e-08 0 1.5192e-08 0.0021 1.5195e-08 0 1.5249e-08 0 1.5252e-08 0.0021 1.5255e-08 0 1.5309e-08 0 1.5312e-08 0.0021 1.5315e-08 0 1.5369e-08 0 1.5372e-08 0.0021 1.5375e-08 0 1.5429e-08 0 1.5432e-08 0.0021 1.5435e-08 0 1.5489e-08 0 1.5492e-08 0.0021 1.5495e-08 0 1.5549e-08 0 1.5552e-08 0.0021 1.5555e-08 0 1.5609e-08 0 1.5612e-08 0.0021 1.5615e-08 0 1.5669e-08 0 1.5672e-08 0.0021 1.5675e-08 0 1.5729e-08 0 1.5732e-08 0.0021 1.5735e-08 0 1.5789e-08 0 1.5792e-08 0.0021 1.5795e-08 0 1.5849e-08 0 1.5852e-08 0.0021 1.5855e-08 0 1.5909e-08 0 1.5912e-08 0.0021 1.5915e-08 0 1.5969e-08 0 1.5972e-08 0.0021 1.5975e-08 0 1.6029e-08 0 1.6032e-08 0.0021 1.6035e-08 0 1.6089e-08 0 1.6092e-08 0.0021 1.6095e-08 0 1.6149e-08 0 1.6152e-08 0.0021 1.6155e-08 0 1.6209e-08 0 1.6212e-08 0.0021 1.6215e-08 0 1.6269e-08 0 1.6272e-08 0.0021 1.6275e-08 0 1.6329e-08 0 1.6332e-08 0.0021 1.6335e-08 0 1.6389e-08 0 1.6392e-08 0.0021 1.6395e-08 0 1.6449e-08 0 1.6452e-08 0.0021 1.6455e-08 0 1.6509e-08 0 1.6512e-08 0.0021 1.6515e-08 0 1.6569e-08 0 1.6572e-08 0.0021 1.6575e-08 0 1.6629e-08 0 1.6632e-08 0.0021 1.6635e-08 0 1.6689e-08 0 1.6692e-08 0.0021 1.6695e-08 0 1.6749e-08 0 1.6752e-08 0.0021 1.6755e-08 0 1.6809e-08 0 1.6812e-08 0.0021 1.6815e-08 0 1.6869e-08 0 1.6872e-08 0.0021 1.6875e-08 0 1.6929e-08 0 1.6932e-08 0.0021 1.6935e-08 0 1.6989e-08 0 1.6992e-08 0.0021 1.6995e-08 0 1.7049e-08 0 1.7052e-08 0.0021 1.7055e-08 0 1.7109e-08 0 1.7112e-08 0.0021 1.7115e-08 0 1.7169e-08 0 1.7172e-08 0.0021 1.7175e-08 0 1.7229e-08 0 1.7232e-08 0.0021 1.7235e-08 0 1.7289e-08 0 1.7292e-08 0.0021 1.7295e-08 0 1.7349e-08 0 1.7352e-08 0.0021 1.7355e-08 0 1.7409e-08 0 1.7412e-08 0.0021 1.7415e-08 0 1.7469e-08 0 1.7472e-08 0.0021 1.7475e-08 0 1.7529e-08 0 1.7532e-08 0.0021 1.7535e-08 0 1.7589e-08 0 1.7592e-08 0.0021 1.7595e-08 0 1.7649e-08 0 1.7652e-08 0.0021 1.7655e-08 0 1.7709e-08 0 1.7712e-08 0.0021 1.7715e-08 0 1.7769e-08 0 1.7772e-08 0.0021 1.7775e-08 0 1.7829e-08 0 1.7832e-08 0.0021 1.7835e-08 0 1.7889e-08 0 1.7892e-08 0.0021 1.7895e-08 0 1.7949e-08 0 1.7952e-08 0.0021 1.7955e-08 0 1.8009e-08 0 1.8012e-08 0.0021 1.8015e-08 0 1.8069e-08 0 1.8072e-08 0.0021 1.8075e-08 0 1.8129e-08 0 1.8132e-08 0.0021 1.8135e-08 0 1.8189e-08 0 1.8192e-08 0.0021 1.8195e-08 0 1.8249e-08 0 1.8252e-08 0.0021 1.8255e-08 0 1.8309e-08 0 1.8312e-08 0.0021 1.8315e-08 0 1.8369e-08 0 1.8372e-08 0.0021 1.8375e-08 0 1.8429e-08 0 1.8432e-08 0.0021 1.8435e-08 0 1.8489e-08 0 1.8492e-08 0.0021 1.8495e-08 0 1.8549e-08 0 1.8552e-08 0.0021 1.8555e-08 0 1.8609e-08 0 1.8612e-08 0.0021 1.8615e-08 0 1.8669e-08 0 1.8672e-08 0.0021 1.8675e-08 0 1.8729e-08 0 1.8732e-08 0.0021 1.8735e-08 0 1.8789e-08 0 1.8792e-08 0.0021 1.8795e-08 0 1.8849e-08 0 1.8852e-08 0.0021 1.8855e-08 0 1.8909e-08 0 1.8912e-08 0.0021 1.8915e-08 0 1.8969e-08 0 1.8972e-08 0.0021 1.8975e-08 0 1.9029e-08 0 1.9032e-08 0.0021 1.9035e-08 0 1.9089e-08 0 1.9092e-08 0.0021 1.9095e-08 0 1.9149e-08 0 1.9152e-08 0.0021 1.9155e-08 0 1.9209e-08 0 1.9212e-08 0.0021 1.9215e-08 0 1.9269e-08 0 1.9272e-08 0.0021 1.9275e-08 0 1.9329e-08 0 1.9332e-08 0.0021 1.9335e-08 0 1.9389e-08 0 1.9392e-08 0.0021 1.9395e-08 0 1.9449e-08 0 1.9452e-08 0.0021 1.9455e-08 0 1.9509e-08 0 1.9512e-08 0.0021 1.9515e-08 0 1.9569e-08 0 1.9572e-08 0.0021 1.9575e-08 0 1.9629e-08 0 1.9632e-08 0.0021 1.9635e-08 0 1.9689e-08 0 1.9692e-08 0.0021 1.9695e-08 0 1.9749e-08 0 1.9752e-08 0.0021 1.9755e-08 0 1.9809e-08 0 1.9812e-08 0.0021 1.9815e-08 0 1.9869e-08 0 1.9872e-08 0.0021 1.9875e-08 0 1.9929e-08 0 1.9932e-08 0.0021 1.9935e-08 0 1.9989e-08 0 1.9992e-08 0.0021 1.9995e-08 0 2.0049e-08 0 2.0052e-08 0.0021 2.0055e-08 0 2.0109e-08 0 2.0112e-08 0.0021 2.0115e-08 0 2.0169e-08 0 2.0172e-08 0.0021 2.0175e-08 0 2.0229e-08 0 2.0232e-08 0.0021 2.0235e-08 0 2.0289e-08 0 2.0292e-08 0.0021 2.0295e-08 0 2.0349e-08 0 2.0352e-08 0.0021 2.0355e-08 0 2.0409e-08 0 2.0412e-08 0.0021 2.0415e-08 0 2.0469e-08 0 2.0472e-08 0.0021 2.0475e-08 0 2.0529e-08 0 2.0532e-08 0.0021 2.0535e-08 0 2.0589e-08 0 2.0592e-08 0.0021 2.0595e-08 0 2.0649e-08 0 2.0652e-08 0.0021 2.0655e-08 0 2.0709e-08 0 2.0712e-08 0.0021 2.0715e-08 0 2.0769e-08 0 2.0772e-08 0.0021 2.0775e-08 0 2.0829e-08 0 2.0832e-08 0.0021 2.0835e-08 0 2.0889e-08 0 2.0892e-08 0.0021 2.0895e-08 0 2.0949e-08 0 2.0952e-08 0.0021 2.0955e-08 0 2.1009e-08 0 2.1012e-08 0.0021 2.1015e-08 0 2.1069e-08 0 2.1072e-08 0.0021 2.1075e-08 0 2.1129e-08 0 2.1132e-08 0.0021 2.1135e-08 0 2.1189e-08 0 2.1192e-08 0.0021 2.1195e-08 0 2.1249e-08 0 2.1252e-08 0.0021 2.1255e-08 0 2.1309e-08 0 2.1312e-08 0.0021 2.1315e-08 0 2.1369e-08 0 2.1372e-08 0.0021 2.1375e-08 0 2.1429e-08 0 2.1432e-08 0.0021 2.1435e-08 0 2.1489e-08 0 2.1492e-08 0.0021 2.1495e-08 0 2.1549e-08 0 2.1552e-08 0.0021 2.1555e-08 0 2.1609e-08 0 2.1612e-08 0.0021 2.1615e-08 0 2.1669e-08 0 2.1672e-08 0.0021 2.1675e-08 0 2.1729e-08 0 2.1732e-08 0.0021 2.1735e-08 0 2.1789e-08 0 2.1792e-08 0.0021 2.1795e-08 0 2.1849e-08 0 2.1852e-08 0.0021 2.1855e-08 0 2.1909e-08 0 2.1912e-08 0.0021 2.1915e-08 0 2.1969e-08 0 2.1972e-08 0.0021 2.1975e-08 0 2.2029e-08 0 2.2032e-08 0.0021 2.2035e-08 0 2.2089e-08 0 2.2092e-08 0.0021 2.2095e-08 0 2.2149e-08 0 2.2152e-08 0.0021 2.2155e-08 0 2.2209e-08 0 2.2212e-08 0.0021 2.2215e-08 0 2.2269e-08 0 2.2272e-08 0.0021 2.2275e-08 0 2.2329e-08 0 2.2332e-08 0.0021 2.2335e-08 0 2.2389e-08 0 2.2392e-08 0.0021 2.2395e-08 0 2.2449e-08 0 2.2452e-08 0.0021 2.2455e-08 0 2.2509e-08 0 2.2512e-08 0.0021 2.2515e-08 0 2.2569e-08 0 2.2572e-08 0.0021 2.2575e-08 0 2.2629e-08 0 2.2632e-08 0.0021 2.2635e-08 0 2.2689e-08 0 2.2692e-08 0.0021 2.2695e-08 0 2.2749e-08 0 2.2752e-08 0.0021 2.2755e-08 0 2.2809e-08 0 2.2812e-08 0.0021 2.2815e-08 0 2.2869e-08 0 2.2872e-08 0.0021 2.2875e-08 0 2.2929e-08 0 2.2932e-08 0.0021 2.2935e-08 0 2.2989e-08 0 2.2992e-08 0.0021 2.2995e-08 0 2.3049e-08 0 2.3052e-08 0.0021 2.3055e-08 0 2.3109e-08 0 2.3112e-08 0.0021 2.3115e-08 0 2.3169e-08 0 2.3172e-08 0.0021 2.3175e-08 0 2.3229e-08 0 2.3232e-08 0.0021 2.3235e-08 0 2.3289e-08 0 2.3292e-08 0.0021 2.3295e-08 0 2.3349e-08 0 2.3352e-08 0.0021 2.3355e-08 0 2.3409e-08 0 2.3412e-08 0.0021 2.3415e-08 0 2.3469e-08 0 2.3472e-08 0.0021 2.3475e-08 0 2.3529e-08 0 2.3532e-08 0.0021 2.3535e-08 0 2.3589e-08 0 2.3592e-08 0.0021 2.3595e-08 0 2.3649e-08 0 2.3652e-08 0.0021 2.3655e-08 0 2.3709e-08 0 2.3712e-08 0.0021 2.3715e-08 0 2.3769e-08 0 2.3772e-08 0.0021 2.3775e-08 0 2.3829e-08 0 2.3832e-08 0.0021 2.3835e-08 0 2.3889e-08 0 2.3892e-08 0.0021 2.3895e-08 0)
IT03|T 0 T03  PWL(0 0 9e-12 0 1.2e-11 0.0021 1.5e-11 0 6.9e-11 0 7.2e-11 0.0021 7.5e-11 0 1.29e-10 0 1.32e-10 0.0021 1.35e-10 0 1.89e-10 0 1.92e-10 0.0021 1.95e-10 0 2.49e-10 0 2.52e-10 0.0021 2.55e-10 0 3.09e-10 0 3.12e-10 0.0021 3.15e-10 0 3.69e-10 0 3.72e-10 0.0021 3.75e-10 0 4.29e-10 0 4.32e-10 0.0021 4.35e-10 0 4.89e-10 0 4.92e-10 0.0021 4.95e-10 0 5.49e-10 0 5.52e-10 0.0021 5.55e-10 0 6.09e-10 0 6.12e-10 0.0021 6.15e-10 0 6.69e-10 0 6.72e-10 0.0021 6.75e-10 0 7.29e-10 0 7.32e-10 0.0021 7.35e-10 0 7.89e-10 0 7.92e-10 0.0021 7.95e-10 0 8.49e-10 0 8.52e-10 0.0021 8.55e-10 0 9.09e-10 0 9.12e-10 0.0021 9.15e-10 0 9.69e-10 0 9.72e-10 0.0021 9.75e-10 0 1.029e-09 0 1.032e-09 0.0021 1.035e-09 0 1.089e-09 0 1.092e-09 0.0021 1.095e-09 0 1.149e-09 0 1.152e-09 0.0021 1.155e-09 0 1.209e-09 0 1.212e-09 0.0021 1.215e-09 0 1.269e-09 0 1.272e-09 0.0021 1.275e-09 0 1.329e-09 0 1.332e-09 0.0021 1.335e-09 0 1.389e-09 0 1.392e-09 0.0021 1.395e-09 0 1.449e-09 0 1.452e-09 0.0021 1.455e-09 0 1.509e-09 0 1.512e-09 0.0021 1.515e-09 0 1.569e-09 0 1.572e-09 0.0021 1.575e-09 0 1.629e-09 0 1.632e-09 0.0021 1.635e-09 0 1.689e-09 0 1.692e-09 0.0021 1.695e-09 0 1.749e-09 0 1.752e-09 0.0021 1.755e-09 0 1.809e-09 0 1.812e-09 0.0021 1.815e-09 0 1.869e-09 0 1.872e-09 0.0021 1.875e-09 0 1.929e-09 0 1.932e-09 0.0021 1.935e-09 0 1.989e-09 0 1.992e-09 0.0021 1.995e-09 0 2.049e-09 0 2.052e-09 0.0021 2.055e-09 0 2.109e-09 0 2.112e-09 0.0021 2.115e-09 0 2.169e-09 0 2.172e-09 0.0021 2.175e-09 0 2.229e-09 0 2.232e-09 0.0021 2.235e-09 0 2.289e-09 0 2.292e-09 0.0021 2.295e-09 0 2.349e-09 0 2.352e-09 0.0021 2.355e-09 0 2.409e-09 0 2.412e-09 0.0021 2.415e-09 0 2.469e-09 0 2.472e-09 0.0021 2.475e-09 0 2.529e-09 0 2.532e-09 0.0021 2.535e-09 0 2.589e-09 0 2.592e-09 0.0021 2.595e-09 0 2.649e-09 0 2.652e-09 0.0021 2.655e-09 0 2.709e-09 0 2.712e-09 0.0021 2.715e-09 0 2.769e-09 0 2.772e-09 0.0021 2.775e-09 0 2.829e-09 0 2.832e-09 0.0021 2.835e-09 0 2.889e-09 0 2.892e-09 0.0021 2.895e-09 0 2.949e-09 0 2.952e-09 0.0021 2.955e-09 0 3.009e-09 0 3.012e-09 0.0021 3.015e-09 0 3.069e-09 0 3.072e-09 0.0021 3.075e-09 0 3.129e-09 0 3.132e-09 0.0021 3.135e-09 0 3.189e-09 0 3.192e-09 0.0021 3.195e-09 0 3.249e-09 0 3.252e-09 0.0021 3.255e-09 0 3.309e-09 0 3.312e-09 0.0021 3.315e-09 0 3.369e-09 0 3.372e-09 0.0021 3.375e-09 0 3.429e-09 0 3.432e-09 0.0021 3.435e-09 0 3.489e-09 0 3.492e-09 0.0021 3.495e-09 0 3.549e-09 0 3.552e-09 0.0021 3.555e-09 0 3.609e-09 0 3.612e-09 0.0021 3.615e-09 0 3.669e-09 0 3.672e-09 0.0021 3.675e-09 0 3.729e-09 0 3.732e-09 0.0021 3.735e-09 0 3.789e-09 0 3.792e-09 0.0021 3.795e-09 0 3.849e-09 0 3.852e-09 0.0021 3.855e-09 0 3.909e-09 0 3.912e-09 0.0021 3.915e-09 0 3.969e-09 0 3.972e-09 0.0021 3.975e-09 0 4.029e-09 0 4.032e-09 0.0021 4.035e-09 0 4.089e-09 0 4.092e-09 0.0021 4.095e-09 0 4.149e-09 0 4.152e-09 0.0021 4.155e-09 0 4.209e-09 0 4.212e-09 0.0021 4.215e-09 0 4.269e-09 0 4.272e-09 0.0021 4.275e-09 0 4.329e-09 0 4.332e-09 0.0021 4.335e-09 0 4.389e-09 0 4.392e-09 0.0021 4.395e-09 0 4.449e-09 0 4.452e-09 0.0021 4.455e-09 0 4.509e-09 0 4.512e-09 0.0021 4.515e-09 0 4.569e-09 0 4.572e-09 0.0021 4.575e-09 0 4.629e-09 0 4.632e-09 0.0021 4.635e-09 0 4.689e-09 0 4.692e-09 0.0021 4.695e-09 0 4.749e-09 0 4.752e-09 0.0021 4.755e-09 0 4.809e-09 0 4.812e-09 0.0021 4.815e-09 0 4.869e-09 0 4.872e-09 0.0021 4.875e-09 0 4.929e-09 0 4.932e-09 0.0021 4.935e-09 0 4.989e-09 0 4.992e-09 0.0021 4.995e-09 0 5.049e-09 0 5.052e-09 0.0021 5.055e-09 0 5.109e-09 0 5.112e-09 0.0021 5.115e-09 0 5.169e-09 0 5.172e-09 0.0021 5.175e-09 0 5.229e-09 0 5.232e-09 0.0021 5.235e-09 0 5.289e-09 0 5.292e-09 0.0021 5.295e-09 0 5.349e-09 0 5.352e-09 0.0021 5.355e-09 0 5.409e-09 0 5.412e-09 0.0021 5.415e-09 0 5.469e-09 0 5.472e-09 0.0021 5.475e-09 0 5.529e-09 0 5.532e-09 0.0021 5.535e-09 0 5.589e-09 0 5.592e-09 0.0021 5.595e-09 0 5.649e-09 0 5.652e-09 0.0021 5.655e-09 0 5.709e-09 0 5.712e-09 0.0021 5.715e-09 0 5.769e-09 0 5.772e-09 0.0021 5.775e-09 0 5.829e-09 0 5.832e-09 0.0021 5.835e-09 0 5.889e-09 0 5.892e-09 0.0021 5.895e-09 0 5.949e-09 0 5.952e-09 0.0021 5.955e-09 0 6.009e-09 0 6.012e-09 0.0021 6.015e-09 0 6.069e-09 0 6.072e-09 0.0021 6.075e-09 0 6.129e-09 0 6.132e-09 0.0021 6.135e-09 0 6.189e-09 0 6.192e-09 0.0021 6.195e-09 0 6.249e-09 0 6.252e-09 0.0021 6.255e-09 0 6.309e-09 0 6.312e-09 0.0021 6.315e-09 0 6.369e-09 0 6.372e-09 0.0021 6.375e-09 0 6.429e-09 0 6.432e-09 0.0021 6.435e-09 0 6.489e-09 0 6.492e-09 0.0021 6.495e-09 0 6.549e-09 0 6.552e-09 0.0021 6.555e-09 0 6.609e-09 0 6.612e-09 0.0021 6.615e-09 0 6.669e-09 0 6.672e-09 0.0021 6.675e-09 0 6.729e-09 0 6.732e-09 0.0021 6.735e-09 0 6.789e-09 0 6.792e-09 0.0021 6.795e-09 0 6.849e-09 0 6.852e-09 0.0021 6.855e-09 0 6.909e-09 0 6.912e-09 0.0021 6.915e-09 0 6.969e-09 0 6.972e-09 0.0021 6.975e-09 0 7.029e-09 0 7.032e-09 0.0021 7.035e-09 0 7.089e-09 0 7.092e-09 0.0021 7.095e-09 0 7.149e-09 0 7.152e-09 0.0021 7.155e-09 0 7.209e-09 0 7.212e-09 0.0021 7.215e-09 0 7.269e-09 0 7.272e-09 0.0021 7.275e-09 0 7.329e-09 0 7.332e-09 0.0021 7.335e-09 0 7.389e-09 0 7.392e-09 0.0021 7.395e-09 0 7.449e-09 0 7.452e-09 0.0021 7.455e-09 0 7.509e-09 0 7.512e-09 0.0021 7.515e-09 0 7.569e-09 0 7.572e-09 0.0021 7.575e-09 0 7.629e-09 0 7.632e-09 0.0021 7.635e-09 0 7.689e-09 0 7.692e-09 0.0021 7.695e-09 0 7.749e-09 0 7.752e-09 0.0021 7.755e-09 0 7.809e-09 0 7.812e-09 0.0021 7.815e-09 0 7.869e-09 0 7.872e-09 0.0021 7.875e-09 0 7.929e-09 0 7.932e-09 0.0021 7.935e-09 0 7.989e-09 0 7.992e-09 0.0021 7.995e-09 0 8.049e-09 0 8.052e-09 0.0021 8.055e-09 0 8.109e-09 0 8.112e-09 0.0021 8.115e-09 0 8.169e-09 0 8.172e-09 0.0021 8.175e-09 0 8.229e-09 0 8.232e-09 0.0021 8.235e-09 0 8.289e-09 0 8.292e-09 0.0021 8.295e-09 0 8.349e-09 0 8.352e-09 0.0021 8.355e-09 0 8.409e-09 0 8.412e-09 0.0021 8.415e-09 0 8.469e-09 0 8.472e-09 0.0021 8.475e-09 0 8.529e-09 0 8.532e-09 0.0021 8.535e-09 0 8.589e-09 0 8.592e-09 0.0021 8.595e-09 0 8.649e-09 0 8.652e-09 0.0021 8.655e-09 0 8.709e-09 0 8.712e-09 0.0021 8.715e-09 0 8.769e-09 0 8.772e-09 0.0021 8.775e-09 0 8.829e-09 0 8.832e-09 0.0021 8.835e-09 0 8.889e-09 0 8.892e-09 0.0021 8.895e-09 0 8.949e-09 0 8.952e-09 0.0021 8.955e-09 0 9.009e-09 0 9.012e-09 0.0021 9.015e-09 0 9.069e-09 0 9.072e-09 0.0021 9.075e-09 0 9.129e-09 0 9.132e-09 0.0021 9.135e-09 0 9.189e-09 0 9.192e-09 0.0021 9.195e-09 0 9.249e-09 0 9.252e-09 0.0021 9.255e-09 0 9.309e-09 0 9.312e-09 0.0021 9.315e-09 0 9.369e-09 0 9.372e-09 0.0021 9.375e-09 0 9.429e-09 0 9.432e-09 0.0021 9.435e-09 0 9.489e-09 0 9.492e-09 0.0021 9.495e-09 0 9.549e-09 0 9.552e-09 0.0021 9.555e-09 0 9.609e-09 0 9.612e-09 0.0021 9.615e-09 0 9.669e-09 0 9.672e-09 0.0021 9.675e-09 0 9.729e-09 0 9.732e-09 0.0021 9.735e-09 0 9.789e-09 0 9.792e-09 0.0021 9.795e-09 0 9.849e-09 0 9.852e-09 0.0021 9.855e-09 0 9.909e-09 0 9.912e-09 0.0021 9.915e-09 0 9.969e-09 0 9.972e-09 0.0021 9.975e-09 0 1.0029e-08 0 1.0032e-08 0.0021 1.0035e-08 0 1.0089e-08 0 1.0092e-08 0.0021 1.0095e-08 0 1.0149e-08 0 1.0152e-08 0.0021 1.0155e-08 0 1.0209e-08 0 1.0212e-08 0.0021 1.0215e-08 0 1.0269e-08 0 1.0272e-08 0.0021 1.0275e-08 0 1.0329e-08 0 1.0332e-08 0.0021 1.0335e-08 0 1.0389e-08 0 1.0392e-08 0.0021 1.0395e-08 0 1.0449e-08 0 1.0452e-08 0.0021 1.0455e-08 0 1.0509e-08 0 1.0512e-08 0.0021 1.0515e-08 0 1.0569e-08 0 1.0572e-08 0.0021 1.0575e-08 0 1.0629e-08 0 1.0632e-08 0.0021 1.0635e-08 0 1.0689e-08 0 1.0692e-08 0.0021 1.0695e-08 0 1.0749e-08 0 1.0752e-08 0.0021 1.0755e-08 0 1.0809e-08 0 1.0812e-08 0.0021 1.0815e-08 0 1.0869e-08 0 1.0872e-08 0.0021 1.0875e-08 0 1.0929e-08 0 1.0932e-08 0.0021 1.0935e-08 0 1.0989e-08 0 1.0992e-08 0.0021 1.0995e-08 0 1.1049e-08 0 1.1052e-08 0.0021 1.1055e-08 0 1.1109e-08 0 1.1112e-08 0.0021 1.1115e-08 0 1.1169e-08 0 1.1172e-08 0.0021 1.1175e-08 0 1.1229e-08 0 1.1232e-08 0.0021 1.1235e-08 0 1.1289e-08 0 1.1292e-08 0.0021 1.1295e-08 0 1.1349e-08 0 1.1352e-08 0.0021 1.1355e-08 0 1.1409e-08 0 1.1412e-08 0.0021 1.1415e-08 0 1.1469e-08 0 1.1472e-08 0.0021 1.1475e-08 0 1.1529e-08 0 1.1532e-08 0.0021 1.1535e-08 0 1.1589e-08 0 1.1592e-08 0.0021 1.1595e-08 0 1.1649e-08 0 1.1652e-08 0.0021 1.1655e-08 0 1.1709e-08 0 1.1712e-08 0.0021 1.1715e-08 0 1.1769e-08 0 1.1772e-08 0.0021 1.1775e-08 0 1.1829e-08 0 1.1832e-08 0.0021 1.1835e-08 0 1.1889e-08 0 1.1892e-08 0.0021 1.1895e-08 0 1.1949e-08 0 1.1952e-08 0.0021 1.1955e-08 0 1.2009e-08 0 1.2012e-08 0.0021 1.2015e-08 0 1.2069e-08 0 1.2072e-08 0.0021 1.2075e-08 0 1.2129e-08 0 1.2132e-08 0.0021 1.2135e-08 0 1.2189e-08 0 1.2192e-08 0.0021 1.2195e-08 0 1.2249e-08 0 1.2252e-08 0.0021 1.2255e-08 0 1.2309e-08 0 1.2312e-08 0.0021 1.2315e-08 0 1.2369e-08 0 1.2372e-08 0.0021 1.2375e-08 0 1.2429e-08 0 1.2432e-08 0.0021 1.2435e-08 0 1.2489e-08 0 1.2492e-08 0.0021 1.2495e-08 0 1.2549e-08 0 1.2552e-08 0.0021 1.2555e-08 0 1.2609e-08 0 1.2612e-08 0.0021 1.2615e-08 0 1.2669e-08 0 1.2672e-08 0.0021 1.2675e-08 0 1.2729e-08 0 1.2732e-08 0.0021 1.2735e-08 0 1.2789e-08 0 1.2792e-08 0.0021 1.2795e-08 0 1.2849e-08 0 1.2852e-08 0.0021 1.2855e-08 0 1.2909e-08 0 1.2912e-08 0.0021 1.2915e-08 0 1.2969e-08 0 1.2972e-08 0.0021 1.2975e-08 0 1.3029e-08 0 1.3032e-08 0.0021 1.3035e-08 0 1.3089e-08 0 1.3092e-08 0.0021 1.3095e-08 0 1.3149e-08 0 1.3152e-08 0.0021 1.3155e-08 0 1.3209e-08 0 1.3212e-08 0.0021 1.3215e-08 0 1.3269e-08 0 1.3272e-08 0.0021 1.3275e-08 0 1.3329e-08 0 1.3332e-08 0.0021 1.3335e-08 0 1.3389e-08 0 1.3392e-08 0.0021 1.3395e-08 0 1.3449e-08 0 1.3452e-08 0.0021 1.3455e-08 0 1.3509e-08 0 1.3512e-08 0.0021 1.3515e-08 0 1.3569e-08 0 1.3572e-08 0.0021 1.3575e-08 0 1.3629e-08 0 1.3632e-08 0.0021 1.3635e-08 0 1.3689e-08 0 1.3692e-08 0.0021 1.3695e-08 0 1.3749e-08 0 1.3752e-08 0.0021 1.3755e-08 0 1.3809e-08 0 1.3812e-08 0.0021 1.3815e-08 0 1.3869e-08 0 1.3872e-08 0.0021 1.3875e-08 0 1.3929e-08 0 1.3932e-08 0.0021 1.3935e-08 0 1.3989e-08 0 1.3992e-08 0.0021 1.3995e-08 0 1.4049e-08 0 1.4052e-08 0.0021 1.4055e-08 0 1.4109e-08 0 1.4112e-08 0.0021 1.4115e-08 0 1.4169e-08 0 1.4172e-08 0.0021 1.4175e-08 0 1.4229e-08 0 1.4232e-08 0.0021 1.4235e-08 0 1.4289e-08 0 1.4292e-08 0.0021 1.4295e-08 0 1.4349e-08 0 1.4352e-08 0.0021 1.4355e-08 0 1.4409e-08 0 1.4412e-08 0.0021 1.4415e-08 0 1.4469e-08 0 1.4472e-08 0.0021 1.4475e-08 0 1.4529e-08 0 1.4532e-08 0.0021 1.4535e-08 0 1.4589e-08 0 1.4592e-08 0.0021 1.4595e-08 0 1.4649e-08 0 1.4652e-08 0.0021 1.4655e-08 0 1.4709e-08 0 1.4712e-08 0.0021 1.4715e-08 0 1.4769e-08 0 1.4772e-08 0.0021 1.4775e-08 0 1.4829e-08 0 1.4832e-08 0.0021 1.4835e-08 0 1.4889e-08 0 1.4892e-08 0.0021 1.4895e-08 0 1.4949e-08 0 1.4952e-08 0.0021 1.4955e-08 0 1.5009e-08 0 1.5012e-08 0.0021 1.5015e-08 0 1.5069e-08 0 1.5072e-08 0.0021 1.5075e-08 0 1.5129e-08 0 1.5132e-08 0.0021 1.5135e-08 0 1.5189e-08 0 1.5192e-08 0.0021 1.5195e-08 0 1.5249e-08 0 1.5252e-08 0.0021 1.5255e-08 0 1.5309e-08 0 1.5312e-08 0.0021 1.5315e-08 0 1.5369e-08 0 1.5372e-08 0.0021 1.5375e-08 0 1.5429e-08 0 1.5432e-08 0.0021 1.5435e-08 0 1.5489e-08 0 1.5492e-08 0.0021 1.5495e-08 0 1.5549e-08 0 1.5552e-08 0.0021 1.5555e-08 0 1.5609e-08 0 1.5612e-08 0.0021 1.5615e-08 0 1.5669e-08 0 1.5672e-08 0.0021 1.5675e-08 0 1.5729e-08 0 1.5732e-08 0.0021 1.5735e-08 0 1.5789e-08 0 1.5792e-08 0.0021 1.5795e-08 0 1.5849e-08 0 1.5852e-08 0.0021 1.5855e-08 0 1.5909e-08 0 1.5912e-08 0.0021 1.5915e-08 0 1.5969e-08 0 1.5972e-08 0.0021 1.5975e-08 0 1.6029e-08 0 1.6032e-08 0.0021 1.6035e-08 0 1.6089e-08 0 1.6092e-08 0.0021 1.6095e-08 0 1.6149e-08 0 1.6152e-08 0.0021 1.6155e-08 0 1.6209e-08 0 1.6212e-08 0.0021 1.6215e-08 0 1.6269e-08 0 1.6272e-08 0.0021 1.6275e-08 0 1.6329e-08 0 1.6332e-08 0.0021 1.6335e-08 0 1.6389e-08 0 1.6392e-08 0.0021 1.6395e-08 0 1.6449e-08 0 1.6452e-08 0.0021 1.6455e-08 0 1.6509e-08 0 1.6512e-08 0.0021 1.6515e-08 0 1.6569e-08 0 1.6572e-08 0.0021 1.6575e-08 0 1.6629e-08 0 1.6632e-08 0.0021 1.6635e-08 0 1.6689e-08 0 1.6692e-08 0.0021 1.6695e-08 0 1.6749e-08 0 1.6752e-08 0.0021 1.6755e-08 0 1.6809e-08 0 1.6812e-08 0.0021 1.6815e-08 0 1.6869e-08 0 1.6872e-08 0.0021 1.6875e-08 0 1.6929e-08 0 1.6932e-08 0.0021 1.6935e-08 0 1.6989e-08 0 1.6992e-08 0.0021 1.6995e-08 0 1.7049e-08 0 1.7052e-08 0.0021 1.7055e-08 0 1.7109e-08 0 1.7112e-08 0.0021 1.7115e-08 0 1.7169e-08 0 1.7172e-08 0.0021 1.7175e-08 0 1.7229e-08 0 1.7232e-08 0.0021 1.7235e-08 0 1.7289e-08 0 1.7292e-08 0.0021 1.7295e-08 0 1.7349e-08 0 1.7352e-08 0.0021 1.7355e-08 0 1.7409e-08 0 1.7412e-08 0.0021 1.7415e-08 0 1.7469e-08 0 1.7472e-08 0.0021 1.7475e-08 0 1.7529e-08 0 1.7532e-08 0.0021 1.7535e-08 0 1.7589e-08 0 1.7592e-08 0.0021 1.7595e-08 0 1.7649e-08 0 1.7652e-08 0.0021 1.7655e-08 0 1.7709e-08 0 1.7712e-08 0.0021 1.7715e-08 0 1.7769e-08 0 1.7772e-08 0.0021 1.7775e-08 0 1.7829e-08 0 1.7832e-08 0.0021 1.7835e-08 0 1.7889e-08 0 1.7892e-08 0.0021 1.7895e-08 0 1.7949e-08 0 1.7952e-08 0.0021 1.7955e-08 0 1.8009e-08 0 1.8012e-08 0.0021 1.8015e-08 0 1.8069e-08 0 1.8072e-08 0.0021 1.8075e-08 0 1.8129e-08 0 1.8132e-08 0.0021 1.8135e-08 0 1.8189e-08 0 1.8192e-08 0.0021 1.8195e-08 0 1.8249e-08 0 1.8252e-08 0.0021 1.8255e-08 0 1.8309e-08 0 1.8312e-08 0.0021 1.8315e-08 0 1.8369e-08 0 1.8372e-08 0.0021 1.8375e-08 0 1.8429e-08 0 1.8432e-08 0.0021 1.8435e-08 0 1.8489e-08 0 1.8492e-08 0.0021 1.8495e-08 0 1.8549e-08 0 1.8552e-08 0.0021 1.8555e-08 0 1.8609e-08 0 1.8612e-08 0.0021 1.8615e-08 0 1.8669e-08 0 1.8672e-08 0.0021 1.8675e-08 0 1.8729e-08 0 1.8732e-08 0.0021 1.8735e-08 0 1.8789e-08 0 1.8792e-08 0.0021 1.8795e-08 0 1.8849e-08 0 1.8852e-08 0.0021 1.8855e-08 0 1.8909e-08 0 1.8912e-08 0.0021 1.8915e-08 0 1.8969e-08 0 1.8972e-08 0.0021 1.8975e-08 0 1.9029e-08 0 1.9032e-08 0.0021 1.9035e-08 0 1.9089e-08 0 1.9092e-08 0.0021 1.9095e-08 0 1.9149e-08 0 1.9152e-08 0.0021 1.9155e-08 0 1.9209e-08 0 1.9212e-08 0.0021 1.9215e-08 0 1.9269e-08 0 1.9272e-08 0.0021 1.9275e-08 0 1.9329e-08 0 1.9332e-08 0.0021 1.9335e-08 0 1.9389e-08 0 1.9392e-08 0.0021 1.9395e-08 0 1.9449e-08 0 1.9452e-08 0.0021 1.9455e-08 0 1.9509e-08 0 1.9512e-08 0.0021 1.9515e-08 0 1.9569e-08 0 1.9572e-08 0.0021 1.9575e-08 0 1.9629e-08 0 1.9632e-08 0.0021 1.9635e-08 0 1.9689e-08 0 1.9692e-08 0.0021 1.9695e-08 0 1.9749e-08 0 1.9752e-08 0.0021 1.9755e-08 0 1.9809e-08 0 1.9812e-08 0.0021 1.9815e-08 0 1.9869e-08 0 1.9872e-08 0.0021 1.9875e-08 0 1.9929e-08 0 1.9932e-08 0.0021 1.9935e-08 0 1.9989e-08 0 1.9992e-08 0.0021 1.9995e-08 0 2.0049e-08 0 2.0052e-08 0.0021 2.0055e-08 0 2.0109e-08 0 2.0112e-08 0.0021 2.0115e-08 0 2.0169e-08 0 2.0172e-08 0.0021 2.0175e-08 0 2.0229e-08 0 2.0232e-08 0.0021 2.0235e-08 0 2.0289e-08 0 2.0292e-08 0.0021 2.0295e-08 0 2.0349e-08 0 2.0352e-08 0.0021 2.0355e-08 0 2.0409e-08 0 2.0412e-08 0.0021 2.0415e-08 0 2.0469e-08 0 2.0472e-08 0.0021 2.0475e-08 0 2.0529e-08 0 2.0532e-08 0.0021 2.0535e-08 0 2.0589e-08 0 2.0592e-08 0.0021 2.0595e-08 0 2.0649e-08 0 2.0652e-08 0.0021 2.0655e-08 0 2.0709e-08 0 2.0712e-08 0.0021 2.0715e-08 0 2.0769e-08 0 2.0772e-08 0.0021 2.0775e-08 0 2.0829e-08 0 2.0832e-08 0.0021 2.0835e-08 0 2.0889e-08 0 2.0892e-08 0.0021 2.0895e-08 0 2.0949e-08 0 2.0952e-08 0.0021 2.0955e-08 0 2.1009e-08 0 2.1012e-08 0.0021 2.1015e-08 0 2.1069e-08 0 2.1072e-08 0.0021 2.1075e-08 0 2.1129e-08 0 2.1132e-08 0.0021 2.1135e-08 0 2.1189e-08 0 2.1192e-08 0.0021 2.1195e-08 0 2.1249e-08 0 2.1252e-08 0.0021 2.1255e-08 0 2.1309e-08 0 2.1312e-08 0.0021 2.1315e-08 0 2.1369e-08 0 2.1372e-08 0.0021 2.1375e-08 0 2.1429e-08 0 2.1432e-08 0.0021 2.1435e-08 0 2.1489e-08 0 2.1492e-08 0.0021 2.1495e-08 0 2.1549e-08 0 2.1552e-08 0.0021 2.1555e-08 0 2.1609e-08 0 2.1612e-08 0.0021 2.1615e-08 0 2.1669e-08 0 2.1672e-08 0.0021 2.1675e-08 0 2.1729e-08 0 2.1732e-08 0.0021 2.1735e-08 0 2.1789e-08 0 2.1792e-08 0.0021 2.1795e-08 0 2.1849e-08 0 2.1852e-08 0.0021 2.1855e-08 0 2.1909e-08 0 2.1912e-08 0.0021 2.1915e-08 0 2.1969e-08 0 2.1972e-08 0.0021 2.1975e-08 0 2.2029e-08 0 2.2032e-08 0.0021 2.2035e-08 0 2.2089e-08 0 2.2092e-08 0.0021 2.2095e-08 0 2.2149e-08 0 2.2152e-08 0.0021 2.2155e-08 0 2.2209e-08 0 2.2212e-08 0.0021 2.2215e-08 0 2.2269e-08 0 2.2272e-08 0.0021 2.2275e-08 0 2.2329e-08 0 2.2332e-08 0.0021 2.2335e-08 0 2.2389e-08 0 2.2392e-08 0.0021 2.2395e-08 0 2.2449e-08 0 2.2452e-08 0.0021 2.2455e-08 0 2.2509e-08 0 2.2512e-08 0.0021 2.2515e-08 0 2.2569e-08 0 2.2572e-08 0.0021 2.2575e-08 0 2.2629e-08 0 2.2632e-08 0.0021 2.2635e-08 0 2.2689e-08 0 2.2692e-08 0.0021 2.2695e-08 0 2.2749e-08 0 2.2752e-08 0.0021 2.2755e-08 0 2.2809e-08 0 2.2812e-08 0.0021 2.2815e-08 0 2.2869e-08 0 2.2872e-08 0.0021 2.2875e-08 0 2.2929e-08 0 2.2932e-08 0.0021 2.2935e-08 0 2.2989e-08 0 2.2992e-08 0.0021 2.2995e-08 0 2.3049e-08 0 2.3052e-08 0.0021 2.3055e-08 0 2.3109e-08 0 2.3112e-08 0.0021 2.3115e-08 0 2.3169e-08 0 2.3172e-08 0.0021 2.3175e-08 0 2.3229e-08 0 2.3232e-08 0.0021 2.3235e-08 0 2.3289e-08 0 2.3292e-08 0.0021 2.3295e-08 0 2.3349e-08 0 2.3352e-08 0.0021 2.3355e-08 0 2.3409e-08 0 2.3412e-08 0.0021 2.3415e-08 0 2.3469e-08 0 2.3472e-08 0.0021 2.3475e-08 0 2.3529e-08 0 2.3532e-08 0.0021 2.3535e-08 0 2.3589e-08 0 2.3592e-08 0.0021 2.3595e-08 0 2.3649e-08 0 2.3652e-08 0.0021 2.3655e-08 0 2.3709e-08 0 2.3712e-08 0.0021 2.3715e-08 0 2.3769e-08 0 2.3772e-08 0.0021 2.3775e-08 0 2.3829e-08 0 2.3832e-08 0.0021 2.3835e-08 0 2.3889e-08 0 2.3892e-08 0.0021 2.3895e-08 0)
LSPL_IG0_0|1 IG0_0_RX SPL_IG0_0|D1  2e-12
LSPL_IG0_0|2 SPL_IG0_0|D1 SPL_IG0_0|D2  4.135667696e-12
LSPL_IG0_0|3 SPL_IG0_0|D2 SPL_IG0_0|JCT  9.84682784761905e-13
LSPL_IG0_0|4 SPL_IG0_0|JCT SPL_IG0_0|QA1  9.84682784761905e-13
LSPL_IG0_0|5 SPL_IG0_0|QA1 IG0_0_TO0  2e-12
LSPL_IG0_0|6 SPL_IG0_0|JCT SPL_IG0_0|QB1  9.84682784761905e-13
LSPL_IG0_0|7 SPL_IG0_0|QB1 IG0_0_TO1  2e-12
LSPL_IP1_0|1 IP1_0_RX SPL_IP1_0|D1  2e-12
LSPL_IP1_0|2 SPL_IP1_0|D1 SPL_IP1_0|D2  4.135667696e-12
LSPL_IP1_0|3 SPL_IP1_0|D2 SPL_IP1_0|JCT  9.84682784761905e-13
LSPL_IP1_0|4 SPL_IP1_0|JCT SPL_IP1_0|QA1  9.84682784761905e-13
LSPL_IP1_0|5 SPL_IP1_0|QA1 IP1_0_TO1  2e-12
LSPL_IP1_0|6 SPL_IP1_0|JCT SPL_IP1_0|QB1  9.84682784761905e-13
LSPL_IP1_0|7 SPL_IP1_0|QB1 IP1_0_OUT  2e-12
LSPL_IG2_0|1 IG2_0_RX SPL_IG2_0|D1  2e-12
LSPL_IG2_0|2 SPL_IG2_0|D1 SPL_IG2_0|D2  4.135667696e-12
LSPL_IG2_0|3 SPL_IG2_0|D2 SPL_IG2_0|JCT  9.84682784761905e-13
LSPL_IG2_0|4 SPL_IG2_0|JCT SPL_IG2_0|QA1  9.84682784761905e-13
LSPL_IG2_0|5 SPL_IG2_0|QA1 IG2_0_TO2  2e-12
LSPL_IG2_0|6 SPL_IG2_0|JCT SPL_IG2_0|QB1  9.84682784761905e-13
LSPL_IG2_0|7 SPL_IG2_0|QB1 IG2_0_TO3  2e-12
LSPL_IP3_0|1 IP3_0_RX SPL_IP3_0|D1  2e-12
LSPL_IP3_0|2 SPL_IP3_0|D1 SPL_IP3_0|D2  4.135667696e-12
LSPL_IP3_0|3 SPL_IP3_0|D2 SPL_IP3_0|JCT  9.84682784761905e-13
LSPL_IP3_0|4 SPL_IP3_0|JCT SPL_IP3_0|QA1  9.84682784761905e-13
LSPL_IP3_0|5 SPL_IP3_0|QA1 IP3_0_TO1  2e-12
LSPL_IP3_0|6 SPL_IP3_0|JCT SPL_IP3_0|QB1  9.84682784761905e-13
LSPL_IP3_0|7 SPL_IP3_0|QB1 IP3_0_OUT  2e-12
IT04|T 0 T04  PWL(0 0 6e-12 0 9e-12 0.0014 1.2e-11 0 6.6e-11 0 6.9e-11 0.0014 7.2e-11 0 1.26e-10 0 1.29e-10 0.0014 1.32e-10 0 1.86e-10 0 1.89e-10 0.0014 1.92e-10 0 2.46e-10 0 2.49e-10 0.0014 2.52e-10 0 3.06e-10 0 3.09e-10 0.0014 3.12e-10 0 3.66e-10 0 3.69e-10 0.0014 3.72e-10 0 4.26e-10 0 4.29e-10 0.0014 4.32e-10 0 4.86e-10 0 4.89e-10 0.0014 4.92e-10 0 5.46e-10 0 5.49e-10 0.0014 5.52e-10 0 6.06e-10 0 6.09e-10 0.0014 6.12e-10 0 6.66e-10 0 6.69e-10 0.0014 6.72e-10 0 7.26e-10 0 7.29e-10 0.0014 7.32e-10 0 7.86e-10 0 7.89e-10 0.0014 7.92e-10 0 8.46e-10 0 8.49e-10 0.0014 8.52e-10 0 9.06e-10 0 9.09e-10 0.0014 9.12e-10 0 9.66e-10 0 9.69e-10 0.0014 9.72e-10 0 1.026e-09 0 1.029e-09 0.0014 1.032e-09 0 1.086e-09 0 1.089e-09 0.0014 1.092e-09 0 1.146e-09 0 1.149e-09 0.0014 1.152e-09 0 1.206e-09 0 1.209e-09 0.0014 1.212e-09 0 1.266e-09 0 1.269e-09 0.0014 1.272e-09 0 1.326e-09 0 1.329e-09 0.0014 1.332e-09 0 1.386e-09 0 1.389e-09 0.0014 1.392e-09 0 1.446e-09 0 1.449e-09 0.0014 1.452e-09 0 1.506e-09 0 1.509e-09 0.0014 1.512e-09 0 1.566e-09 0 1.569e-09 0.0014 1.572e-09 0 1.626e-09 0 1.629e-09 0.0014 1.632e-09 0 1.686e-09 0 1.689e-09 0.0014 1.692e-09 0 1.746e-09 0 1.749e-09 0.0014 1.752e-09 0 1.806e-09 0 1.809e-09 0.0014 1.812e-09 0 1.866e-09 0 1.869e-09 0.0014 1.872e-09 0 1.926e-09 0 1.929e-09 0.0014 1.932e-09 0 1.986e-09 0 1.989e-09 0.0014 1.992e-09 0 2.046e-09 0 2.049e-09 0.0014 2.052e-09 0 2.106e-09 0 2.109e-09 0.0014 2.112e-09 0 2.166e-09 0 2.169e-09 0.0014 2.172e-09 0 2.226e-09 0 2.229e-09 0.0014 2.232e-09 0 2.286e-09 0 2.289e-09 0.0014 2.292e-09 0 2.346e-09 0 2.349e-09 0.0014 2.352e-09 0 2.406e-09 0 2.409e-09 0.0014 2.412e-09 0 2.466e-09 0 2.469e-09 0.0014 2.472e-09 0 2.526e-09 0 2.529e-09 0.0014 2.532e-09 0 2.586e-09 0 2.589e-09 0.0014 2.592e-09 0 2.646e-09 0 2.649e-09 0.0014 2.652e-09 0 2.706e-09 0 2.709e-09 0.0014 2.712e-09 0 2.766e-09 0 2.769e-09 0.0014 2.772e-09 0 2.826e-09 0 2.829e-09 0.0014 2.832e-09 0 2.886e-09 0 2.889e-09 0.0014 2.892e-09 0 2.946e-09 0 2.949e-09 0.0014 2.952e-09 0 3.006e-09 0 3.009e-09 0.0014 3.012e-09 0 3.066e-09 0 3.069e-09 0.0014 3.072e-09 0 3.126e-09 0 3.129e-09 0.0014 3.132e-09 0 3.186e-09 0 3.189e-09 0.0014 3.192e-09 0 3.246e-09 0 3.249e-09 0.0014 3.252e-09 0 3.306e-09 0 3.309e-09 0.0014 3.312e-09 0 3.366e-09 0 3.369e-09 0.0014 3.372e-09 0 3.426e-09 0 3.429e-09 0.0014 3.432e-09 0 3.486e-09 0 3.489e-09 0.0014 3.492e-09 0 3.546e-09 0 3.549e-09 0.0014 3.552e-09 0 3.606e-09 0 3.609e-09 0.0014 3.612e-09 0 3.666e-09 0 3.669e-09 0.0014 3.672e-09 0 3.726e-09 0 3.729e-09 0.0014 3.732e-09 0 3.786e-09 0 3.789e-09 0.0014 3.792e-09 0 3.846e-09 0 3.849e-09 0.0014 3.852e-09 0 3.906e-09 0 3.909e-09 0.0014 3.912e-09 0 3.966e-09 0 3.969e-09 0.0014 3.972e-09 0 4.026e-09 0 4.029e-09 0.0014 4.032e-09 0 4.086e-09 0 4.089e-09 0.0014 4.092e-09 0 4.146e-09 0 4.149e-09 0.0014 4.152e-09 0 4.206e-09 0 4.209e-09 0.0014 4.212e-09 0 4.266e-09 0 4.269e-09 0.0014 4.272e-09 0 4.326e-09 0 4.329e-09 0.0014 4.332e-09 0 4.386e-09 0 4.389e-09 0.0014 4.392e-09 0 4.446e-09 0 4.449e-09 0.0014 4.452e-09 0 4.506e-09 0 4.509e-09 0.0014 4.512e-09 0 4.566e-09 0 4.569e-09 0.0014 4.572e-09 0 4.626e-09 0 4.629e-09 0.0014 4.632e-09 0 4.686e-09 0 4.689e-09 0.0014 4.692e-09 0 4.746e-09 0 4.749e-09 0.0014 4.752e-09 0 4.806e-09 0 4.809e-09 0.0014 4.812e-09 0 4.866e-09 0 4.869e-09 0.0014 4.872e-09 0 4.926e-09 0 4.929e-09 0.0014 4.932e-09 0 4.986e-09 0 4.989e-09 0.0014 4.992e-09 0 5.046e-09 0 5.049e-09 0.0014 5.052e-09 0 5.106e-09 0 5.109e-09 0.0014 5.112e-09 0 5.166e-09 0 5.169e-09 0.0014 5.172e-09 0 5.226e-09 0 5.229e-09 0.0014 5.232e-09 0 5.286e-09 0 5.289e-09 0.0014 5.292e-09 0 5.346e-09 0 5.349e-09 0.0014 5.352e-09 0 5.406e-09 0 5.409e-09 0.0014 5.412e-09 0 5.466e-09 0 5.469e-09 0.0014 5.472e-09 0 5.526e-09 0 5.529e-09 0.0014 5.532e-09 0 5.586e-09 0 5.589e-09 0.0014 5.592e-09 0 5.646e-09 0 5.649e-09 0.0014 5.652e-09 0 5.706e-09 0 5.709e-09 0.0014 5.712e-09 0 5.766e-09 0 5.769e-09 0.0014 5.772e-09 0 5.826e-09 0 5.829e-09 0.0014 5.832e-09 0 5.886e-09 0 5.889e-09 0.0014 5.892e-09 0 5.946e-09 0 5.949e-09 0.0014 5.952e-09 0 6.006e-09 0 6.009e-09 0.0014 6.012e-09 0 6.066e-09 0 6.069e-09 0.0014 6.072e-09 0 6.126e-09 0 6.129e-09 0.0014 6.132e-09 0 6.186e-09 0 6.189e-09 0.0014 6.192e-09 0 6.246e-09 0 6.249e-09 0.0014 6.252e-09 0 6.306e-09 0 6.309e-09 0.0014 6.312e-09 0 6.366e-09 0 6.369e-09 0.0014 6.372e-09 0 6.426e-09 0 6.429e-09 0.0014 6.432e-09 0 6.486e-09 0 6.489e-09 0.0014 6.492e-09 0 6.546e-09 0 6.549e-09 0.0014 6.552e-09 0 6.606e-09 0 6.609e-09 0.0014 6.612e-09 0 6.666e-09 0 6.669e-09 0.0014 6.672e-09 0 6.726e-09 0 6.729e-09 0.0014 6.732e-09 0 6.786e-09 0 6.789e-09 0.0014 6.792e-09 0 6.846e-09 0 6.849e-09 0.0014 6.852e-09 0 6.906e-09 0 6.909e-09 0.0014 6.912e-09 0 6.966e-09 0 6.969e-09 0.0014 6.972e-09 0 7.026e-09 0 7.029e-09 0.0014 7.032e-09 0 7.086e-09 0 7.089e-09 0.0014 7.092e-09 0 7.146e-09 0 7.149e-09 0.0014 7.152e-09 0 7.206e-09 0 7.209e-09 0.0014 7.212e-09 0 7.266e-09 0 7.269e-09 0.0014 7.272e-09 0 7.326e-09 0 7.329e-09 0.0014 7.332e-09 0 7.386e-09 0 7.389e-09 0.0014 7.392e-09 0 7.446e-09 0 7.449e-09 0.0014 7.452e-09 0 7.506e-09 0 7.509e-09 0.0014 7.512e-09 0 7.566e-09 0 7.569e-09 0.0014 7.572e-09 0 7.626e-09 0 7.629e-09 0.0014 7.632e-09 0 7.686e-09 0 7.689e-09 0.0014 7.692e-09 0 7.746e-09 0 7.749e-09 0.0014 7.752e-09 0 7.806e-09 0 7.809e-09 0.0014 7.812e-09 0 7.866e-09 0 7.869e-09 0.0014 7.872e-09 0 7.926e-09 0 7.929e-09 0.0014 7.932e-09 0 7.986e-09 0 7.989e-09 0.0014 7.992e-09 0 8.046e-09 0 8.049e-09 0.0014 8.052e-09 0 8.106e-09 0 8.109e-09 0.0014 8.112e-09 0 8.166e-09 0 8.169e-09 0.0014 8.172e-09 0 8.226e-09 0 8.229e-09 0.0014 8.232e-09 0 8.286e-09 0 8.289e-09 0.0014 8.292e-09 0 8.346e-09 0 8.349e-09 0.0014 8.352e-09 0 8.406e-09 0 8.409e-09 0.0014 8.412e-09 0 8.466e-09 0 8.469e-09 0.0014 8.472e-09 0 8.526e-09 0 8.529e-09 0.0014 8.532e-09 0 8.586e-09 0 8.589e-09 0.0014 8.592e-09 0 8.646e-09 0 8.649e-09 0.0014 8.652e-09 0 8.706e-09 0 8.709e-09 0.0014 8.712e-09 0 8.766e-09 0 8.769e-09 0.0014 8.772e-09 0 8.826e-09 0 8.829e-09 0.0014 8.832e-09 0 8.886e-09 0 8.889e-09 0.0014 8.892e-09 0 8.946e-09 0 8.949e-09 0.0014 8.952e-09 0 9.006e-09 0 9.009e-09 0.0014 9.012e-09 0 9.066e-09 0 9.069e-09 0.0014 9.072e-09 0 9.126e-09 0 9.129e-09 0.0014 9.132e-09 0 9.186e-09 0 9.189e-09 0.0014 9.192e-09 0 9.246e-09 0 9.249e-09 0.0014 9.252e-09 0 9.306e-09 0 9.309e-09 0.0014 9.312e-09 0 9.366e-09 0 9.369e-09 0.0014 9.372e-09 0 9.426e-09 0 9.429e-09 0.0014 9.432e-09 0 9.486e-09 0 9.489e-09 0.0014 9.492e-09 0 9.546e-09 0 9.549e-09 0.0014 9.552e-09 0 9.606e-09 0 9.609e-09 0.0014 9.612e-09 0 9.666e-09 0 9.669e-09 0.0014 9.672e-09 0 9.726e-09 0 9.729e-09 0.0014 9.732e-09 0 9.786e-09 0 9.789e-09 0.0014 9.792e-09 0 9.846e-09 0 9.849e-09 0.0014 9.852e-09 0 9.906e-09 0 9.909e-09 0.0014 9.912e-09 0 9.966e-09 0 9.969e-09 0.0014 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0014 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0014 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0014 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0014 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0014 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0014 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0014 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0014 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0014 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0014 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0014 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0014 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0014 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0014 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0014 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0014 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0014 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0014 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0014 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0014 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0014 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0014 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0014 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0014 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0014 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0014 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0014 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0014 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0014 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0014 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0014 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0014 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0014 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0014 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0014 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0014 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0014 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0014 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0014 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0014 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0014 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0014 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0014 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0014 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0014 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0014 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0014 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0014 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0014 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0014 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0014 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0014 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0014 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0014 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0014 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0014 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0014 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0014 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0014 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0014 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0014 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0014 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0014 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0014 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0014 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0014 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0014 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0014 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0014 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0014 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0014 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0014 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0014 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0014 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0014 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0014 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0014 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0014 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0014 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0014 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0014 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0014 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0014 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0014 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0014 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0014 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0014 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0014 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0014 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0014 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0014 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0014 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0014 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0014 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0014 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0014 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0014 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0014 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0014 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0014 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0014 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0014 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0014 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0014 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0014 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0014 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0014 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0014 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0014 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0014 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0014 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0014 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0014 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0014 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0014 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0014 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0014 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0014 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0014 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0014 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0014 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0014 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0014 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0014 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0014 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0014 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0014 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0014 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0014 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0014 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0014 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0014 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0014 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0014 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0014 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0014 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0014 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0014 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0014 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0014 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0014 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0014 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0014 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0014 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0014 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0014 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0014 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0014 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0014 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0014 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0014 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0014 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0014 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0014 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0014 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0014 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0014 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0014 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0014 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0014 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0014 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0014 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0014 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0014 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0014 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0014 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0014 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0014 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0014 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0014 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0014 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0014 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0014 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0014 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0014 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0014 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0014 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0014 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0014 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0014 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0014 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0014 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0014 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0014 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0014 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0014 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0014 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0014 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0014 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0014 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0014 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0014 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0014 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0014 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0014 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0014 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0014 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0014 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0014 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0014 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0014 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0014 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0014 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0014 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0014 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0014 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0014 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0014 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0014 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0014 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0014 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0014 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0014 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0014 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0014 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0014 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0014 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0014 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0014 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0014 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0014 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0014 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0014 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0014 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0014 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0014 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0014 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0014 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0014 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0014 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0014 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0014 2.3892e-08 0)
IT05|T 0 T05  PWL(0 0 6e-12 0 9e-12 0.0014 1.2e-11 0 6.6e-11 0 6.9e-11 0.0014 7.2e-11 0 1.26e-10 0 1.29e-10 0.0014 1.32e-10 0 1.86e-10 0 1.89e-10 0.0014 1.92e-10 0 2.46e-10 0 2.49e-10 0.0014 2.52e-10 0 3.06e-10 0 3.09e-10 0.0014 3.12e-10 0 3.66e-10 0 3.69e-10 0.0014 3.72e-10 0 4.26e-10 0 4.29e-10 0.0014 4.32e-10 0 4.86e-10 0 4.89e-10 0.0014 4.92e-10 0 5.46e-10 0 5.49e-10 0.0014 5.52e-10 0 6.06e-10 0 6.09e-10 0.0014 6.12e-10 0 6.66e-10 0 6.69e-10 0.0014 6.72e-10 0 7.26e-10 0 7.29e-10 0.0014 7.32e-10 0 7.86e-10 0 7.89e-10 0.0014 7.92e-10 0 8.46e-10 0 8.49e-10 0.0014 8.52e-10 0 9.06e-10 0 9.09e-10 0.0014 9.12e-10 0 9.66e-10 0 9.69e-10 0.0014 9.72e-10 0 1.026e-09 0 1.029e-09 0.0014 1.032e-09 0 1.086e-09 0 1.089e-09 0.0014 1.092e-09 0 1.146e-09 0 1.149e-09 0.0014 1.152e-09 0 1.206e-09 0 1.209e-09 0.0014 1.212e-09 0 1.266e-09 0 1.269e-09 0.0014 1.272e-09 0 1.326e-09 0 1.329e-09 0.0014 1.332e-09 0 1.386e-09 0 1.389e-09 0.0014 1.392e-09 0 1.446e-09 0 1.449e-09 0.0014 1.452e-09 0 1.506e-09 0 1.509e-09 0.0014 1.512e-09 0 1.566e-09 0 1.569e-09 0.0014 1.572e-09 0 1.626e-09 0 1.629e-09 0.0014 1.632e-09 0 1.686e-09 0 1.689e-09 0.0014 1.692e-09 0 1.746e-09 0 1.749e-09 0.0014 1.752e-09 0 1.806e-09 0 1.809e-09 0.0014 1.812e-09 0 1.866e-09 0 1.869e-09 0.0014 1.872e-09 0 1.926e-09 0 1.929e-09 0.0014 1.932e-09 0 1.986e-09 0 1.989e-09 0.0014 1.992e-09 0 2.046e-09 0 2.049e-09 0.0014 2.052e-09 0 2.106e-09 0 2.109e-09 0.0014 2.112e-09 0 2.166e-09 0 2.169e-09 0.0014 2.172e-09 0 2.226e-09 0 2.229e-09 0.0014 2.232e-09 0 2.286e-09 0 2.289e-09 0.0014 2.292e-09 0 2.346e-09 0 2.349e-09 0.0014 2.352e-09 0 2.406e-09 0 2.409e-09 0.0014 2.412e-09 0 2.466e-09 0 2.469e-09 0.0014 2.472e-09 0 2.526e-09 0 2.529e-09 0.0014 2.532e-09 0 2.586e-09 0 2.589e-09 0.0014 2.592e-09 0 2.646e-09 0 2.649e-09 0.0014 2.652e-09 0 2.706e-09 0 2.709e-09 0.0014 2.712e-09 0 2.766e-09 0 2.769e-09 0.0014 2.772e-09 0 2.826e-09 0 2.829e-09 0.0014 2.832e-09 0 2.886e-09 0 2.889e-09 0.0014 2.892e-09 0 2.946e-09 0 2.949e-09 0.0014 2.952e-09 0 3.006e-09 0 3.009e-09 0.0014 3.012e-09 0 3.066e-09 0 3.069e-09 0.0014 3.072e-09 0 3.126e-09 0 3.129e-09 0.0014 3.132e-09 0 3.186e-09 0 3.189e-09 0.0014 3.192e-09 0 3.246e-09 0 3.249e-09 0.0014 3.252e-09 0 3.306e-09 0 3.309e-09 0.0014 3.312e-09 0 3.366e-09 0 3.369e-09 0.0014 3.372e-09 0 3.426e-09 0 3.429e-09 0.0014 3.432e-09 0 3.486e-09 0 3.489e-09 0.0014 3.492e-09 0 3.546e-09 0 3.549e-09 0.0014 3.552e-09 0 3.606e-09 0 3.609e-09 0.0014 3.612e-09 0 3.666e-09 0 3.669e-09 0.0014 3.672e-09 0 3.726e-09 0 3.729e-09 0.0014 3.732e-09 0 3.786e-09 0 3.789e-09 0.0014 3.792e-09 0 3.846e-09 0 3.849e-09 0.0014 3.852e-09 0 3.906e-09 0 3.909e-09 0.0014 3.912e-09 0 3.966e-09 0 3.969e-09 0.0014 3.972e-09 0 4.026e-09 0 4.029e-09 0.0014 4.032e-09 0 4.086e-09 0 4.089e-09 0.0014 4.092e-09 0 4.146e-09 0 4.149e-09 0.0014 4.152e-09 0 4.206e-09 0 4.209e-09 0.0014 4.212e-09 0 4.266e-09 0 4.269e-09 0.0014 4.272e-09 0 4.326e-09 0 4.329e-09 0.0014 4.332e-09 0 4.386e-09 0 4.389e-09 0.0014 4.392e-09 0 4.446e-09 0 4.449e-09 0.0014 4.452e-09 0 4.506e-09 0 4.509e-09 0.0014 4.512e-09 0 4.566e-09 0 4.569e-09 0.0014 4.572e-09 0 4.626e-09 0 4.629e-09 0.0014 4.632e-09 0 4.686e-09 0 4.689e-09 0.0014 4.692e-09 0 4.746e-09 0 4.749e-09 0.0014 4.752e-09 0 4.806e-09 0 4.809e-09 0.0014 4.812e-09 0 4.866e-09 0 4.869e-09 0.0014 4.872e-09 0 4.926e-09 0 4.929e-09 0.0014 4.932e-09 0 4.986e-09 0 4.989e-09 0.0014 4.992e-09 0 5.046e-09 0 5.049e-09 0.0014 5.052e-09 0 5.106e-09 0 5.109e-09 0.0014 5.112e-09 0 5.166e-09 0 5.169e-09 0.0014 5.172e-09 0 5.226e-09 0 5.229e-09 0.0014 5.232e-09 0 5.286e-09 0 5.289e-09 0.0014 5.292e-09 0 5.346e-09 0 5.349e-09 0.0014 5.352e-09 0 5.406e-09 0 5.409e-09 0.0014 5.412e-09 0 5.466e-09 0 5.469e-09 0.0014 5.472e-09 0 5.526e-09 0 5.529e-09 0.0014 5.532e-09 0 5.586e-09 0 5.589e-09 0.0014 5.592e-09 0 5.646e-09 0 5.649e-09 0.0014 5.652e-09 0 5.706e-09 0 5.709e-09 0.0014 5.712e-09 0 5.766e-09 0 5.769e-09 0.0014 5.772e-09 0 5.826e-09 0 5.829e-09 0.0014 5.832e-09 0 5.886e-09 0 5.889e-09 0.0014 5.892e-09 0 5.946e-09 0 5.949e-09 0.0014 5.952e-09 0 6.006e-09 0 6.009e-09 0.0014 6.012e-09 0 6.066e-09 0 6.069e-09 0.0014 6.072e-09 0 6.126e-09 0 6.129e-09 0.0014 6.132e-09 0 6.186e-09 0 6.189e-09 0.0014 6.192e-09 0 6.246e-09 0 6.249e-09 0.0014 6.252e-09 0 6.306e-09 0 6.309e-09 0.0014 6.312e-09 0 6.366e-09 0 6.369e-09 0.0014 6.372e-09 0 6.426e-09 0 6.429e-09 0.0014 6.432e-09 0 6.486e-09 0 6.489e-09 0.0014 6.492e-09 0 6.546e-09 0 6.549e-09 0.0014 6.552e-09 0 6.606e-09 0 6.609e-09 0.0014 6.612e-09 0 6.666e-09 0 6.669e-09 0.0014 6.672e-09 0 6.726e-09 0 6.729e-09 0.0014 6.732e-09 0 6.786e-09 0 6.789e-09 0.0014 6.792e-09 0 6.846e-09 0 6.849e-09 0.0014 6.852e-09 0 6.906e-09 0 6.909e-09 0.0014 6.912e-09 0 6.966e-09 0 6.969e-09 0.0014 6.972e-09 0 7.026e-09 0 7.029e-09 0.0014 7.032e-09 0 7.086e-09 0 7.089e-09 0.0014 7.092e-09 0 7.146e-09 0 7.149e-09 0.0014 7.152e-09 0 7.206e-09 0 7.209e-09 0.0014 7.212e-09 0 7.266e-09 0 7.269e-09 0.0014 7.272e-09 0 7.326e-09 0 7.329e-09 0.0014 7.332e-09 0 7.386e-09 0 7.389e-09 0.0014 7.392e-09 0 7.446e-09 0 7.449e-09 0.0014 7.452e-09 0 7.506e-09 0 7.509e-09 0.0014 7.512e-09 0 7.566e-09 0 7.569e-09 0.0014 7.572e-09 0 7.626e-09 0 7.629e-09 0.0014 7.632e-09 0 7.686e-09 0 7.689e-09 0.0014 7.692e-09 0 7.746e-09 0 7.749e-09 0.0014 7.752e-09 0 7.806e-09 0 7.809e-09 0.0014 7.812e-09 0 7.866e-09 0 7.869e-09 0.0014 7.872e-09 0 7.926e-09 0 7.929e-09 0.0014 7.932e-09 0 7.986e-09 0 7.989e-09 0.0014 7.992e-09 0 8.046e-09 0 8.049e-09 0.0014 8.052e-09 0 8.106e-09 0 8.109e-09 0.0014 8.112e-09 0 8.166e-09 0 8.169e-09 0.0014 8.172e-09 0 8.226e-09 0 8.229e-09 0.0014 8.232e-09 0 8.286e-09 0 8.289e-09 0.0014 8.292e-09 0 8.346e-09 0 8.349e-09 0.0014 8.352e-09 0 8.406e-09 0 8.409e-09 0.0014 8.412e-09 0 8.466e-09 0 8.469e-09 0.0014 8.472e-09 0 8.526e-09 0 8.529e-09 0.0014 8.532e-09 0 8.586e-09 0 8.589e-09 0.0014 8.592e-09 0 8.646e-09 0 8.649e-09 0.0014 8.652e-09 0 8.706e-09 0 8.709e-09 0.0014 8.712e-09 0 8.766e-09 0 8.769e-09 0.0014 8.772e-09 0 8.826e-09 0 8.829e-09 0.0014 8.832e-09 0 8.886e-09 0 8.889e-09 0.0014 8.892e-09 0 8.946e-09 0 8.949e-09 0.0014 8.952e-09 0 9.006e-09 0 9.009e-09 0.0014 9.012e-09 0 9.066e-09 0 9.069e-09 0.0014 9.072e-09 0 9.126e-09 0 9.129e-09 0.0014 9.132e-09 0 9.186e-09 0 9.189e-09 0.0014 9.192e-09 0 9.246e-09 0 9.249e-09 0.0014 9.252e-09 0 9.306e-09 0 9.309e-09 0.0014 9.312e-09 0 9.366e-09 0 9.369e-09 0.0014 9.372e-09 0 9.426e-09 0 9.429e-09 0.0014 9.432e-09 0 9.486e-09 0 9.489e-09 0.0014 9.492e-09 0 9.546e-09 0 9.549e-09 0.0014 9.552e-09 0 9.606e-09 0 9.609e-09 0.0014 9.612e-09 0 9.666e-09 0 9.669e-09 0.0014 9.672e-09 0 9.726e-09 0 9.729e-09 0.0014 9.732e-09 0 9.786e-09 0 9.789e-09 0.0014 9.792e-09 0 9.846e-09 0 9.849e-09 0.0014 9.852e-09 0 9.906e-09 0 9.909e-09 0.0014 9.912e-09 0 9.966e-09 0 9.969e-09 0.0014 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0014 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0014 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0014 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0014 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0014 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0014 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0014 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0014 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0014 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0014 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0014 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0014 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0014 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0014 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0014 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0014 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0014 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0014 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0014 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0014 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0014 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0014 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0014 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0014 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0014 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0014 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0014 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0014 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0014 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0014 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0014 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0014 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0014 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0014 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0014 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0014 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0014 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0014 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0014 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0014 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0014 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0014 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0014 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0014 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0014 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0014 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0014 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0014 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0014 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0014 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0014 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0014 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0014 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0014 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0014 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0014 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0014 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0014 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0014 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0014 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0014 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0014 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0014 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0014 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0014 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0014 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0014 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0014 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0014 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0014 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0014 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0014 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0014 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0014 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0014 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0014 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0014 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0014 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0014 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0014 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0014 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0014 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0014 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0014 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0014 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0014 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0014 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0014 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0014 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0014 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0014 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0014 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0014 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0014 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0014 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0014 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0014 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0014 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0014 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0014 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0014 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0014 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0014 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0014 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0014 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0014 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0014 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0014 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0014 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0014 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0014 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0014 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0014 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0014 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0014 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0014 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0014 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0014 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0014 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0014 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0014 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0014 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0014 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0014 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0014 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0014 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0014 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0014 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0014 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0014 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0014 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0014 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0014 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0014 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0014 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0014 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0014 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0014 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0014 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0014 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0014 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0014 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0014 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0014 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0014 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0014 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0014 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0014 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0014 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0014 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0014 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0014 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0014 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0014 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0014 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0014 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0014 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0014 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0014 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0014 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0014 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0014 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0014 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0014 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0014 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0014 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0014 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0014 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0014 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0014 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0014 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0014 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0014 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0014 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0014 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0014 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0014 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0014 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0014 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0014 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0014 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0014 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0014 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0014 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0014 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0014 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0014 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0014 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0014 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0014 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0014 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0014 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0014 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0014 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0014 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0014 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0014 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0014 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0014 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0014 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0014 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0014 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0014 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0014 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0014 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0014 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0014 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0014 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0014 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0014 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0014 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0014 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0014 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0014 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0014 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0014 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0014 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0014 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0014 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0014 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0014 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0014 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0014 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0014 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0014 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0014 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0014 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0014 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0014 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0014 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0014 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0014 2.3892e-08 0)
IT06|T 0 T06  PWL(0 0 6e-12 0 9e-12 0.0014 1.2e-11 0 6.6e-11 0 6.9e-11 0.0014 7.2e-11 0 1.26e-10 0 1.29e-10 0.0014 1.32e-10 0 1.86e-10 0 1.89e-10 0.0014 1.92e-10 0 2.46e-10 0 2.49e-10 0.0014 2.52e-10 0 3.06e-10 0 3.09e-10 0.0014 3.12e-10 0 3.66e-10 0 3.69e-10 0.0014 3.72e-10 0 4.26e-10 0 4.29e-10 0.0014 4.32e-10 0 4.86e-10 0 4.89e-10 0.0014 4.92e-10 0 5.46e-10 0 5.49e-10 0.0014 5.52e-10 0 6.06e-10 0 6.09e-10 0.0014 6.12e-10 0 6.66e-10 0 6.69e-10 0.0014 6.72e-10 0 7.26e-10 0 7.29e-10 0.0014 7.32e-10 0 7.86e-10 0 7.89e-10 0.0014 7.92e-10 0 8.46e-10 0 8.49e-10 0.0014 8.52e-10 0 9.06e-10 0 9.09e-10 0.0014 9.12e-10 0 9.66e-10 0 9.69e-10 0.0014 9.72e-10 0 1.026e-09 0 1.029e-09 0.0014 1.032e-09 0 1.086e-09 0 1.089e-09 0.0014 1.092e-09 0 1.146e-09 0 1.149e-09 0.0014 1.152e-09 0 1.206e-09 0 1.209e-09 0.0014 1.212e-09 0 1.266e-09 0 1.269e-09 0.0014 1.272e-09 0 1.326e-09 0 1.329e-09 0.0014 1.332e-09 0 1.386e-09 0 1.389e-09 0.0014 1.392e-09 0 1.446e-09 0 1.449e-09 0.0014 1.452e-09 0 1.506e-09 0 1.509e-09 0.0014 1.512e-09 0 1.566e-09 0 1.569e-09 0.0014 1.572e-09 0 1.626e-09 0 1.629e-09 0.0014 1.632e-09 0 1.686e-09 0 1.689e-09 0.0014 1.692e-09 0 1.746e-09 0 1.749e-09 0.0014 1.752e-09 0 1.806e-09 0 1.809e-09 0.0014 1.812e-09 0 1.866e-09 0 1.869e-09 0.0014 1.872e-09 0 1.926e-09 0 1.929e-09 0.0014 1.932e-09 0 1.986e-09 0 1.989e-09 0.0014 1.992e-09 0 2.046e-09 0 2.049e-09 0.0014 2.052e-09 0 2.106e-09 0 2.109e-09 0.0014 2.112e-09 0 2.166e-09 0 2.169e-09 0.0014 2.172e-09 0 2.226e-09 0 2.229e-09 0.0014 2.232e-09 0 2.286e-09 0 2.289e-09 0.0014 2.292e-09 0 2.346e-09 0 2.349e-09 0.0014 2.352e-09 0 2.406e-09 0 2.409e-09 0.0014 2.412e-09 0 2.466e-09 0 2.469e-09 0.0014 2.472e-09 0 2.526e-09 0 2.529e-09 0.0014 2.532e-09 0 2.586e-09 0 2.589e-09 0.0014 2.592e-09 0 2.646e-09 0 2.649e-09 0.0014 2.652e-09 0 2.706e-09 0 2.709e-09 0.0014 2.712e-09 0 2.766e-09 0 2.769e-09 0.0014 2.772e-09 0 2.826e-09 0 2.829e-09 0.0014 2.832e-09 0 2.886e-09 0 2.889e-09 0.0014 2.892e-09 0 2.946e-09 0 2.949e-09 0.0014 2.952e-09 0 3.006e-09 0 3.009e-09 0.0014 3.012e-09 0 3.066e-09 0 3.069e-09 0.0014 3.072e-09 0 3.126e-09 0 3.129e-09 0.0014 3.132e-09 0 3.186e-09 0 3.189e-09 0.0014 3.192e-09 0 3.246e-09 0 3.249e-09 0.0014 3.252e-09 0 3.306e-09 0 3.309e-09 0.0014 3.312e-09 0 3.366e-09 0 3.369e-09 0.0014 3.372e-09 0 3.426e-09 0 3.429e-09 0.0014 3.432e-09 0 3.486e-09 0 3.489e-09 0.0014 3.492e-09 0 3.546e-09 0 3.549e-09 0.0014 3.552e-09 0 3.606e-09 0 3.609e-09 0.0014 3.612e-09 0 3.666e-09 0 3.669e-09 0.0014 3.672e-09 0 3.726e-09 0 3.729e-09 0.0014 3.732e-09 0 3.786e-09 0 3.789e-09 0.0014 3.792e-09 0 3.846e-09 0 3.849e-09 0.0014 3.852e-09 0 3.906e-09 0 3.909e-09 0.0014 3.912e-09 0 3.966e-09 0 3.969e-09 0.0014 3.972e-09 0 4.026e-09 0 4.029e-09 0.0014 4.032e-09 0 4.086e-09 0 4.089e-09 0.0014 4.092e-09 0 4.146e-09 0 4.149e-09 0.0014 4.152e-09 0 4.206e-09 0 4.209e-09 0.0014 4.212e-09 0 4.266e-09 0 4.269e-09 0.0014 4.272e-09 0 4.326e-09 0 4.329e-09 0.0014 4.332e-09 0 4.386e-09 0 4.389e-09 0.0014 4.392e-09 0 4.446e-09 0 4.449e-09 0.0014 4.452e-09 0 4.506e-09 0 4.509e-09 0.0014 4.512e-09 0 4.566e-09 0 4.569e-09 0.0014 4.572e-09 0 4.626e-09 0 4.629e-09 0.0014 4.632e-09 0 4.686e-09 0 4.689e-09 0.0014 4.692e-09 0 4.746e-09 0 4.749e-09 0.0014 4.752e-09 0 4.806e-09 0 4.809e-09 0.0014 4.812e-09 0 4.866e-09 0 4.869e-09 0.0014 4.872e-09 0 4.926e-09 0 4.929e-09 0.0014 4.932e-09 0 4.986e-09 0 4.989e-09 0.0014 4.992e-09 0 5.046e-09 0 5.049e-09 0.0014 5.052e-09 0 5.106e-09 0 5.109e-09 0.0014 5.112e-09 0 5.166e-09 0 5.169e-09 0.0014 5.172e-09 0 5.226e-09 0 5.229e-09 0.0014 5.232e-09 0 5.286e-09 0 5.289e-09 0.0014 5.292e-09 0 5.346e-09 0 5.349e-09 0.0014 5.352e-09 0 5.406e-09 0 5.409e-09 0.0014 5.412e-09 0 5.466e-09 0 5.469e-09 0.0014 5.472e-09 0 5.526e-09 0 5.529e-09 0.0014 5.532e-09 0 5.586e-09 0 5.589e-09 0.0014 5.592e-09 0 5.646e-09 0 5.649e-09 0.0014 5.652e-09 0 5.706e-09 0 5.709e-09 0.0014 5.712e-09 0 5.766e-09 0 5.769e-09 0.0014 5.772e-09 0 5.826e-09 0 5.829e-09 0.0014 5.832e-09 0 5.886e-09 0 5.889e-09 0.0014 5.892e-09 0 5.946e-09 0 5.949e-09 0.0014 5.952e-09 0 6.006e-09 0 6.009e-09 0.0014 6.012e-09 0 6.066e-09 0 6.069e-09 0.0014 6.072e-09 0 6.126e-09 0 6.129e-09 0.0014 6.132e-09 0 6.186e-09 0 6.189e-09 0.0014 6.192e-09 0 6.246e-09 0 6.249e-09 0.0014 6.252e-09 0 6.306e-09 0 6.309e-09 0.0014 6.312e-09 0 6.366e-09 0 6.369e-09 0.0014 6.372e-09 0 6.426e-09 0 6.429e-09 0.0014 6.432e-09 0 6.486e-09 0 6.489e-09 0.0014 6.492e-09 0 6.546e-09 0 6.549e-09 0.0014 6.552e-09 0 6.606e-09 0 6.609e-09 0.0014 6.612e-09 0 6.666e-09 0 6.669e-09 0.0014 6.672e-09 0 6.726e-09 0 6.729e-09 0.0014 6.732e-09 0 6.786e-09 0 6.789e-09 0.0014 6.792e-09 0 6.846e-09 0 6.849e-09 0.0014 6.852e-09 0 6.906e-09 0 6.909e-09 0.0014 6.912e-09 0 6.966e-09 0 6.969e-09 0.0014 6.972e-09 0 7.026e-09 0 7.029e-09 0.0014 7.032e-09 0 7.086e-09 0 7.089e-09 0.0014 7.092e-09 0 7.146e-09 0 7.149e-09 0.0014 7.152e-09 0 7.206e-09 0 7.209e-09 0.0014 7.212e-09 0 7.266e-09 0 7.269e-09 0.0014 7.272e-09 0 7.326e-09 0 7.329e-09 0.0014 7.332e-09 0 7.386e-09 0 7.389e-09 0.0014 7.392e-09 0 7.446e-09 0 7.449e-09 0.0014 7.452e-09 0 7.506e-09 0 7.509e-09 0.0014 7.512e-09 0 7.566e-09 0 7.569e-09 0.0014 7.572e-09 0 7.626e-09 0 7.629e-09 0.0014 7.632e-09 0 7.686e-09 0 7.689e-09 0.0014 7.692e-09 0 7.746e-09 0 7.749e-09 0.0014 7.752e-09 0 7.806e-09 0 7.809e-09 0.0014 7.812e-09 0 7.866e-09 0 7.869e-09 0.0014 7.872e-09 0 7.926e-09 0 7.929e-09 0.0014 7.932e-09 0 7.986e-09 0 7.989e-09 0.0014 7.992e-09 0 8.046e-09 0 8.049e-09 0.0014 8.052e-09 0 8.106e-09 0 8.109e-09 0.0014 8.112e-09 0 8.166e-09 0 8.169e-09 0.0014 8.172e-09 0 8.226e-09 0 8.229e-09 0.0014 8.232e-09 0 8.286e-09 0 8.289e-09 0.0014 8.292e-09 0 8.346e-09 0 8.349e-09 0.0014 8.352e-09 0 8.406e-09 0 8.409e-09 0.0014 8.412e-09 0 8.466e-09 0 8.469e-09 0.0014 8.472e-09 0 8.526e-09 0 8.529e-09 0.0014 8.532e-09 0 8.586e-09 0 8.589e-09 0.0014 8.592e-09 0 8.646e-09 0 8.649e-09 0.0014 8.652e-09 0 8.706e-09 0 8.709e-09 0.0014 8.712e-09 0 8.766e-09 0 8.769e-09 0.0014 8.772e-09 0 8.826e-09 0 8.829e-09 0.0014 8.832e-09 0 8.886e-09 0 8.889e-09 0.0014 8.892e-09 0 8.946e-09 0 8.949e-09 0.0014 8.952e-09 0 9.006e-09 0 9.009e-09 0.0014 9.012e-09 0 9.066e-09 0 9.069e-09 0.0014 9.072e-09 0 9.126e-09 0 9.129e-09 0.0014 9.132e-09 0 9.186e-09 0 9.189e-09 0.0014 9.192e-09 0 9.246e-09 0 9.249e-09 0.0014 9.252e-09 0 9.306e-09 0 9.309e-09 0.0014 9.312e-09 0 9.366e-09 0 9.369e-09 0.0014 9.372e-09 0 9.426e-09 0 9.429e-09 0.0014 9.432e-09 0 9.486e-09 0 9.489e-09 0.0014 9.492e-09 0 9.546e-09 0 9.549e-09 0.0014 9.552e-09 0 9.606e-09 0 9.609e-09 0.0014 9.612e-09 0 9.666e-09 0 9.669e-09 0.0014 9.672e-09 0 9.726e-09 0 9.729e-09 0.0014 9.732e-09 0 9.786e-09 0 9.789e-09 0.0014 9.792e-09 0 9.846e-09 0 9.849e-09 0.0014 9.852e-09 0 9.906e-09 0 9.909e-09 0.0014 9.912e-09 0 9.966e-09 0 9.969e-09 0.0014 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0014 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0014 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0014 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0014 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0014 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0014 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0014 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0014 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0014 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0014 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0014 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0014 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0014 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0014 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0014 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0014 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0014 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0014 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0014 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0014 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0014 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0014 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0014 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0014 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0014 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0014 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0014 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0014 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0014 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0014 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0014 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0014 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0014 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0014 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0014 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0014 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0014 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0014 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0014 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0014 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0014 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0014 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0014 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0014 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0014 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0014 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0014 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0014 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0014 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0014 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0014 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0014 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0014 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0014 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0014 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0014 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0014 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0014 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0014 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0014 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0014 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0014 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0014 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0014 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0014 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0014 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0014 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0014 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0014 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0014 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0014 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0014 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0014 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0014 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0014 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0014 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0014 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0014 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0014 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0014 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0014 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0014 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0014 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0014 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0014 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0014 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0014 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0014 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0014 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0014 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0014 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0014 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0014 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0014 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0014 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0014 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0014 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0014 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0014 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0014 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0014 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0014 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0014 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0014 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0014 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0014 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0014 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0014 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0014 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0014 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0014 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0014 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0014 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0014 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0014 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0014 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0014 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0014 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0014 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0014 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0014 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0014 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0014 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0014 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0014 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0014 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0014 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0014 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0014 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0014 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0014 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0014 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0014 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0014 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0014 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0014 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0014 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0014 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0014 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0014 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0014 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0014 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0014 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0014 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0014 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0014 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0014 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0014 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0014 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0014 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0014 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0014 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0014 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0014 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0014 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0014 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0014 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0014 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0014 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0014 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0014 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0014 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0014 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0014 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0014 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0014 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0014 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0014 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0014 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0014 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0014 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0014 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0014 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0014 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0014 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0014 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0014 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0014 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0014 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0014 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0014 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0014 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0014 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0014 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0014 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0014 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0014 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0014 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0014 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0014 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0014 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0014 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0014 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0014 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0014 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0014 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0014 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0014 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0014 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0014 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0014 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0014 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0014 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0014 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0014 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0014 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0014 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0014 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0014 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0014 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0014 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0014 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0014 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0014 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0014 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0014 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0014 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0014 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0014 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0014 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0014 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0014 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0014 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0014 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0014 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0014 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0014 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0014 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0014 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0014 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0014 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0014 2.3892e-08 0)
IT07|T 0 T07  PWL(0 0 6e-12 0 9e-12 0.0028 1.2e-11 0 6.6e-11 0 6.9e-11 0.0028 7.2e-11 0 1.26e-10 0 1.29e-10 0.0028 1.32e-10 0 1.86e-10 0 1.89e-10 0.0028 1.92e-10 0 2.46e-10 0 2.49e-10 0.0028 2.52e-10 0 3.06e-10 0 3.09e-10 0.0028 3.12e-10 0 3.66e-10 0 3.69e-10 0.0028 3.72e-10 0 4.26e-10 0 4.29e-10 0.0028 4.32e-10 0 4.86e-10 0 4.89e-10 0.0028 4.92e-10 0 5.46e-10 0 5.49e-10 0.0028 5.52e-10 0 6.06e-10 0 6.09e-10 0.0028 6.12e-10 0 6.66e-10 0 6.69e-10 0.0028 6.72e-10 0 7.26e-10 0 7.29e-10 0.0028 7.32e-10 0 7.86e-10 0 7.89e-10 0.0028 7.92e-10 0 8.46e-10 0 8.49e-10 0.0028 8.52e-10 0 9.06e-10 0 9.09e-10 0.0028 9.12e-10 0 9.66e-10 0 9.69e-10 0.0028 9.72e-10 0 1.026e-09 0 1.029e-09 0.0028 1.032e-09 0 1.086e-09 0 1.089e-09 0.0028 1.092e-09 0 1.146e-09 0 1.149e-09 0.0028 1.152e-09 0 1.206e-09 0 1.209e-09 0.0028 1.212e-09 0 1.266e-09 0 1.269e-09 0.0028 1.272e-09 0 1.326e-09 0 1.329e-09 0.0028 1.332e-09 0 1.386e-09 0 1.389e-09 0.0028 1.392e-09 0 1.446e-09 0 1.449e-09 0.0028 1.452e-09 0 1.506e-09 0 1.509e-09 0.0028 1.512e-09 0 1.566e-09 0 1.569e-09 0.0028 1.572e-09 0 1.626e-09 0 1.629e-09 0.0028 1.632e-09 0 1.686e-09 0 1.689e-09 0.0028 1.692e-09 0 1.746e-09 0 1.749e-09 0.0028 1.752e-09 0 1.806e-09 0 1.809e-09 0.0028 1.812e-09 0 1.866e-09 0 1.869e-09 0.0028 1.872e-09 0 1.926e-09 0 1.929e-09 0.0028 1.932e-09 0 1.986e-09 0 1.989e-09 0.0028 1.992e-09 0 2.046e-09 0 2.049e-09 0.0028 2.052e-09 0 2.106e-09 0 2.109e-09 0.0028 2.112e-09 0 2.166e-09 0 2.169e-09 0.0028 2.172e-09 0 2.226e-09 0 2.229e-09 0.0028 2.232e-09 0 2.286e-09 0 2.289e-09 0.0028 2.292e-09 0 2.346e-09 0 2.349e-09 0.0028 2.352e-09 0 2.406e-09 0 2.409e-09 0.0028 2.412e-09 0 2.466e-09 0 2.469e-09 0.0028 2.472e-09 0 2.526e-09 0 2.529e-09 0.0028 2.532e-09 0 2.586e-09 0 2.589e-09 0.0028 2.592e-09 0 2.646e-09 0 2.649e-09 0.0028 2.652e-09 0 2.706e-09 0 2.709e-09 0.0028 2.712e-09 0 2.766e-09 0 2.769e-09 0.0028 2.772e-09 0 2.826e-09 0 2.829e-09 0.0028 2.832e-09 0 2.886e-09 0 2.889e-09 0.0028 2.892e-09 0 2.946e-09 0 2.949e-09 0.0028 2.952e-09 0 3.006e-09 0 3.009e-09 0.0028 3.012e-09 0 3.066e-09 0 3.069e-09 0.0028 3.072e-09 0 3.126e-09 0 3.129e-09 0.0028 3.132e-09 0 3.186e-09 0 3.189e-09 0.0028 3.192e-09 0 3.246e-09 0 3.249e-09 0.0028 3.252e-09 0 3.306e-09 0 3.309e-09 0.0028 3.312e-09 0 3.366e-09 0 3.369e-09 0.0028 3.372e-09 0 3.426e-09 0 3.429e-09 0.0028 3.432e-09 0 3.486e-09 0 3.489e-09 0.0028 3.492e-09 0 3.546e-09 0 3.549e-09 0.0028 3.552e-09 0 3.606e-09 0 3.609e-09 0.0028 3.612e-09 0 3.666e-09 0 3.669e-09 0.0028 3.672e-09 0 3.726e-09 0 3.729e-09 0.0028 3.732e-09 0 3.786e-09 0 3.789e-09 0.0028 3.792e-09 0 3.846e-09 0 3.849e-09 0.0028 3.852e-09 0 3.906e-09 0 3.909e-09 0.0028 3.912e-09 0 3.966e-09 0 3.969e-09 0.0028 3.972e-09 0 4.026e-09 0 4.029e-09 0.0028 4.032e-09 0 4.086e-09 0 4.089e-09 0.0028 4.092e-09 0 4.146e-09 0 4.149e-09 0.0028 4.152e-09 0 4.206e-09 0 4.209e-09 0.0028 4.212e-09 0 4.266e-09 0 4.269e-09 0.0028 4.272e-09 0 4.326e-09 0 4.329e-09 0.0028 4.332e-09 0 4.386e-09 0 4.389e-09 0.0028 4.392e-09 0 4.446e-09 0 4.449e-09 0.0028 4.452e-09 0 4.506e-09 0 4.509e-09 0.0028 4.512e-09 0 4.566e-09 0 4.569e-09 0.0028 4.572e-09 0 4.626e-09 0 4.629e-09 0.0028 4.632e-09 0 4.686e-09 0 4.689e-09 0.0028 4.692e-09 0 4.746e-09 0 4.749e-09 0.0028 4.752e-09 0 4.806e-09 0 4.809e-09 0.0028 4.812e-09 0 4.866e-09 0 4.869e-09 0.0028 4.872e-09 0 4.926e-09 0 4.929e-09 0.0028 4.932e-09 0 4.986e-09 0 4.989e-09 0.0028 4.992e-09 0 5.046e-09 0 5.049e-09 0.0028 5.052e-09 0 5.106e-09 0 5.109e-09 0.0028 5.112e-09 0 5.166e-09 0 5.169e-09 0.0028 5.172e-09 0 5.226e-09 0 5.229e-09 0.0028 5.232e-09 0 5.286e-09 0 5.289e-09 0.0028 5.292e-09 0 5.346e-09 0 5.349e-09 0.0028 5.352e-09 0 5.406e-09 0 5.409e-09 0.0028 5.412e-09 0 5.466e-09 0 5.469e-09 0.0028 5.472e-09 0 5.526e-09 0 5.529e-09 0.0028 5.532e-09 0 5.586e-09 0 5.589e-09 0.0028 5.592e-09 0 5.646e-09 0 5.649e-09 0.0028 5.652e-09 0 5.706e-09 0 5.709e-09 0.0028 5.712e-09 0 5.766e-09 0 5.769e-09 0.0028 5.772e-09 0 5.826e-09 0 5.829e-09 0.0028 5.832e-09 0 5.886e-09 0 5.889e-09 0.0028 5.892e-09 0 5.946e-09 0 5.949e-09 0.0028 5.952e-09 0 6.006e-09 0 6.009e-09 0.0028 6.012e-09 0 6.066e-09 0 6.069e-09 0.0028 6.072e-09 0 6.126e-09 0 6.129e-09 0.0028 6.132e-09 0 6.186e-09 0 6.189e-09 0.0028 6.192e-09 0 6.246e-09 0 6.249e-09 0.0028 6.252e-09 0 6.306e-09 0 6.309e-09 0.0028 6.312e-09 0 6.366e-09 0 6.369e-09 0.0028 6.372e-09 0 6.426e-09 0 6.429e-09 0.0028 6.432e-09 0 6.486e-09 0 6.489e-09 0.0028 6.492e-09 0 6.546e-09 0 6.549e-09 0.0028 6.552e-09 0 6.606e-09 0 6.609e-09 0.0028 6.612e-09 0 6.666e-09 0 6.669e-09 0.0028 6.672e-09 0 6.726e-09 0 6.729e-09 0.0028 6.732e-09 0 6.786e-09 0 6.789e-09 0.0028 6.792e-09 0 6.846e-09 0 6.849e-09 0.0028 6.852e-09 0 6.906e-09 0 6.909e-09 0.0028 6.912e-09 0 6.966e-09 0 6.969e-09 0.0028 6.972e-09 0 7.026e-09 0 7.029e-09 0.0028 7.032e-09 0 7.086e-09 0 7.089e-09 0.0028 7.092e-09 0 7.146e-09 0 7.149e-09 0.0028 7.152e-09 0 7.206e-09 0 7.209e-09 0.0028 7.212e-09 0 7.266e-09 0 7.269e-09 0.0028 7.272e-09 0 7.326e-09 0 7.329e-09 0.0028 7.332e-09 0 7.386e-09 0 7.389e-09 0.0028 7.392e-09 0 7.446e-09 0 7.449e-09 0.0028 7.452e-09 0 7.506e-09 0 7.509e-09 0.0028 7.512e-09 0 7.566e-09 0 7.569e-09 0.0028 7.572e-09 0 7.626e-09 0 7.629e-09 0.0028 7.632e-09 0 7.686e-09 0 7.689e-09 0.0028 7.692e-09 0 7.746e-09 0 7.749e-09 0.0028 7.752e-09 0 7.806e-09 0 7.809e-09 0.0028 7.812e-09 0 7.866e-09 0 7.869e-09 0.0028 7.872e-09 0 7.926e-09 0 7.929e-09 0.0028 7.932e-09 0 7.986e-09 0 7.989e-09 0.0028 7.992e-09 0 8.046e-09 0 8.049e-09 0.0028 8.052e-09 0 8.106e-09 0 8.109e-09 0.0028 8.112e-09 0 8.166e-09 0 8.169e-09 0.0028 8.172e-09 0 8.226e-09 0 8.229e-09 0.0028 8.232e-09 0 8.286e-09 0 8.289e-09 0.0028 8.292e-09 0 8.346e-09 0 8.349e-09 0.0028 8.352e-09 0 8.406e-09 0 8.409e-09 0.0028 8.412e-09 0 8.466e-09 0 8.469e-09 0.0028 8.472e-09 0 8.526e-09 0 8.529e-09 0.0028 8.532e-09 0 8.586e-09 0 8.589e-09 0.0028 8.592e-09 0 8.646e-09 0 8.649e-09 0.0028 8.652e-09 0 8.706e-09 0 8.709e-09 0.0028 8.712e-09 0 8.766e-09 0 8.769e-09 0.0028 8.772e-09 0 8.826e-09 0 8.829e-09 0.0028 8.832e-09 0 8.886e-09 0 8.889e-09 0.0028 8.892e-09 0 8.946e-09 0 8.949e-09 0.0028 8.952e-09 0 9.006e-09 0 9.009e-09 0.0028 9.012e-09 0 9.066e-09 0 9.069e-09 0.0028 9.072e-09 0 9.126e-09 0 9.129e-09 0.0028 9.132e-09 0 9.186e-09 0 9.189e-09 0.0028 9.192e-09 0 9.246e-09 0 9.249e-09 0.0028 9.252e-09 0 9.306e-09 0 9.309e-09 0.0028 9.312e-09 0 9.366e-09 0 9.369e-09 0.0028 9.372e-09 0 9.426e-09 0 9.429e-09 0.0028 9.432e-09 0 9.486e-09 0 9.489e-09 0.0028 9.492e-09 0 9.546e-09 0 9.549e-09 0.0028 9.552e-09 0 9.606e-09 0 9.609e-09 0.0028 9.612e-09 0 9.666e-09 0 9.669e-09 0.0028 9.672e-09 0 9.726e-09 0 9.729e-09 0.0028 9.732e-09 0 9.786e-09 0 9.789e-09 0.0028 9.792e-09 0 9.846e-09 0 9.849e-09 0.0028 9.852e-09 0 9.906e-09 0 9.909e-09 0.0028 9.912e-09 0 9.966e-09 0 9.969e-09 0.0028 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0028 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0028 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0028 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0028 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0028 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0028 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0028 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0028 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0028 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0028 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0028 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0028 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0028 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0028 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0028 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0028 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0028 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0028 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0028 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0028 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0028 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0028 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0028 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0028 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0028 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0028 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0028 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0028 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0028 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0028 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0028 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0028 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0028 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0028 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0028 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0028 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0028 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0028 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0028 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0028 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0028 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0028 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0028 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0028 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0028 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0028 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0028 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0028 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0028 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0028 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0028 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0028 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0028 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0028 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0028 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0028 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0028 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0028 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0028 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0028 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0028 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0028 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0028 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0028 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0028 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0028 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0028 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0028 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0028 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0028 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0028 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0028 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0028 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0028 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0028 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0028 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0028 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0028 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0028 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0028 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0028 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0028 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0028 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0028 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0028 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0028 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0028 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0028 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0028 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0028 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0028 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0028 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0028 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0028 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0028 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0028 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0028 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0028 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0028 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0028 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0028 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0028 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0028 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0028 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0028 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0028 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0028 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0028 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0028 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0028 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0028 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0028 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0028 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0028 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0028 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0028 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0028 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0028 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0028 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0028 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0028 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0028 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0028 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0028 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0028 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0028 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0028 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0028 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0028 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0028 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0028 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0028 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0028 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0028 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0028 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0028 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0028 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0028 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0028 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0028 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0028 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0028 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0028 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0028 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0028 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0028 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0028 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0028 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0028 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0028 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0028 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0028 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0028 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0028 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0028 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0028 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0028 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0028 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0028 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0028 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0028 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0028 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0028 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0028 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0028 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0028 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0028 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0028 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0028 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0028 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0028 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0028 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0028 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0028 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0028 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0028 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0028 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0028 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0028 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0028 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0028 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0028 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0028 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0028 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0028 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0028 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0028 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0028 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0028 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0028 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0028 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0028 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0028 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0028 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0028 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0028 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0028 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0028 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0028 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0028 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0028 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0028 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0028 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0028 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0028 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0028 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0028 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0028 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0028 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0028 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0028 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0028 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0028 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0028 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0028 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0028 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0028 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0028 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0028 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0028 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0028 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0028 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0028 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0028 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0028 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0028 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0028 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0028 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0028 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0028 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0028 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0028 2.3892e-08 0)
ID01|T 0 D01  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 6.6e-11 0 6.9e-11 0.0007 7.2e-11 0 1.26e-10 0 1.29e-10 0.0007 1.32e-10 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 2.46e-10 0 2.49e-10 0.0007 2.52e-10 0 3.06e-10 0 3.09e-10 0.0007 3.12e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 4.26e-10 0 4.29e-10 0.0007 4.32e-10 0 4.86e-10 0 4.89e-10 0.0007 4.92e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 6.06e-10 0 6.09e-10 0.0007 6.12e-10 0 6.66e-10 0 6.69e-10 0.0007 6.72e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 7.86e-10 0 7.89e-10 0.0007 7.92e-10 0 8.46e-10 0 8.49e-10 0.0007 8.52e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 9.66e-10 0 9.69e-10 0.0007 9.72e-10 0 1.026e-09 0 1.029e-09 0.0007 1.032e-09 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.146e-09 0 1.149e-09 0.0007 1.152e-09 0 1.206e-09 0 1.209e-09 0.0007 1.212e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.326e-09 0 1.329e-09 0.0007 1.332e-09 0 1.386e-09 0 1.389e-09 0.0007 1.392e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.506e-09 0 1.509e-09 0.0007 1.512e-09 0 1.566e-09 0 1.569e-09 0.0007 1.572e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.686e-09 0 1.689e-09 0.0007 1.692e-09 0 1.746e-09 0 1.749e-09 0.0007 1.752e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.866e-09 0 1.869e-09 0.0007 1.872e-09 0 1.926e-09 0 1.929e-09 0.0007 1.932e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.046e-09 0 2.049e-09 0.0007 2.052e-09 0 2.106e-09 0 2.109e-09 0.0007 2.112e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.226e-09 0 2.229e-09 0.0007 2.232e-09 0 2.286e-09 0 2.289e-09 0.0007 2.292e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.406e-09 0 2.409e-09 0.0007 2.412e-09 0 2.466e-09 0 2.469e-09 0.0007 2.472e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.586e-09 0 2.589e-09 0.0007 2.592e-09 0 2.646e-09 0 2.649e-09 0.0007 2.652e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.766e-09 0 2.769e-09 0.0007 2.772e-09 0 2.826e-09 0 2.829e-09 0.0007 2.832e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 2.946e-09 0 2.949e-09 0.0007 2.952e-09 0 3.006e-09 0 3.009e-09 0.0007 3.012e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.126e-09 0 3.129e-09 0.0007 3.132e-09 0 3.186e-09 0 3.189e-09 0.0007 3.192e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.306e-09 0 3.309e-09 0.0007 3.312e-09 0 3.366e-09 0 3.369e-09 0.0007 3.372e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.486e-09 0 3.489e-09 0.0007 3.492e-09 0 3.546e-09 0 3.549e-09 0.0007 3.552e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.666e-09 0 3.669e-09 0.0007 3.672e-09 0 3.726e-09 0 3.729e-09 0.0007 3.732e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.846e-09 0 3.849e-09 0.0007 3.852e-09 0 3.906e-09 0 3.909e-09 0.0007 3.912e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.026e-09 0 4.029e-09 0.0007 4.032e-09 0 4.086e-09 0 4.089e-09 0.0007 4.092e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.206e-09 0 4.209e-09 0.0007 4.212e-09 0 4.266e-09 0 4.269e-09 0.0007 4.272e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.386e-09 0 4.389e-09 0.0007 4.392e-09 0 4.446e-09 0 4.449e-09 0.0007 4.452e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.566e-09 0 4.569e-09 0.0007 4.572e-09 0 4.626e-09 0 4.629e-09 0.0007 4.632e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.746e-09 0 4.749e-09 0.0007 4.752e-09 0 4.806e-09 0 4.809e-09 0.0007 4.812e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 4.926e-09 0 4.929e-09 0.0007 4.932e-09 0 4.986e-09 0 4.989e-09 0.0007 4.992e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.106e-09 0 5.109e-09 0.0007 5.112e-09 0 5.166e-09 0 5.169e-09 0.0007 5.172e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.286e-09 0 5.289e-09 0.0007 5.292e-09 0 5.346e-09 0 5.349e-09 0.0007 5.352e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.466e-09 0 5.469e-09 0.0007 5.472e-09 0 5.526e-09 0 5.529e-09 0.0007 5.532e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.646e-09 0 5.649e-09 0.0007 5.652e-09 0 5.706e-09 0 5.709e-09 0.0007 5.712e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.826e-09 0 5.829e-09 0.0007 5.832e-09 0 5.886e-09 0 5.889e-09 0.0007 5.892e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.006e-09 0 6.009e-09 0.0007 6.012e-09 0 6.066e-09 0 6.069e-09 0.0007 6.072e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.186e-09 0 6.189e-09 0.0007 6.192e-09 0 6.246e-09 0 6.249e-09 0.0007 6.252e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.366e-09 0 6.369e-09 0.0007 6.372e-09 0 6.426e-09 0 6.429e-09 0.0007 6.432e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.546e-09 0 6.549e-09 0.0007 6.552e-09 0 6.606e-09 0 6.609e-09 0.0007 6.612e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.726e-09 0 6.729e-09 0.0007 6.732e-09 0 6.786e-09 0 6.789e-09 0.0007 6.792e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 6.906e-09 0 6.909e-09 0.0007 6.912e-09 0 6.966e-09 0 6.969e-09 0.0007 6.972e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.086e-09 0 7.089e-09 0.0007 7.092e-09 0 7.146e-09 0 7.149e-09 0.0007 7.152e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.266e-09 0 7.269e-09 0.0007 7.272e-09 0 7.326e-09 0 7.329e-09 0.0007 7.332e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.446e-09 0 7.449e-09 0.0007 7.452e-09 0 7.506e-09 0 7.509e-09 0.0007 7.512e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.626e-09 0 7.629e-09 0.0007 7.632e-09 0 7.686e-09 0 7.689e-09 0.0007 7.692e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.806e-09 0 7.809e-09 0.0007 7.812e-09 0 7.866e-09 0 7.869e-09 0.0007 7.872e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 7.986e-09 0 7.989e-09 0.0007 7.992e-09 0 8.046e-09 0 8.049e-09 0.0007 8.052e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.166e-09 0 8.169e-09 0.0007 8.172e-09 0 8.226e-09 0 8.229e-09 0.0007 8.232e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.346e-09 0 8.349e-09 0.0007 8.352e-09 0 8.406e-09 0 8.409e-09 0.0007 8.412e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.526e-09 0 8.529e-09 0.0007 8.532e-09 0 8.586e-09 0 8.589e-09 0.0007 8.592e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.706e-09 0 8.709e-09 0.0007 8.712e-09 0 8.766e-09 0 8.769e-09 0.0007 8.772e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 8.886e-09 0 8.889e-09 0.0007 8.892e-09 0 8.946e-09 0 8.949e-09 0.0007 8.952e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.066e-09 0 9.069e-09 0.0007 9.072e-09 0 9.126e-09 0 9.129e-09 0.0007 9.132e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.246e-09 0 9.249e-09 0.0007 9.252e-09 0 9.306e-09 0 9.309e-09 0.0007 9.312e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.426e-09 0 9.429e-09 0.0007 9.432e-09 0 9.486e-09 0 9.489e-09 0.0007 9.492e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.606e-09 0 9.609e-09 0.0007 9.612e-09 0 9.666e-09 0 9.669e-09 0.0007 9.672e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.786e-09 0 9.789e-09 0.0007 9.792e-09 0 9.846e-09 0 9.849e-09 0.0007 9.852e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 9.966e-09 0 9.969e-09 0.0007 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0007 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0007 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0007 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0007 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0007 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0007 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0007 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0007 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0007 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0007 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0007 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0007 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0007 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0007 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0007 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0007 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0007 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0007 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0007 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0007 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0007 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0007 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0007 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0007 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0007 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0007 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0007 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0007 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0007 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0007 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0007 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0007 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0007 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0007 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0007 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0007 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0007 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0007 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0007 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0007 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0007 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0007 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0007 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0007 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0007 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0007 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0007 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0007 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0007 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0007 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0007 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0007 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0007 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0007 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0007 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0007 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0007 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0007 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0007 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0007 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0007 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0007 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0007 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0007 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0007 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0007 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0007 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0007 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0007 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0007 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0007 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0007 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0007 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0007 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0007 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0007 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0007 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0007 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0007 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0007 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0007 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0007 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0007 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0007 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0007 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0007 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0007 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0007 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0007 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0007 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0007 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0007 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0007 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0007 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0007 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0007 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0007 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0007 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0007 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0007 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0007 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0007 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0007 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0007 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0007 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0007 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0007 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0007 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0007 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0007 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0007 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0007 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0007 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0007 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0007 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0007 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0007 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0007 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0007 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0007 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0007 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0007 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0007 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0007 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0007 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0007 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0007 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0007 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0007 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0007 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0007 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0007 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0007 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0007 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0007 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0007 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0007 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0007 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0007 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0007 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0007 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0007 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0007 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0007 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0007 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0007 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0007 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0007 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0007 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0007 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0007 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0007 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0007 2.3892e-08 0)
L_DFF_IP1_01|1 IP1_0_OUT _DFF_IP1_01|A1  2.067833848e-12
L_DFF_IP1_01|2 _DFF_IP1_01|A1 _DFF_IP1_01|A2  4.135667696e-12
L_DFF_IP1_01|3 _DFF_IP1_01|A3 _DFF_IP1_01|A4  8.271335392e-12
L_DFF_IP1_01|T D01 _DFF_IP1_01|T1  2.067833848e-12
L_DFF_IP1_01|4 _DFF_IP1_01|T1 _DFF_IP1_01|T2  4.135667696e-12
L_DFF_IP1_01|5 _DFF_IP1_01|A4 _DFF_IP1_01|Q1  4.135667696e-12
L_DFF_IP1_01|6 _DFF_IP1_01|Q1 IP1_1_OUT  2.067833848e-12
ID02|T 0 D02  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 6.6e-11 0 6.9e-11 0.0007 7.2e-11 0 1.26e-10 0 1.29e-10 0.0007 1.32e-10 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 2.46e-10 0 2.49e-10 0.0007 2.52e-10 0 3.06e-10 0 3.09e-10 0.0007 3.12e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 4.26e-10 0 4.29e-10 0.0007 4.32e-10 0 4.86e-10 0 4.89e-10 0.0007 4.92e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 6.06e-10 0 6.09e-10 0.0007 6.12e-10 0 6.66e-10 0 6.69e-10 0.0007 6.72e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 7.86e-10 0 7.89e-10 0.0007 7.92e-10 0 8.46e-10 0 8.49e-10 0.0007 8.52e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 9.66e-10 0 9.69e-10 0.0007 9.72e-10 0 1.026e-09 0 1.029e-09 0.0007 1.032e-09 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.146e-09 0 1.149e-09 0.0007 1.152e-09 0 1.206e-09 0 1.209e-09 0.0007 1.212e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.326e-09 0 1.329e-09 0.0007 1.332e-09 0 1.386e-09 0 1.389e-09 0.0007 1.392e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.506e-09 0 1.509e-09 0.0007 1.512e-09 0 1.566e-09 0 1.569e-09 0.0007 1.572e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.686e-09 0 1.689e-09 0.0007 1.692e-09 0 1.746e-09 0 1.749e-09 0.0007 1.752e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.866e-09 0 1.869e-09 0.0007 1.872e-09 0 1.926e-09 0 1.929e-09 0.0007 1.932e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.046e-09 0 2.049e-09 0.0007 2.052e-09 0 2.106e-09 0 2.109e-09 0.0007 2.112e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.226e-09 0 2.229e-09 0.0007 2.232e-09 0 2.286e-09 0 2.289e-09 0.0007 2.292e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.406e-09 0 2.409e-09 0.0007 2.412e-09 0 2.466e-09 0 2.469e-09 0.0007 2.472e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.586e-09 0 2.589e-09 0.0007 2.592e-09 0 2.646e-09 0 2.649e-09 0.0007 2.652e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.766e-09 0 2.769e-09 0.0007 2.772e-09 0 2.826e-09 0 2.829e-09 0.0007 2.832e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 2.946e-09 0 2.949e-09 0.0007 2.952e-09 0 3.006e-09 0 3.009e-09 0.0007 3.012e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.126e-09 0 3.129e-09 0.0007 3.132e-09 0 3.186e-09 0 3.189e-09 0.0007 3.192e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.306e-09 0 3.309e-09 0.0007 3.312e-09 0 3.366e-09 0 3.369e-09 0.0007 3.372e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.486e-09 0 3.489e-09 0.0007 3.492e-09 0 3.546e-09 0 3.549e-09 0.0007 3.552e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.666e-09 0 3.669e-09 0.0007 3.672e-09 0 3.726e-09 0 3.729e-09 0.0007 3.732e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.846e-09 0 3.849e-09 0.0007 3.852e-09 0 3.906e-09 0 3.909e-09 0.0007 3.912e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.026e-09 0 4.029e-09 0.0007 4.032e-09 0 4.086e-09 0 4.089e-09 0.0007 4.092e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.206e-09 0 4.209e-09 0.0007 4.212e-09 0 4.266e-09 0 4.269e-09 0.0007 4.272e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.386e-09 0 4.389e-09 0.0007 4.392e-09 0 4.446e-09 0 4.449e-09 0.0007 4.452e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.566e-09 0 4.569e-09 0.0007 4.572e-09 0 4.626e-09 0 4.629e-09 0.0007 4.632e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.746e-09 0 4.749e-09 0.0007 4.752e-09 0 4.806e-09 0 4.809e-09 0.0007 4.812e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 4.926e-09 0 4.929e-09 0.0007 4.932e-09 0 4.986e-09 0 4.989e-09 0.0007 4.992e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.106e-09 0 5.109e-09 0.0007 5.112e-09 0 5.166e-09 0 5.169e-09 0.0007 5.172e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.286e-09 0 5.289e-09 0.0007 5.292e-09 0 5.346e-09 0 5.349e-09 0.0007 5.352e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.466e-09 0 5.469e-09 0.0007 5.472e-09 0 5.526e-09 0 5.529e-09 0.0007 5.532e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.646e-09 0 5.649e-09 0.0007 5.652e-09 0 5.706e-09 0 5.709e-09 0.0007 5.712e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.826e-09 0 5.829e-09 0.0007 5.832e-09 0 5.886e-09 0 5.889e-09 0.0007 5.892e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.006e-09 0 6.009e-09 0.0007 6.012e-09 0 6.066e-09 0 6.069e-09 0.0007 6.072e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.186e-09 0 6.189e-09 0.0007 6.192e-09 0 6.246e-09 0 6.249e-09 0.0007 6.252e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.366e-09 0 6.369e-09 0.0007 6.372e-09 0 6.426e-09 0 6.429e-09 0.0007 6.432e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.546e-09 0 6.549e-09 0.0007 6.552e-09 0 6.606e-09 0 6.609e-09 0.0007 6.612e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.726e-09 0 6.729e-09 0.0007 6.732e-09 0 6.786e-09 0 6.789e-09 0.0007 6.792e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 6.906e-09 0 6.909e-09 0.0007 6.912e-09 0 6.966e-09 0 6.969e-09 0.0007 6.972e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.086e-09 0 7.089e-09 0.0007 7.092e-09 0 7.146e-09 0 7.149e-09 0.0007 7.152e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.266e-09 0 7.269e-09 0.0007 7.272e-09 0 7.326e-09 0 7.329e-09 0.0007 7.332e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.446e-09 0 7.449e-09 0.0007 7.452e-09 0 7.506e-09 0 7.509e-09 0.0007 7.512e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.626e-09 0 7.629e-09 0.0007 7.632e-09 0 7.686e-09 0 7.689e-09 0.0007 7.692e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.806e-09 0 7.809e-09 0.0007 7.812e-09 0 7.866e-09 0 7.869e-09 0.0007 7.872e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 7.986e-09 0 7.989e-09 0.0007 7.992e-09 0 8.046e-09 0 8.049e-09 0.0007 8.052e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.166e-09 0 8.169e-09 0.0007 8.172e-09 0 8.226e-09 0 8.229e-09 0.0007 8.232e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.346e-09 0 8.349e-09 0.0007 8.352e-09 0 8.406e-09 0 8.409e-09 0.0007 8.412e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.526e-09 0 8.529e-09 0.0007 8.532e-09 0 8.586e-09 0 8.589e-09 0.0007 8.592e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.706e-09 0 8.709e-09 0.0007 8.712e-09 0 8.766e-09 0 8.769e-09 0.0007 8.772e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 8.886e-09 0 8.889e-09 0.0007 8.892e-09 0 8.946e-09 0 8.949e-09 0.0007 8.952e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.066e-09 0 9.069e-09 0.0007 9.072e-09 0 9.126e-09 0 9.129e-09 0.0007 9.132e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.246e-09 0 9.249e-09 0.0007 9.252e-09 0 9.306e-09 0 9.309e-09 0.0007 9.312e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.426e-09 0 9.429e-09 0.0007 9.432e-09 0 9.486e-09 0 9.489e-09 0.0007 9.492e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.606e-09 0 9.609e-09 0.0007 9.612e-09 0 9.666e-09 0 9.669e-09 0.0007 9.672e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.786e-09 0 9.789e-09 0.0007 9.792e-09 0 9.846e-09 0 9.849e-09 0.0007 9.852e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 9.966e-09 0 9.969e-09 0.0007 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0007 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0007 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0007 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0007 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0007 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0007 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0007 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0007 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0007 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0007 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0007 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0007 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0007 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0007 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0007 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0007 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0007 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0007 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0007 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0007 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0007 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0007 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0007 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0007 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0007 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0007 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0007 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0007 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0007 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0007 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0007 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0007 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0007 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0007 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0007 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0007 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0007 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0007 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0007 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0007 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0007 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0007 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0007 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0007 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0007 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0007 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0007 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0007 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0007 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0007 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0007 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0007 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0007 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0007 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0007 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0007 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0007 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0007 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0007 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0007 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0007 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0007 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0007 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0007 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0007 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0007 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0007 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0007 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0007 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0007 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0007 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0007 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0007 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0007 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0007 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0007 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0007 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0007 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0007 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0007 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0007 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0007 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0007 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0007 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0007 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0007 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0007 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0007 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0007 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0007 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0007 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0007 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0007 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0007 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0007 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0007 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0007 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0007 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0007 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0007 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0007 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0007 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0007 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0007 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0007 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0007 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0007 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0007 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0007 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0007 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0007 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0007 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0007 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0007 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0007 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0007 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0007 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0007 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0007 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0007 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0007 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0007 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0007 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0007 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0007 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0007 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0007 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0007 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0007 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0007 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0007 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0007 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0007 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0007 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0007 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0007 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0007 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0007 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0007 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0007 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0007 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0007 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0007 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0007 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0007 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0007 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0007 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0007 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0007 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0007 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0007 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0007 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0007 2.3892e-08 0)
L_DFF_IP2_01|1 IP2_0_OUT _DFF_IP2_01|A1  2.067833848e-12
L_DFF_IP2_01|2 _DFF_IP2_01|A1 _DFF_IP2_01|A2  4.135667696e-12
L_DFF_IP2_01|3 _DFF_IP2_01|A3 _DFF_IP2_01|A4  8.271335392e-12
L_DFF_IP2_01|T D02 _DFF_IP2_01|T1  2.067833848e-12
L_DFF_IP2_01|4 _DFF_IP2_01|T1 _DFF_IP2_01|T2  4.135667696e-12
L_DFF_IP2_01|5 _DFF_IP2_01|A4 _DFF_IP2_01|Q1  4.135667696e-12
L_DFF_IP2_01|6 _DFF_IP2_01|Q1 IP2_1_OUT  2.067833848e-12
ID03|T 0 D03  PWL(0 0 6e-12 0 9e-12 0.0007 1.2e-11 0 6.6e-11 0 6.9e-11 0.0007 7.2e-11 0 1.26e-10 0 1.29e-10 0.0007 1.32e-10 0 1.86e-10 0 1.89e-10 0.0007 1.92e-10 0 2.46e-10 0 2.49e-10 0.0007 2.52e-10 0 3.06e-10 0 3.09e-10 0.0007 3.12e-10 0 3.66e-10 0 3.69e-10 0.0007 3.72e-10 0 4.26e-10 0 4.29e-10 0.0007 4.32e-10 0 4.86e-10 0 4.89e-10 0.0007 4.92e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 6.06e-10 0 6.09e-10 0.0007 6.12e-10 0 6.66e-10 0 6.69e-10 0.0007 6.72e-10 0 7.26e-10 0 7.29e-10 0.0007 7.32e-10 0 7.86e-10 0 7.89e-10 0.0007 7.92e-10 0 8.46e-10 0 8.49e-10 0.0007 8.52e-10 0 9.06e-10 0 9.09e-10 0.0007 9.12e-10 0 9.66e-10 0 9.69e-10 0.0007 9.72e-10 0 1.026e-09 0 1.029e-09 0.0007 1.032e-09 0 1.086e-09 0 1.089e-09 0.0007 1.092e-09 0 1.146e-09 0 1.149e-09 0.0007 1.152e-09 0 1.206e-09 0 1.209e-09 0.0007 1.212e-09 0 1.266e-09 0 1.269e-09 0.0007 1.272e-09 0 1.326e-09 0 1.329e-09 0.0007 1.332e-09 0 1.386e-09 0 1.389e-09 0.0007 1.392e-09 0 1.446e-09 0 1.449e-09 0.0007 1.452e-09 0 1.506e-09 0 1.509e-09 0.0007 1.512e-09 0 1.566e-09 0 1.569e-09 0.0007 1.572e-09 0 1.626e-09 0 1.629e-09 0.0007 1.632e-09 0 1.686e-09 0 1.689e-09 0.0007 1.692e-09 0 1.746e-09 0 1.749e-09 0.0007 1.752e-09 0 1.806e-09 0 1.809e-09 0.0007 1.812e-09 0 1.866e-09 0 1.869e-09 0.0007 1.872e-09 0 1.926e-09 0 1.929e-09 0.0007 1.932e-09 0 1.986e-09 0 1.989e-09 0.0007 1.992e-09 0 2.046e-09 0 2.049e-09 0.0007 2.052e-09 0 2.106e-09 0 2.109e-09 0.0007 2.112e-09 0 2.166e-09 0 2.169e-09 0.0007 2.172e-09 0 2.226e-09 0 2.229e-09 0.0007 2.232e-09 0 2.286e-09 0 2.289e-09 0.0007 2.292e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.406e-09 0 2.409e-09 0.0007 2.412e-09 0 2.466e-09 0 2.469e-09 0.0007 2.472e-09 0 2.526e-09 0 2.529e-09 0.0007 2.532e-09 0 2.586e-09 0 2.589e-09 0.0007 2.592e-09 0 2.646e-09 0 2.649e-09 0.0007 2.652e-09 0 2.706e-09 0 2.709e-09 0.0007 2.712e-09 0 2.766e-09 0 2.769e-09 0.0007 2.772e-09 0 2.826e-09 0 2.829e-09 0.0007 2.832e-09 0 2.886e-09 0 2.889e-09 0.0007 2.892e-09 0 2.946e-09 0 2.949e-09 0.0007 2.952e-09 0 3.006e-09 0 3.009e-09 0.0007 3.012e-09 0 3.066e-09 0 3.069e-09 0.0007 3.072e-09 0 3.126e-09 0 3.129e-09 0.0007 3.132e-09 0 3.186e-09 0 3.189e-09 0.0007 3.192e-09 0 3.246e-09 0 3.249e-09 0.0007 3.252e-09 0 3.306e-09 0 3.309e-09 0.0007 3.312e-09 0 3.366e-09 0 3.369e-09 0.0007 3.372e-09 0 3.426e-09 0 3.429e-09 0.0007 3.432e-09 0 3.486e-09 0 3.489e-09 0.0007 3.492e-09 0 3.546e-09 0 3.549e-09 0.0007 3.552e-09 0 3.606e-09 0 3.609e-09 0.0007 3.612e-09 0 3.666e-09 0 3.669e-09 0.0007 3.672e-09 0 3.726e-09 0 3.729e-09 0.0007 3.732e-09 0 3.786e-09 0 3.789e-09 0.0007 3.792e-09 0 3.846e-09 0 3.849e-09 0.0007 3.852e-09 0 3.906e-09 0 3.909e-09 0.0007 3.912e-09 0 3.966e-09 0 3.969e-09 0.0007 3.972e-09 0 4.026e-09 0 4.029e-09 0.0007 4.032e-09 0 4.086e-09 0 4.089e-09 0.0007 4.092e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.206e-09 0 4.209e-09 0.0007 4.212e-09 0 4.266e-09 0 4.269e-09 0.0007 4.272e-09 0 4.326e-09 0 4.329e-09 0.0007 4.332e-09 0 4.386e-09 0 4.389e-09 0.0007 4.392e-09 0 4.446e-09 0 4.449e-09 0.0007 4.452e-09 0 4.506e-09 0 4.509e-09 0.0007 4.512e-09 0 4.566e-09 0 4.569e-09 0.0007 4.572e-09 0 4.626e-09 0 4.629e-09 0.0007 4.632e-09 0 4.686e-09 0 4.689e-09 0.0007 4.692e-09 0 4.746e-09 0 4.749e-09 0.0007 4.752e-09 0 4.806e-09 0 4.809e-09 0.0007 4.812e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 4.926e-09 0 4.929e-09 0.0007 4.932e-09 0 4.986e-09 0 4.989e-09 0.0007 4.992e-09 0 5.046e-09 0 5.049e-09 0.0007 5.052e-09 0 5.106e-09 0 5.109e-09 0.0007 5.112e-09 0 5.166e-09 0 5.169e-09 0.0007 5.172e-09 0 5.226e-09 0 5.229e-09 0.0007 5.232e-09 0 5.286e-09 0 5.289e-09 0.0007 5.292e-09 0 5.346e-09 0 5.349e-09 0.0007 5.352e-09 0 5.406e-09 0 5.409e-09 0.0007 5.412e-09 0 5.466e-09 0 5.469e-09 0.0007 5.472e-09 0 5.526e-09 0 5.529e-09 0.0007 5.532e-09 0 5.586e-09 0 5.589e-09 0.0007 5.592e-09 0 5.646e-09 0 5.649e-09 0.0007 5.652e-09 0 5.706e-09 0 5.709e-09 0.0007 5.712e-09 0 5.766e-09 0 5.769e-09 0.0007 5.772e-09 0 5.826e-09 0 5.829e-09 0.0007 5.832e-09 0 5.886e-09 0 5.889e-09 0.0007 5.892e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.006e-09 0 6.009e-09 0.0007 6.012e-09 0 6.066e-09 0 6.069e-09 0.0007 6.072e-09 0 6.126e-09 0 6.129e-09 0.0007 6.132e-09 0 6.186e-09 0 6.189e-09 0.0007 6.192e-09 0 6.246e-09 0 6.249e-09 0.0007 6.252e-09 0 6.306e-09 0 6.309e-09 0.0007 6.312e-09 0 6.366e-09 0 6.369e-09 0.0007 6.372e-09 0 6.426e-09 0 6.429e-09 0.0007 6.432e-09 0 6.486e-09 0 6.489e-09 0.0007 6.492e-09 0 6.546e-09 0 6.549e-09 0.0007 6.552e-09 0 6.606e-09 0 6.609e-09 0.0007 6.612e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.726e-09 0 6.729e-09 0.0007 6.732e-09 0 6.786e-09 0 6.789e-09 0.0007 6.792e-09 0 6.846e-09 0 6.849e-09 0.0007 6.852e-09 0 6.906e-09 0 6.909e-09 0.0007 6.912e-09 0 6.966e-09 0 6.969e-09 0.0007 6.972e-09 0 7.026e-09 0 7.029e-09 0.0007 7.032e-09 0 7.086e-09 0 7.089e-09 0.0007 7.092e-09 0 7.146e-09 0 7.149e-09 0.0007 7.152e-09 0 7.206e-09 0 7.209e-09 0.0007 7.212e-09 0 7.266e-09 0 7.269e-09 0.0007 7.272e-09 0 7.326e-09 0 7.329e-09 0.0007 7.332e-09 0 7.386e-09 0 7.389e-09 0.0007 7.392e-09 0 7.446e-09 0 7.449e-09 0.0007 7.452e-09 0 7.506e-09 0 7.509e-09 0.0007 7.512e-09 0 7.566e-09 0 7.569e-09 0.0007 7.572e-09 0 7.626e-09 0 7.629e-09 0.0007 7.632e-09 0 7.686e-09 0 7.689e-09 0.0007 7.692e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.806e-09 0 7.809e-09 0.0007 7.812e-09 0 7.866e-09 0 7.869e-09 0.0007 7.872e-09 0 7.926e-09 0 7.929e-09 0.0007 7.932e-09 0 7.986e-09 0 7.989e-09 0.0007 7.992e-09 0 8.046e-09 0 8.049e-09 0.0007 8.052e-09 0 8.106e-09 0 8.109e-09 0.0007 8.112e-09 0 8.166e-09 0 8.169e-09 0.0007 8.172e-09 0 8.226e-09 0 8.229e-09 0.0007 8.232e-09 0 8.286e-09 0 8.289e-09 0.0007 8.292e-09 0 8.346e-09 0 8.349e-09 0.0007 8.352e-09 0 8.406e-09 0 8.409e-09 0.0007 8.412e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.526e-09 0 8.529e-09 0.0007 8.532e-09 0 8.586e-09 0 8.589e-09 0.0007 8.592e-09 0 8.646e-09 0 8.649e-09 0.0007 8.652e-09 0 8.706e-09 0 8.709e-09 0.0007 8.712e-09 0 8.766e-09 0 8.769e-09 0.0007 8.772e-09 0 8.826e-09 0 8.829e-09 0.0007 8.832e-09 0 8.886e-09 0 8.889e-09 0.0007 8.892e-09 0 8.946e-09 0 8.949e-09 0.0007 8.952e-09 0 9.006e-09 0 9.009e-09 0.0007 9.012e-09 0 9.066e-09 0 9.069e-09 0.0007 9.072e-09 0 9.126e-09 0 9.129e-09 0.0007 9.132e-09 0 9.186e-09 0 9.189e-09 0.0007 9.192e-09 0 9.246e-09 0 9.249e-09 0.0007 9.252e-09 0 9.306e-09 0 9.309e-09 0.0007 9.312e-09 0 9.366e-09 0 9.369e-09 0.0007 9.372e-09 0 9.426e-09 0 9.429e-09 0.0007 9.432e-09 0 9.486e-09 0 9.489e-09 0.0007 9.492e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.606e-09 0 9.609e-09 0.0007 9.612e-09 0 9.666e-09 0 9.669e-09 0.0007 9.672e-09 0 9.726e-09 0 9.729e-09 0.0007 9.732e-09 0 9.786e-09 0 9.789e-09 0.0007 9.792e-09 0 9.846e-09 0 9.849e-09 0.0007 9.852e-09 0 9.906e-09 0 9.909e-09 0.0007 9.912e-09 0 9.966e-09 0 9.969e-09 0.0007 9.972e-09 0 1.0026e-08 0 1.0029e-08 0.0007 1.0032e-08 0 1.0086e-08 0 1.0089e-08 0.0007 1.0092e-08 0 1.0146e-08 0 1.0149e-08 0.0007 1.0152e-08 0 1.0206e-08 0 1.0209e-08 0.0007 1.0212e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.0326e-08 0 1.0329e-08 0.0007 1.0332e-08 0 1.0386e-08 0 1.0389e-08 0.0007 1.0392e-08 0 1.0446e-08 0 1.0449e-08 0.0007 1.0452e-08 0 1.0506e-08 0 1.0509e-08 0.0007 1.0512e-08 0 1.0566e-08 0 1.0569e-08 0.0007 1.0572e-08 0 1.0626e-08 0 1.0629e-08 0.0007 1.0632e-08 0 1.0686e-08 0 1.0689e-08 0.0007 1.0692e-08 0 1.0746e-08 0 1.0749e-08 0.0007 1.0752e-08 0 1.0806e-08 0 1.0809e-08 0.0007 1.0812e-08 0 1.0866e-08 0 1.0869e-08 0.0007 1.0872e-08 0 1.0926e-08 0 1.0929e-08 0.0007 1.0932e-08 0 1.0986e-08 0 1.0989e-08 0.0007 1.0992e-08 0 1.1046e-08 0 1.1049e-08 0.0007 1.1052e-08 0 1.1106e-08 0 1.1109e-08 0.0007 1.1112e-08 0 1.1166e-08 0 1.1169e-08 0.0007 1.1172e-08 0 1.1226e-08 0 1.1229e-08 0.0007 1.1232e-08 0 1.1286e-08 0 1.1289e-08 0.0007 1.1292e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1406e-08 0 1.1409e-08 0.0007 1.1412e-08 0 1.1466e-08 0 1.1469e-08 0.0007 1.1472e-08 0 1.1526e-08 0 1.1529e-08 0.0007 1.1532e-08 0 1.1586e-08 0 1.1589e-08 0.0007 1.1592e-08 0 1.1646e-08 0 1.1649e-08 0.0007 1.1652e-08 0 1.1706e-08 0 1.1709e-08 0.0007 1.1712e-08 0 1.1766e-08 0 1.1769e-08 0.0007 1.1772e-08 0 1.1826e-08 0 1.1829e-08 0.0007 1.1832e-08 0 1.1886e-08 0 1.1889e-08 0.0007 1.1892e-08 0 1.1946e-08 0 1.1949e-08 0.0007 1.1952e-08 0 1.2006e-08 0 1.2009e-08 0.0007 1.2012e-08 0 1.2066e-08 0 1.2069e-08 0.0007 1.2072e-08 0 1.2126e-08 0 1.2129e-08 0.0007 1.2132e-08 0 1.2186e-08 0 1.2189e-08 0.0007 1.2192e-08 0 1.2246e-08 0 1.2249e-08 0.0007 1.2252e-08 0 1.2306e-08 0 1.2309e-08 0.0007 1.2312e-08 0 1.2366e-08 0 1.2369e-08 0.0007 1.2372e-08 0 1.2426e-08 0 1.2429e-08 0.0007 1.2432e-08 0 1.2486e-08 0 1.2489e-08 0.0007 1.2492e-08 0 1.2546e-08 0 1.2549e-08 0.0007 1.2552e-08 0 1.2606e-08 0 1.2609e-08 0.0007 1.2612e-08 0 1.2666e-08 0 1.2669e-08 0.0007 1.2672e-08 0 1.2726e-08 0 1.2729e-08 0.0007 1.2732e-08 0 1.2786e-08 0 1.2789e-08 0.0007 1.2792e-08 0 1.2846e-08 0 1.2849e-08 0.0007 1.2852e-08 0 1.2906e-08 0 1.2909e-08 0.0007 1.2912e-08 0 1.2966e-08 0 1.2969e-08 0.0007 1.2972e-08 0 1.3026e-08 0 1.3029e-08 0.0007 1.3032e-08 0 1.3086e-08 0 1.3089e-08 0.0007 1.3092e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3206e-08 0 1.3209e-08 0.0007 1.3212e-08 0 1.3266e-08 0 1.3269e-08 0.0007 1.3272e-08 0 1.3326e-08 0 1.3329e-08 0.0007 1.3332e-08 0 1.3386e-08 0 1.3389e-08 0.0007 1.3392e-08 0 1.3446e-08 0 1.3449e-08 0.0007 1.3452e-08 0 1.3506e-08 0 1.3509e-08 0.0007 1.3512e-08 0 1.3566e-08 0 1.3569e-08 0.0007 1.3572e-08 0 1.3626e-08 0 1.3629e-08 0.0007 1.3632e-08 0 1.3686e-08 0 1.3689e-08 0.0007 1.3692e-08 0 1.3746e-08 0 1.3749e-08 0.0007 1.3752e-08 0 1.3806e-08 0 1.3809e-08 0.0007 1.3812e-08 0 1.3866e-08 0 1.3869e-08 0.0007 1.3872e-08 0 1.3926e-08 0 1.3929e-08 0.0007 1.3932e-08 0 1.3986e-08 0 1.3989e-08 0.0007 1.3992e-08 0 1.4046e-08 0 1.4049e-08 0.0007 1.4052e-08 0 1.4106e-08 0 1.4109e-08 0.0007 1.4112e-08 0 1.4166e-08 0 1.4169e-08 0.0007 1.4172e-08 0 1.4226e-08 0 1.4229e-08 0.0007 1.4232e-08 0 1.4286e-08 0 1.4289e-08 0.0007 1.4292e-08 0 1.4346e-08 0 1.4349e-08 0.0007 1.4352e-08 0 1.4406e-08 0 1.4409e-08 0.0007 1.4412e-08 0 1.4466e-08 0 1.4469e-08 0.0007 1.4472e-08 0 1.4526e-08 0 1.4529e-08 0.0007 1.4532e-08 0 1.4586e-08 0 1.4589e-08 0.0007 1.4592e-08 0 1.4646e-08 0 1.4649e-08 0.0007 1.4652e-08 0 1.4706e-08 0 1.4709e-08 0.0007 1.4712e-08 0 1.4766e-08 0 1.4769e-08 0.0007 1.4772e-08 0 1.4826e-08 0 1.4829e-08 0.0007 1.4832e-08 0 1.4886e-08 0 1.4889e-08 0.0007 1.4892e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5066e-08 0 1.5069e-08 0.0007 1.5072e-08 0 1.5126e-08 0 1.5129e-08 0.0007 1.5132e-08 0 1.5186e-08 0 1.5189e-08 0.0007 1.5192e-08 0 1.5246e-08 0 1.5249e-08 0.0007 1.5252e-08 0 1.5306e-08 0 1.5309e-08 0.0007 1.5312e-08 0 1.5366e-08 0 1.5369e-08 0.0007 1.5372e-08 0 1.5426e-08 0 1.5429e-08 0.0007 1.5432e-08 0 1.5486e-08 0 1.5489e-08 0.0007 1.5492e-08 0 1.5546e-08 0 1.5549e-08 0.0007 1.5552e-08 0 1.5606e-08 0 1.5609e-08 0.0007 1.5612e-08 0 1.5666e-08 0 1.5669e-08 0.0007 1.5672e-08 0 1.5726e-08 0 1.5729e-08 0.0007 1.5732e-08 0 1.5786e-08 0 1.5789e-08 0.0007 1.5792e-08 0 1.5846e-08 0 1.5849e-08 0.0007 1.5852e-08 0 1.5906e-08 0 1.5909e-08 0.0007 1.5912e-08 0 1.5966e-08 0 1.5969e-08 0.0007 1.5972e-08 0 1.6026e-08 0 1.6029e-08 0.0007 1.6032e-08 0 1.6086e-08 0 1.6089e-08 0.0007 1.6092e-08 0 1.6146e-08 0 1.6149e-08 0.0007 1.6152e-08 0 1.6206e-08 0 1.6209e-08 0.0007 1.6212e-08 0 1.6266e-08 0 1.6269e-08 0.0007 1.6272e-08 0 1.6326e-08 0 1.6329e-08 0.0007 1.6332e-08 0 1.6386e-08 0 1.6389e-08 0.0007 1.6392e-08 0 1.6446e-08 0 1.6449e-08 0.0007 1.6452e-08 0 1.6506e-08 0 1.6509e-08 0.0007 1.6512e-08 0 1.6566e-08 0 1.6569e-08 0.0007 1.6572e-08 0 1.6626e-08 0 1.6629e-08 0.0007 1.6632e-08 0 1.6686e-08 0 1.6689e-08 0.0007 1.6692e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6806e-08 0 1.6809e-08 0.0007 1.6812e-08 0 1.6866e-08 0 1.6869e-08 0.0007 1.6872e-08 0 1.6926e-08 0 1.6929e-08 0.0007 1.6932e-08 0 1.6986e-08 0 1.6989e-08 0.0007 1.6992e-08 0 1.7046e-08 0 1.7049e-08 0.0007 1.7052e-08 0 1.7106e-08 0 1.7109e-08 0.0007 1.7112e-08 0 1.7166e-08 0 1.7169e-08 0.0007 1.7172e-08 0 1.7226e-08 0 1.7229e-08 0.0007 1.7232e-08 0 1.7286e-08 0 1.7289e-08 0.0007 1.7292e-08 0 1.7346e-08 0 1.7349e-08 0.0007 1.7352e-08 0 1.7406e-08 0 1.7409e-08 0.0007 1.7412e-08 0 1.7466e-08 0 1.7469e-08 0.0007 1.7472e-08 0 1.7526e-08 0 1.7529e-08 0.0007 1.7532e-08 0 1.7586e-08 0 1.7589e-08 0.0007 1.7592e-08 0 1.7646e-08 0 1.7649e-08 0.0007 1.7652e-08 0 1.7706e-08 0 1.7709e-08 0.0007 1.7712e-08 0 1.7766e-08 0 1.7769e-08 0.0007 1.7772e-08 0 1.7826e-08 0 1.7829e-08 0.0007 1.7832e-08 0 1.7886e-08 0 1.7889e-08 0.0007 1.7892e-08 0 1.7946e-08 0 1.7949e-08 0.0007 1.7952e-08 0 1.8006e-08 0 1.8009e-08 0.0007 1.8012e-08 0 1.8066e-08 0 1.8069e-08 0.0007 1.8072e-08 0 1.8126e-08 0 1.8129e-08 0.0007 1.8132e-08 0 1.8186e-08 0 1.8189e-08 0.0007 1.8192e-08 0 1.8246e-08 0 1.8249e-08 0.0007 1.8252e-08 0 1.8306e-08 0 1.8309e-08 0.0007 1.8312e-08 0 1.8366e-08 0 1.8369e-08 0.0007 1.8372e-08 0 1.8426e-08 0 1.8429e-08 0.0007 1.8432e-08 0 1.8486e-08 0 1.8489e-08 0.0007 1.8492e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8606e-08 0 1.8609e-08 0.0007 1.8612e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8726e-08 0 1.8729e-08 0.0007 1.8732e-08 0 1.8786e-08 0 1.8789e-08 0.0007 1.8792e-08 0 1.8846e-08 0 1.8849e-08 0.0007 1.8852e-08 0 1.8906e-08 0 1.8909e-08 0.0007 1.8912e-08 0 1.8966e-08 0 1.8969e-08 0.0007 1.8972e-08 0 1.9026e-08 0 1.9029e-08 0.0007 1.9032e-08 0 1.9086e-08 0 1.9089e-08 0.0007 1.9092e-08 0 1.9146e-08 0 1.9149e-08 0.0007 1.9152e-08 0 1.9206e-08 0 1.9209e-08 0.0007 1.9212e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9326e-08 0 1.9329e-08 0.0007 1.9332e-08 0 1.9386e-08 0 1.9389e-08 0.0007 1.9392e-08 0 1.9446e-08 0 1.9449e-08 0.0007 1.9452e-08 0 1.9506e-08 0 1.9509e-08 0.0007 1.9512e-08 0 1.9566e-08 0 1.9569e-08 0.0007 1.9572e-08 0 1.9626e-08 0 1.9629e-08 0.0007 1.9632e-08 0 1.9686e-08 0 1.9689e-08 0.0007 1.9692e-08 0 1.9746e-08 0 1.9749e-08 0.0007 1.9752e-08 0 1.9806e-08 0 1.9809e-08 0.0007 1.9812e-08 0 1.9866e-08 0 1.9869e-08 0.0007 1.9872e-08 0 1.9926e-08 0 1.9929e-08 0.0007 1.9932e-08 0 1.9986e-08 0 1.9989e-08 0.0007 1.9992e-08 0 2.0046e-08 0 2.0049e-08 0.0007 2.0052e-08 0 2.0106e-08 0 2.0109e-08 0.0007 2.0112e-08 0 2.0166e-08 0 2.0169e-08 0.0007 2.0172e-08 0 2.0226e-08 0 2.0229e-08 0.0007 2.0232e-08 0 2.0286e-08 0 2.0289e-08 0.0007 2.0292e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0406e-08 0 2.0409e-08 0.0007 2.0412e-08 0 2.0466e-08 0 2.0469e-08 0.0007 2.0472e-08 0 2.0526e-08 0 2.0529e-08 0.0007 2.0532e-08 0 2.0586e-08 0 2.0589e-08 0.0007 2.0592e-08 0 2.0646e-08 0 2.0649e-08 0.0007 2.0652e-08 0 2.0706e-08 0 2.0709e-08 0.0007 2.0712e-08 0 2.0766e-08 0 2.0769e-08 0.0007 2.0772e-08 0 2.0826e-08 0 2.0829e-08 0.0007 2.0832e-08 0 2.0886e-08 0 2.0889e-08 0.0007 2.0892e-08 0 2.0946e-08 0 2.0949e-08 0.0007 2.0952e-08 0 2.1006e-08 0 2.1009e-08 0.0007 2.1012e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1126e-08 0 2.1129e-08 0.0007 2.1132e-08 0 2.1186e-08 0 2.1189e-08 0.0007 2.1192e-08 0 2.1246e-08 0 2.1249e-08 0.0007 2.1252e-08 0 2.1306e-08 0 2.1309e-08 0.0007 2.1312e-08 0 2.1366e-08 0 2.1369e-08 0.0007 2.1372e-08 0 2.1426e-08 0 2.1429e-08 0.0007 2.1432e-08 0 2.1486e-08 0 2.1489e-08 0.0007 2.1492e-08 0 2.1546e-08 0 2.1549e-08 0.0007 2.1552e-08 0 2.1606e-08 0 2.1609e-08 0.0007 2.1612e-08 0 2.1666e-08 0 2.1669e-08 0.0007 2.1672e-08 0 2.1726e-08 0 2.1729e-08 0.0007 2.1732e-08 0 2.1786e-08 0 2.1789e-08 0.0007 2.1792e-08 0 2.1846e-08 0 2.1849e-08 0.0007 2.1852e-08 0 2.1906e-08 0 2.1909e-08 0.0007 2.1912e-08 0 2.1966e-08 0 2.1969e-08 0.0007 2.1972e-08 0 2.2026e-08 0 2.2029e-08 0.0007 2.2032e-08 0 2.2086e-08 0 2.2089e-08 0.0007 2.2092e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2206e-08 0 2.2209e-08 0.0007 2.2212e-08 0 2.2266e-08 0 2.2269e-08 0.0007 2.2272e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2386e-08 0 2.2389e-08 0.0007 2.2392e-08 0 2.2446e-08 0 2.2449e-08 0.0007 2.2452e-08 0 2.2506e-08 0 2.2509e-08 0.0007 2.2512e-08 0 2.2566e-08 0 2.2569e-08 0.0007 2.2572e-08 0 2.2626e-08 0 2.2629e-08 0.0007 2.2632e-08 0 2.2686e-08 0 2.2689e-08 0.0007 2.2692e-08 0 2.2746e-08 0 2.2749e-08 0.0007 2.2752e-08 0 2.2806e-08 0 2.2809e-08 0.0007 2.2812e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.2926e-08 0 2.2929e-08 0.0007 2.2932e-08 0 2.2986e-08 0 2.2989e-08 0.0007 2.2992e-08 0 2.3046e-08 0 2.3049e-08 0.0007 2.3052e-08 0 2.3106e-08 0 2.3109e-08 0.0007 2.3112e-08 0 2.3166e-08 0 2.3169e-08 0.0007 2.3172e-08 0 2.3226e-08 0 2.3229e-08 0.0007 2.3232e-08 0 2.3286e-08 0 2.3289e-08 0.0007 2.3292e-08 0 2.3346e-08 0 2.3349e-08 0.0007 2.3352e-08 0 2.3406e-08 0 2.3409e-08 0.0007 2.3412e-08 0 2.3466e-08 0 2.3469e-08 0.0007 2.3472e-08 0 2.3526e-08 0 2.3529e-08 0.0007 2.3532e-08 0 2.3586e-08 0 2.3589e-08 0.0007 2.3592e-08 0 2.3646e-08 0 2.3649e-08 0.0007 2.3652e-08 0 2.3706e-08 0 2.3709e-08 0.0007 2.3712e-08 0 2.3766e-08 0 2.3769e-08 0.0007 2.3772e-08 0 2.3826e-08 0 2.3829e-08 0.0007 2.3832e-08 0 2.3886e-08 0 2.3889e-08 0.0007 2.3892e-08 0)
L_DFF_IP3_01|1 IP3_0_OUT _DFF_IP3_01|A1  2.067833848e-12
L_DFF_IP3_01|2 _DFF_IP3_01|A1 _DFF_IP3_01|A2  4.135667696e-12
L_DFF_IP3_01|3 _DFF_IP3_01|A3 _DFF_IP3_01|A4  8.271335392e-12
L_DFF_IP3_01|T D03 _DFF_IP3_01|T1  2.067833848e-12
L_DFF_IP3_01|4 _DFF_IP3_01|T1 _DFF_IP3_01|T2  4.135667696e-12
L_DFF_IP3_01|5 _DFF_IP3_01|A4 _DFF_IP3_01|Q1  4.135667696e-12
L_DFF_IP3_01|6 _DFF_IP3_01|Q1 IP3_1_OUT  2.067833848e-12
IT08|T 0 T08  PWL(0 0 3e-12 0 6e-12 0.0014 9e-12 0 6.3e-11 0 6.6e-11 0.0014 6.9e-11 0 1.23e-10 0 1.26e-10 0.0014 1.29e-10 0 1.83e-10 0 1.86e-10 0.0014 1.89e-10 0 2.43e-10 0 2.46e-10 0.0014 2.49e-10 0 3.03e-10 0 3.06e-10 0.0014 3.09e-10 0 3.63e-10 0 3.66e-10 0.0014 3.69e-10 0 4.23e-10 0 4.26e-10 0.0014 4.29e-10 0 4.83e-10 0 4.86e-10 0.0014 4.89e-10 0 5.43e-10 0 5.46e-10 0.0014 5.49e-10 0 6.03e-10 0 6.06e-10 0.0014 6.09e-10 0 6.63e-10 0 6.66e-10 0.0014 6.69e-10 0 7.23e-10 0 7.26e-10 0.0014 7.29e-10 0 7.83e-10 0 7.86e-10 0.0014 7.89e-10 0 8.43e-10 0 8.46e-10 0.0014 8.49e-10 0 9.03e-10 0 9.06e-10 0.0014 9.09e-10 0 9.63e-10 0 9.66e-10 0.0014 9.69e-10 0 1.023e-09 0 1.026e-09 0.0014 1.029e-09 0 1.083e-09 0 1.086e-09 0.0014 1.089e-09 0 1.143e-09 0 1.146e-09 0.0014 1.149e-09 0 1.203e-09 0 1.206e-09 0.0014 1.209e-09 0 1.263e-09 0 1.266e-09 0.0014 1.269e-09 0 1.323e-09 0 1.326e-09 0.0014 1.329e-09 0 1.383e-09 0 1.386e-09 0.0014 1.389e-09 0 1.443e-09 0 1.446e-09 0.0014 1.449e-09 0 1.503e-09 0 1.506e-09 0.0014 1.509e-09 0 1.563e-09 0 1.566e-09 0.0014 1.569e-09 0 1.623e-09 0 1.626e-09 0.0014 1.629e-09 0 1.683e-09 0 1.686e-09 0.0014 1.689e-09 0 1.743e-09 0 1.746e-09 0.0014 1.749e-09 0 1.803e-09 0 1.806e-09 0.0014 1.809e-09 0 1.863e-09 0 1.866e-09 0.0014 1.869e-09 0 1.923e-09 0 1.926e-09 0.0014 1.929e-09 0 1.983e-09 0 1.986e-09 0.0014 1.989e-09 0 2.043e-09 0 2.046e-09 0.0014 2.049e-09 0 2.103e-09 0 2.106e-09 0.0014 2.109e-09 0 2.163e-09 0 2.166e-09 0.0014 2.169e-09 0 2.223e-09 0 2.226e-09 0.0014 2.229e-09 0 2.283e-09 0 2.286e-09 0.0014 2.289e-09 0 2.343e-09 0 2.346e-09 0.0014 2.349e-09 0 2.403e-09 0 2.406e-09 0.0014 2.409e-09 0 2.463e-09 0 2.466e-09 0.0014 2.469e-09 0 2.523e-09 0 2.526e-09 0.0014 2.529e-09 0 2.583e-09 0 2.586e-09 0.0014 2.589e-09 0 2.643e-09 0 2.646e-09 0.0014 2.649e-09 0 2.703e-09 0 2.706e-09 0.0014 2.709e-09 0 2.763e-09 0 2.766e-09 0.0014 2.769e-09 0 2.823e-09 0 2.826e-09 0.0014 2.829e-09 0 2.883e-09 0 2.886e-09 0.0014 2.889e-09 0 2.943e-09 0 2.946e-09 0.0014 2.949e-09 0 3.003e-09 0 3.006e-09 0.0014 3.009e-09 0 3.063e-09 0 3.066e-09 0.0014 3.069e-09 0 3.123e-09 0 3.126e-09 0.0014 3.129e-09 0 3.183e-09 0 3.186e-09 0.0014 3.189e-09 0 3.243e-09 0 3.246e-09 0.0014 3.249e-09 0 3.303e-09 0 3.306e-09 0.0014 3.309e-09 0 3.363e-09 0 3.366e-09 0.0014 3.369e-09 0 3.423e-09 0 3.426e-09 0.0014 3.429e-09 0 3.483e-09 0 3.486e-09 0.0014 3.489e-09 0 3.543e-09 0 3.546e-09 0.0014 3.549e-09 0 3.603e-09 0 3.606e-09 0.0014 3.609e-09 0 3.663e-09 0 3.666e-09 0.0014 3.669e-09 0 3.723e-09 0 3.726e-09 0.0014 3.729e-09 0 3.783e-09 0 3.786e-09 0.0014 3.789e-09 0 3.843e-09 0 3.846e-09 0.0014 3.849e-09 0 3.903e-09 0 3.906e-09 0.0014 3.909e-09 0 3.963e-09 0 3.966e-09 0.0014 3.969e-09 0 4.023e-09 0 4.026e-09 0.0014 4.029e-09 0 4.083e-09 0 4.086e-09 0.0014 4.089e-09 0 4.143e-09 0 4.146e-09 0.0014 4.149e-09 0 4.203e-09 0 4.206e-09 0.0014 4.209e-09 0 4.263e-09 0 4.266e-09 0.0014 4.269e-09 0 4.323e-09 0 4.326e-09 0.0014 4.329e-09 0 4.383e-09 0 4.386e-09 0.0014 4.389e-09 0 4.443e-09 0 4.446e-09 0.0014 4.449e-09 0 4.503e-09 0 4.506e-09 0.0014 4.509e-09 0 4.563e-09 0 4.566e-09 0.0014 4.569e-09 0 4.623e-09 0 4.626e-09 0.0014 4.629e-09 0 4.683e-09 0 4.686e-09 0.0014 4.689e-09 0 4.743e-09 0 4.746e-09 0.0014 4.749e-09 0 4.803e-09 0 4.806e-09 0.0014 4.809e-09 0 4.863e-09 0 4.866e-09 0.0014 4.869e-09 0 4.923e-09 0 4.926e-09 0.0014 4.929e-09 0 4.983e-09 0 4.986e-09 0.0014 4.989e-09 0 5.043e-09 0 5.046e-09 0.0014 5.049e-09 0 5.103e-09 0 5.106e-09 0.0014 5.109e-09 0 5.163e-09 0 5.166e-09 0.0014 5.169e-09 0 5.223e-09 0 5.226e-09 0.0014 5.229e-09 0 5.283e-09 0 5.286e-09 0.0014 5.289e-09 0 5.343e-09 0 5.346e-09 0.0014 5.349e-09 0 5.403e-09 0 5.406e-09 0.0014 5.409e-09 0 5.463e-09 0 5.466e-09 0.0014 5.469e-09 0 5.523e-09 0 5.526e-09 0.0014 5.529e-09 0 5.583e-09 0 5.586e-09 0.0014 5.589e-09 0 5.643e-09 0 5.646e-09 0.0014 5.649e-09 0 5.703e-09 0 5.706e-09 0.0014 5.709e-09 0 5.763e-09 0 5.766e-09 0.0014 5.769e-09 0 5.823e-09 0 5.826e-09 0.0014 5.829e-09 0 5.883e-09 0 5.886e-09 0.0014 5.889e-09 0 5.943e-09 0 5.946e-09 0.0014 5.949e-09 0 6.003e-09 0 6.006e-09 0.0014 6.009e-09 0 6.063e-09 0 6.066e-09 0.0014 6.069e-09 0 6.123e-09 0 6.126e-09 0.0014 6.129e-09 0 6.183e-09 0 6.186e-09 0.0014 6.189e-09 0 6.243e-09 0 6.246e-09 0.0014 6.249e-09 0 6.303e-09 0 6.306e-09 0.0014 6.309e-09 0 6.363e-09 0 6.366e-09 0.0014 6.369e-09 0 6.423e-09 0 6.426e-09 0.0014 6.429e-09 0 6.483e-09 0 6.486e-09 0.0014 6.489e-09 0 6.543e-09 0 6.546e-09 0.0014 6.549e-09 0 6.603e-09 0 6.606e-09 0.0014 6.609e-09 0 6.663e-09 0 6.666e-09 0.0014 6.669e-09 0 6.723e-09 0 6.726e-09 0.0014 6.729e-09 0 6.783e-09 0 6.786e-09 0.0014 6.789e-09 0 6.843e-09 0 6.846e-09 0.0014 6.849e-09 0 6.903e-09 0 6.906e-09 0.0014 6.909e-09 0 6.963e-09 0 6.966e-09 0.0014 6.969e-09 0 7.023e-09 0 7.026e-09 0.0014 7.029e-09 0 7.083e-09 0 7.086e-09 0.0014 7.089e-09 0 7.143e-09 0 7.146e-09 0.0014 7.149e-09 0 7.203e-09 0 7.206e-09 0.0014 7.209e-09 0 7.263e-09 0 7.266e-09 0.0014 7.269e-09 0 7.323e-09 0 7.326e-09 0.0014 7.329e-09 0 7.383e-09 0 7.386e-09 0.0014 7.389e-09 0 7.443e-09 0 7.446e-09 0.0014 7.449e-09 0 7.503e-09 0 7.506e-09 0.0014 7.509e-09 0 7.563e-09 0 7.566e-09 0.0014 7.569e-09 0 7.623e-09 0 7.626e-09 0.0014 7.629e-09 0 7.683e-09 0 7.686e-09 0.0014 7.689e-09 0 7.743e-09 0 7.746e-09 0.0014 7.749e-09 0 7.803e-09 0 7.806e-09 0.0014 7.809e-09 0 7.863e-09 0 7.866e-09 0.0014 7.869e-09 0 7.923e-09 0 7.926e-09 0.0014 7.929e-09 0 7.983e-09 0 7.986e-09 0.0014 7.989e-09 0 8.043e-09 0 8.046e-09 0.0014 8.049e-09 0 8.103e-09 0 8.106e-09 0.0014 8.109e-09 0 8.163e-09 0 8.166e-09 0.0014 8.169e-09 0 8.223e-09 0 8.226e-09 0.0014 8.229e-09 0 8.283e-09 0 8.286e-09 0.0014 8.289e-09 0 8.343e-09 0 8.346e-09 0.0014 8.349e-09 0 8.403e-09 0 8.406e-09 0.0014 8.409e-09 0 8.463e-09 0 8.466e-09 0.0014 8.469e-09 0 8.523e-09 0 8.526e-09 0.0014 8.529e-09 0 8.583e-09 0 8.586e-09 0.0014 8.589e-09 0 8.643e-09 0 8.646e-09 0.0014 8.649e-09 0 8.703e-09 0 8.706e-09 0.0014 8.709e-09 0 8.763e-09 0 8.766e-09 0.0014 8.769e-09 0 8.823e-09 0 8.826e-09 0.0014 8.829e-09 0 8.883e-09 0 8.886e-09 0.0014 8.889e-09 0 8.943e-09 0 8.946e-09 0.0014 8.949e-09 0 9.003e-09 0 9.006e-09 0.0014 9.009e-09 0 9.063e-09 0 9.066e-09 0.0014 9.069e-09 0 9.123e-09 0 9.126e-09 0.0014 9.129e-09 0 9.183e-09 0 9.186e-09 0.0014 9.189e-09 0 9.243e-09 0 9.246e-09 0.0014 9.249e-09 0 9.303e-09 0 9.306e-09 0.0014 9.309e-09 0 9.363e-09 0 9.366e-09 0.0014 9.369e-09 0 9.423e-09 0 9.426e-09 0.0014 9.429e-09 0 9.483e-09 0 9.486e-09 0.0014 9.489e-09 0 9.543e-09 0 9.546e-09 0.0014 9.549e-09 0 9.603e-09 0 9.606e-09 0.0014 9.609e-09 0 9.663e-09 0 9.666e-09 0.0014 9.669e-09 0 9.723e-09 0 9.726e-09 0.0014 9.729e-09 0 9.783e-09 0 9.786e-09 0.0014 9.789e-09 0 9.843e-09 0 9.846e-09 0.0014 9.849e-09 0 9.903e-09 0 9.906e-09 0.0014 9.909e-09 0 9.963e-09 0 9.966e-09 0.0014 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0014 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0014 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0014 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0014 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0014 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0014 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0014 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0014 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0014 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0014 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0014 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0014 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0014 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0014 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0014 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0014 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0014 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0014 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0014 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0014 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0014 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0014 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0014 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0014 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0014 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0014 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0014 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0014 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0014 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0014 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0014 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0014 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0014 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0014 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0014 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0014 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0014 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0014 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0014 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0014 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0014 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0014 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0014 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0014 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0014 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0014 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0014 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0014 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0014 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0014 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0014 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0014 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0014 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0014 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0014 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0014 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0014 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0014 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0014 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0014 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0014 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0014 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0014 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0014 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0014 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0014 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0014 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0014 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0014 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0014 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0014 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0014 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0014 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0014 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0014 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0014 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0014 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0014 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0014 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0014 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0014 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0014 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0014 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0014 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0014 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0014 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0014 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0014 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0014 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0014 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0014 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0014 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0014 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0014 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0014 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0014 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0014 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0014 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0014 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0014 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0014 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0014 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0014 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0014 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0014 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0014 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0014 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0014 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0014 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0014 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0014 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0014 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0014 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0014 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0014 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0014 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0014 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0014 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0014 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0014 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0014 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0014 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0014 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0014 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0014 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0014 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0014 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0014 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0014 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0014 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0014 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0014 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0014 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0014 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0014 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0014 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0014 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0014 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0014 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0014 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0014 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0014 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0014 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0014 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0014 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0014 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0014 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0014 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0014 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0014 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0014 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0014 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0014 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0014 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0014 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0014 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0014 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0014 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0014 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0014 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0014 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0014 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0014 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0014 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0014 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0014 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0014 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0014 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0014 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0014 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0014 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0014 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0014 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0014 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0014 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0014 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0014 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0014 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0014 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0014 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0014 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0014 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0014 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0014 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0014 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0014 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0014 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0014 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0014 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0014 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0014 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0014 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0014 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0014 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0014 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0014 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0014 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0014 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0014 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0014 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0014 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0014 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0014 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0014 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0014 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0014 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0014 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0014 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0014 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0014 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0014 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0014 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0014 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0014 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0014 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0014 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0014 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0014 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0014 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0014 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0014 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0014 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0014 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0014 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0014 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0014 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0014 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0014 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0014 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0014 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0014 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0014 2.3889e-08 0)
IT09|T 0 T09  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 6.3e-11 0 6.6e-11 0.0007 6.9e-11 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 1.83e-10 0 1.86e-10 0.0007 1.89e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.03e-10 0 3.06e-10 0.0007 3.09e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.23e-10 0 4.26e-10 0.0007 4.29e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 5.43e-10 0 5.46e-10 0.0007 5.49e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 6.63e-10 0 6.66e-10 0.0007 6.69e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 7.83e-10 0 7.86e-10 0.0007 7.89e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.03e-10 0 9.06e-10 0.0007 9.09e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.023e-09 0 1.026e-09 0.0007 1.029e-09 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.143e-09 0 1.146e-09 0.0007 1.149e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.263e-09 0 1.266e-09 0.0007 1.269e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.383e-09 0 1.386e-09 0.0007 1.389e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.503e-09 0 1.506e-09 0.0007 1.509e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.623e-09 0 1.626e-09 0.0007 1.629e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.743e-09 0 1.746e-09 0.0007 1.749e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.863e-09 0 1.866e-09 0.0007 1.869e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 1.983e-09 0 1.986e-09 0.0007 1.989e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.103e-09 0 2.106e-09 0.0007 2.109e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.223e-09 0 2.226e-09 0.0007 2.229e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.343e-09 0 2.346e-09 0.0007 2.349e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.463e-09 0 2.466e-09 0.0007 2.469e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.583e-09 0 2.586e-09 0.0007 2.589e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.703e-09 0 2.706e-09 0.0007 2.709e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.823e-09 0 2.826e-09 0.0007 2.829e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 2.943e-09 0 2.946e-09 0.0007 2.949e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.183e-09 0 3.186e-09 0.0007 3.189e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.303e-09 0 3.306e-09 0.0007 3.309e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.423e-09 0 3.426e-09 0.0007 3.429e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.543e-09 0 3.546e-09 0.0007 3.549e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.663e-09 0 3.666e-09 0.0007 3.669e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.783e-09 0 3.786e-09 0.0007 3.789e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.903e-09 0 3.906e-09 0.0007 3.909e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.023e-09 0 4.026e-09 0.0007 4.029e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.143e-09 0 4.146e-09 0.0007 4.149e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.383e-09 0 4.386e-09 0.0007 4.389e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.503e-09 0 4.506e-09 0.0007 4.509e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.623e-09 0 4.626e-09 0.0007 4.629e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.743e-09 0 4.746e-09 0.0007 4.749e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.863e-09 0 4.866e-09 0.0007 4.869e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 4.983e-09 0 4.986e-09 0.0007 4.989e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.103e-09 0 5.106e-09 0.0007 5.109e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.223e-09 0 5.226e-09 0.0007 5.229e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.343e-09 0 5.346e-09 0.0007 5.349e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.583e-09 0 5.586e-09 0.0007 5.589e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.703e-09 0 5.706e-09 0.0007 5.709e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.823e-09 0 5.826e-09 0.0007 5.829e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 5.943e-09 0 5.946e-09 0.0007 5.949e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.183e-09 0 6.186e-09 0.0007 6.189e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.303e-09 0 6.306e-09 0.0007 6.309e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.423e-09 0 6.426e-09 0.0007 6.429e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.543e-09 0 6.546e-09 0.0007 6.549e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.663e-09 0 6.666e-09 0.0007 6.669e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.783e-09 0 6.786e-09 0.0007 6.789e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.903e-09 0 6.906e-09 0.0007 6.909e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.023e-09 0 7.026e-09 0.0007 7.029e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.143e-09 0 7.146e-09 0.0007 7.149e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.263e-09 0 7.266e-09 0.0007 7.269e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.383e-09 0 7.386e-09 0.0007 7.389e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.503e-09 0 7.506e-09 0.0007 7.509e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.623e-09 0 7.626e-09 0.0007 7.629e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.743e-09 0 7.746e-09 0.0007 7.749e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 7.983e-09 0 7.986e-09 0.0007 7.989e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.103e-09 0 8.106e-09 0.0007 8.109e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.223e-09 0 8.226e-09 0.0007 8.229e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.343e-09 0 8.346e-09 0.0007 8.349e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.583e-09 0 8.586e-09 0.0007 8.589e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.703e-09 0 8.706e-09 0.0007 8.709e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.823e-09 0 8.826e-09 0.0007 8.829e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 8.943e-09 0 8.946e-09 0.0007 8.949e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.183e-09 0 9.186e-09 0.0007 9.189e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.303e-09 0 9.306e-09 0.0007 9.309e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.423e-09 0 9.426e-09 0.0007 9.429e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.543e-09 0 9.546e-09 0.0007 9.549e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.663e-09 0 9.666e-09 0.0007 9.669e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.783e-09 0 9.786e-09 0.0007 9.789e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.903e-09 0 9.906e-09 0.0007 9.909e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0007 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0007 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0007 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0007 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0007 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0007 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0007 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0007 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0007 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0007 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0007 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0007 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0007 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0007 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0007 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0007 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0007 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0007 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0007 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0007 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0007 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0007 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0007 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0007 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0007 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0007 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0007 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0007 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0007 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0007 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0007 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0007 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0007 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0007 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0007 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0007 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0007 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0007 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0007 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0007 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0007 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0007 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0007 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0007 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0007 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0007 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0007 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0007 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0007 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0007 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0007 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0007 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0007 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0007 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0007 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0007 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0007 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0007 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0007 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0007 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0007 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0007 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0007 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0007 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0007 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0007 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0007 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0007 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0007 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0007 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0007 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0007 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0007 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0007 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0007 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0007 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0007 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0007 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0007 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0007 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0007 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0007 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0007 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0007 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0007 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0007 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0007 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0007 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0007 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0007 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0007 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0007 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0007 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0007 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0)
L_PG1_12|1 G1_1_TO1 _PG1_12|A1  2.067833848e-12
L_PG1_12|2 _PG1_12|A1 _PG1_12|A2  4.135667696e-12
L_PG1_12|3 _PG1_12|A3 _PG1_12|A4  8.271335392e-12
L_PG1_12|T T09 _PG1_12|T1  2.067833848e-12
L_PG1_12|4 _PG1_12|T1 _PG1_12|T2  4.135667696e-12
L_PG1_12|5 _PG1_12|A4 _PG1_12|Q1  4.135667696e-12
L_PG1_12|6 _PG1_12|Q1 G1_2  2.067833848e-12
IT10|T 0 T10  PWL(0 0 3e-12 0 6e-12 0.0014 9e-12 0 6.3e-11 0 6.6e-11 0.0014 6.9e-11 0 1.23e-10 0 1.26e-10 0.0014 1.29e-10 0 1.83e-10 0 1.86e-10 0.0014 1.89e-10 0 2.43e-10 0 2.46e-10 0.0014 2.49e-10 0 3.03e-10 0 3.06e-10 0.0014 3.09e-10 0 3.63e-10 0 3.66e-10 0.0014 3.69e-10 0 4.23e-10 0 4.26e-10 0.0014 4.29e-10 0 4.83e-10 0 4.86e-10 0.0014 4.89e-10 0 5.43e-10 0 5.46e-10 0.0014 5.49e-10 0 6.03e-10 0 6.06e-10 0.0014 6.09e-10 0 6.63e-10 0 6.66e-10 0.0014 6.69e-10 0 7.23e-10 0 7.26e-10 0.0014 7.29e-10 0 7.83e-10 0 7.86e-10 0.0014 7.89e-10 0 8.43e-10 0 8.46e-10 0.0014 8.49e-10 0 9.03e-10 0 9.06e-10 0.0014 9.09e-10 0 9.63e-10 0 9.66e-10 0.0014 9.69e-10 0 1.023e-09 0 1.026e-09 0.0014 1.029e-09 0 1.083e-09 0 1.086e-09 0.0014 1.089e-09 0 1.143e-09 0 1.146e-09 0.0014 1.149e-09 0 1.203e-09 0 1.206e-09 0.0014 1.209e-09 0 1.263e-09 0 1.266e-09 0.0014 1.269e-09 0 1.323e-09 0 1.326e-09 0.0014 1.329e-09 0 1.383e-09 0 1.386e-09 0.0014 1.389e-09 0 1.443e-09 0 1.446e-09 0.0014 1.449e-09 0 1.503e-09 0 1.506e-09 0.0014 1.509e-09 0 1.563e-09 0 1.566e-09 0.0014 1.569e-09 0 1.623e-09 0 1.626e-09 0.0014 1.629e-09 0 1.683e-09 0 1.686e-09 0.0014 1.689e-09 0 1.743e-09 0 1.746e-09 0.0014 1.749e-09 0 1.803e-09 0 1.806e-09 0.0014 1.809e-09 0 1.863e-09 0 1.866e-09 0.0014 1.869e-09 0 1.923e-09 0 1.926e-09 0.0014 1.929e-09 0 1.983e-09 0 1.986e-09 0.0014 1.989e-09 0 2.043e-09 0 2.046e-09 0.0014 2.049e-09 0 2.103e-09 0 2.106e-09 0.0014 2.109e-09 0 2.163e-09 0 2.166e-09 0.0014 2.169e-09 0 2.223e-09 0 2.226e-09 0.0014 2.229e-09 0 2.283e-09 0 2.286e-09 0.0014 2.289e-09 0 2.343e-09 0 2.346e-09 0.0014 2.349e-09 0 2.403e-09 0 2.406e-09 0.0014 2.409e-09 0 2.463e-09 0 2.466e-09 0.0014 2.469e-09 0 2.523e-09 0 2.526e-09 0.0014 2.529e-09 0 2.583e-09 0 2.586e-09 0.0014 2.589e-09 0 2.643e-09 0 2.646e-09 0.0014 2.649e-09 0 2.703e-09 0 2.706e-09 0.0014 2.709e-09 0 2.763e-09 0 2.766e-09 0.0014 2.769e-09 0 2.823e-09 0 2.826e-09 0.0014 2.829e-09 0 2.883e-09 0 2.886e-09 0.0014 2.889e-09 0 2.943e-09 0 2.946e-09 0.0014 2.949e-09 0 3.003e-09 0 3.006e-09 0.0014 3.009e-09 0 3.063e-09 0 3.066e-09 0.0014 3.069e-09 0 3.123e-09 0 3.126e-09 0.0014 3.129e-09 0 3.183e-09 0 3.186e-09 0.0014 3.189e-09 0 3.243e-09 0 3.246e-09 0.0014 3.249e-09 0 3.303e-09 0 3.306e-09 0.0014 3.309e-09 0 3.363e-09 0 3.366e-09 0.0014 3.369e-09 0 3.423e-09 0 3.426e-09 0.0014 3.429e-09 0 3.483e-09 0 3.486e-09 0.0014 3.489e-09 0 3.543e-09 0 3.546e-09 0.0014 3.549e-09 0 3.603e-09 0 3.606e-09 0.0014 3.609e-09 0 3.663e-09 0 3.666e-09 0.0014 3.669e-09 0 3.723e-09 0 3.726e-09 0.0014 3.729e-09 0 3.783e-09 0 3.786e-09 0.0014 3.789e-09 0 3.843e-09 0 3.846e-09 0.0014 3.849e-09 0 3.903e-09 0 3.906e-09 0.0014 3.909e-09 0 3.963e-09 0 3.966e-09 0.0014 3.969e-09 0 4.023e-09 0 4.026e-09 0.0014 4.029e-09 0 4.083e-09 0 4.086e-09 0.0014 4.089e-09 0 4.143e-09 0 4.146e-09 0.0014 4.149e-09 0 4.203e-09 0 4.206e-09 0.0014 4.209e-09 0 4.263e-09 0 4.266e-09 0.0014 4.269e-09 0 4.323e-09 0 4.326e-09 0.0014 4.329e-09 0 4.383e-09 0 4.386e-09 0.0014 4.389e-09 0 4.443e-09 0 4.446e-09 0.0014 4.449e-09 0 4.503e-09 0 4.506e-09 0.0014 4.509e-09 0 4.563e-09 0 4.566e-09 0.0014 4.569e-09 0 4.623e-09 0 4.626e-09 0.0014 4.629e-09 0 4.683e-09 0 4.686e-09 0.0014 4.689e-09 0 4.743e-09 0 4.746e-09 0.0014 4.749e-09 0 4.803e-09 0 4.806e-09 0.0014 4.809e-09 0 4.863e-09 0 4.866e-09 0.0014 4.869e-09 0 4.923e-09 0 4.926e-09 0.0014 4.929e-09 0 4.983e-09 0 4.986e-09 0.0014 4.989e-09 0 5.043e-09 0 5.046e-09 0.0014 5.049e-09 0 5.103e-09 0 5.106e-09 0.0014 5.109e-09 0 5.163e-09 0 5.166e-09 0.0014 5.169e-09 0 5.223e-09 0 5.226e-09 0.0014 5.229e-09 0 5.283e-09 0 5.286e-09 0.0014 5.289e-09 0 5.343e-09 0 5.346e-09 0.0014 5.349e-09 0 5.403e-09 0 5.406e-09 0.0014 5.409e-09 0 5.463e-09 0 5.466e-09 0.0014 5.469e-09 0 5.523e-09 0 5.526e-09 0.0014 5.529e-09 0 5.583e-09 0 5.586e-09 0.0014 5.589e-09 0 5.643e-09 0 5.646e-09 0.0014 5.649e-09 0 5.703e-09 0 5.706e-09 0.0014 5.709e-09 0 5.763e-09 0 5.766e-09 0.0014 5.769e-09 0 5.823e-09 0 5.826e-09 0.0014 5.829e-09 0 5.883e-09 0 5.886e-09 0.0014 5.889e-09 0 5.943e-09 0 5.946e-09 0.0014 5.949e-09 0 6.003e-09 0 6.006e-09 0.0014 6.009e-09 0 6.063e-09 0 6.066e-09 0.0014 6.069e-09 0 6.123e-09 0 6.126e-09 0.0014 6.129e-09 0 6.183e-09 0 6.186e-09 0.0014 6.189e-09 0 6.243e-09 0 6.246e-09 0.0014 6.249e-09 0 6.303e-09 0 6.306e-09 0.0014 6.309e-09 0 6.363e-09 0 6.366e-09 0.0014 6.369e-09 0 6.423e-09 0 6.426e-09 0.0014 6.429e-09 0 6.483e-09 0 6.486e-09 0.0014 6.489e-09 0 6.543e-09 0 6.546e-09 0.0014 6.549e-09 0 6.603e-09 0 6.606e-09 0.0014 6.609e-09 0 6.663e-09 0 6.666e-09 0.0014 6.669e-09 0 6.723e-09 0 6.726e-09 0.0014 6.729e-09 0 6.783e-09 0 6.786e-09 0.0014 6.789e-09 0 6.843e-09 0 6.846e-09 0.0014 6.849e-09 0 6.903e-09 0 6.906e-09 0.0014 6.909e-09 0 6.963e-09 0 6.966e-09 0.0014 6.969e-09 0 7.023e-09 0 7.026e-09 0.0014 7.029e-09 0 7.083e-09 0 7.086e-09 0.0014 7.089e-09 0 7.143e-09 0 7.146e-09 0.0014 7.149e-09 0 7.203e-09 0 7.206e-09 0.0014 7.209e-09 0 7.263e-09 0 7.266e-09 0.0014 7.269e-09 0 7.323e-09 0 7.326e-09 0.0014 7.329e-09 0 7.383e-09 0 7.386e-09 0.0014 7.389e-09 0 7.443e-09 0 7.446e-09 0.0014 7.449e-09 0 7.503e-09 0 7.506e-09 0.0014 7.509e-09 0 7.563e-09 0 7.566e-09 0.0014 7.569e-09 0 7.623e-09 0 7.626e-09 0.0014 7.629e-09 0 7.683e-09 0 7.686e-09 0.0014 7.689e-09 0 7.743e-09 0 7.746e-09 0.0014 7.749e-09 0 7.803e-09 0 7.806e-09 0.0014 7.809e-09 0 7.863e-09 0 7.866e-09 0.0014 7.869e-09 0 7.923e-09 0 7.926e-09 0.0014 7.929e-09 0 7.983e-09 0 7.986e-09 0.0014 7.989e-09 0 8.043e-09 0 8.046e-09 0.0014 8.049e-09 0 8.103e-09 0 8.106e-09 0.0014 8.109e-09 0 8.163e-09 0 8.166e-09 0.0014 8.169e-09 0 8.223e-09 0 8.226e-09 0.0014 8.229e-09 0 8.283e-09 0 8.286e-09 0.0014 8.289e-09 0 8.343e-09 0 8.346e-09 0.0014 8.349e-09 0 8.403e-09 0 8.406e-09 0.0014 8.409e-09 0 8.463e-09 0 8.466e-09 0.0014 8.469e-09 0 8.523e-09 0 8.526e-09 0.0014 8.529e-09 0 8.583e-09 0 8.586e-09 0.0014 8.589e-09 0 8.643e-09 0 8.646e-09 0.0014 8.649e-09 0 8.703e-09 0 8.706e-09 0.0014 8.709e-09 0 8.763e-09 0 8.766e-09 0.0014 8.769e-09 0 8.823e-09 0 8.826e-09 0.0014 8.829e-09 0 8.883e-09 0 8.886e-09 0.0014 8.889e-09 0 8.943e-09 0 8.946e-09 0.0014 8.949e-09 0 9.003e-09 0 9.006e-09 0.0014 9.009e-09 0 9.063e-09 0 9.066e-09 0.0014 9.069e-09 0 9.123e-09 0 9.126e-09 0.0014 9.129e-09 0 9.183e-09 0 9.186e-09 0.0014 9.189e-09 0 9.243e-09 0 9.246e-09 0.0014 9.249e-09 0 9.303e-09 0 9.306e-09 0.0014 9.309e-09 0 9.363e-09 0 9.366e-09 0.0014 9.369e-09 0 9.423e-09 0 9.426e-09 0.0014 9.429e-09 0 9.483e-09 0 9.486e-09 0.0014 9.489e-09 0 9.543e-09 0 9.546e-09 0.0014 9.549e-09 0 9.603e-09 0 9.606e-09 0.0014 9.609e-09 0 9.663e-09 0 9.666e-09 0.0014 9.669e-09 0 9.723e-09 0 9.726e-09 0.0014 9.729e-09 0 9.783e-09 0 9.786e-09 0.0014 9.789e-09 0 9.843e-09 0 9.846e-09 0.0014 9.849e-09 0 9.903e-09 0 9.906e-09 0.0014 9.909e-09 0 9.963e-09 0 9.966e-09 0.0014 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0014 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0014 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0014 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0014 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0014 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0014 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0014 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0014 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0014 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0014 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0014 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0014 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0014 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0014 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0014 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0014 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0014 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0014 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0014 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0014 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0014 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0014 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0014 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0014 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0014 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0014 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0014 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0014 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0014 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0014 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0014 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0014 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0014 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0014 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0014 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0014 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0014 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0014 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0014 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0014 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0014 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0014 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0014 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0014 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0014 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0014 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0014 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0014 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0014 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0014 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0014 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0014 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0014 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0014 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0014 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0014 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0014 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0014 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0014 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0014 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0014 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0014 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0014 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0014 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0014 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0014 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0014 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0014 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0014 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0014 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0014 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0014 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0014 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0014 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0014 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0014 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0014 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0014 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0014 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0014 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0014 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0014 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0014 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0014 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0014 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0014 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0014 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0014 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0014 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0014 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0014 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0014 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0014 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0014 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0014 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0014 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0014 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0014 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0014 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0014 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0014 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0014 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0014 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0014 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0014 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0014 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0014 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0014 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0014 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0014 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0014 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0014 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0014 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0014 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0014 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0014 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0014 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0014 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0014 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0014 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0014 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0014 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0014 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0014 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0014 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0014 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0014 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0014 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0014 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0014 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0014 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0014 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0014 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0014 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0014 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0014 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0014 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0014 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0014 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0014 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0014 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0014 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0014 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0014 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0014 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0014 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0014 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0014 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0014 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0014 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0014 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0014 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0014 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0014 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0014 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0014 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0014 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0014 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0014 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0014 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0014 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0014 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0014 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0014 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0014 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0014 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0014 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0014 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0014 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0014 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0014 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0014 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0014 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0014 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0014 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0014 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0014 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0014 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0014 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0014 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0014 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0014 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0014 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0014 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0014 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0014 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0014 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0014 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0014 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0014 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0014 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0014 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0014 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0014 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0014 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0014 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0014 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0014 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0014 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0014 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0014 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0014 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0014 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0014 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0014 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0014 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0014 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0014 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0014 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0014 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0014 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0014 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0014 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0014 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0014 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0014 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0014 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0014 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0014 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0014 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0014 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0014 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0014 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0014 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0014 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0014 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0014 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0014 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0014 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0014 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0014 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0014 2.3889e-08 0)
IT11|T 0 T11  PWL(0 0 3e-12 0 6e-12 0.0014 9e-12 0 6.3e-11 0 6.6e-11 0.0014 6.9e-11 0 1.23e-10 0 1.26e-10 0.0014 1.29e-10 0 1.83e-10 0 1.86e-10 0.0014 1.89e-10 0 2.43e-10 0 2.46e-10 0.0014 2.49e-10 0 3.03e-10 0 3.06e-10 0.0014 3.09e-10 0 3.63e-10 0 3.66e-10 0.0014 3.69e-10 0 4.23e-10 0 4.26e-10 0.0014 4.29e-10 0 4.83e-10 0 4.86e-10 0.0014 4.89e-10 0 5.43e-10 0 5.46e-10 0.0014 5.49e-10 0 6.03e-10 0 6.06e-10 0.0014 6.09e-10 0 6.63e-10 0 6.66e-10 0.0014 6.69e-10 0 7.23e-10 0 7.26e-10 0.0014 7.29e-10 0 7.83e-10 0 7.86e-10 0.0014 7.89e-10 0 8.43e-10 0 8.46e-10 0.0014 8.49e-10 0 9.03e-10 0 9.06e-10 0.0014 9.09e-10 0 9.63e-10 0 9.66e-10 0.0014 9.69e-10 0 1.023e-09 0 1.026e-09 0.0014 1.029e-09 0 1.083e-09 0 1.086e-09 0.0014 1.089e-09 0 1.143e-09 0 1.146e-09 0.0014 1.149e-09 0 1.203e-09 0 1.206e-09 0.0014 1.209e-09 0 1.263e-09 0 1.266e-09 0.0014 1.269e-09 0 1.323e-09 0 1.326e-09 0.0014 1.329e-09 0 1.383e-09 0 1.386e-09 0.0014 1.389e-09 0 1.443e-09 0 1.446e-09 0.0014 1.449e-09 0 1.503e-09 0 1.506e-09 0.0014 1.509e-09 0 1.563e-09 0 1.566e-09 0.0014 1.569e-09 0 1.623e-09 0 1.626e-09 0.0014 1.629e-09 0 1.683e-09 0 1.686e-09 0.0014 1.689e-09 0 1.743e-09 0 1.746e-09 0.0014 1.749e-09 0 1.803e-09 0 1.806e-09 0.0014 1.809e-09 0 1.863e-09 0 1.866e-09 0.0014 1.869e-09 0 1.923e-09 0 1.926e-09 0.0014 1.929e-09 0 1.983e-09 0 1.986e-09 0.0014 1.989e-09 0 2.043e-09 0 2.046e-09 0.0014 2.049e-09 0 2.103e-09 0 2.106e-09 0.0014 2.109e-09 0 2.163e-09 0 2.166e-09 0.0014 2.169e-09 0 2.223e-09 0 2.226e-09 0.0014 2.229e-09 0 2.283e-09 0 2.286e-09 0.0014 2.289e-09 0 2.343e-09 0 2.346e-09 0.0014 2.349e-09 0 2.403e-09 0 2.406e-09 0.0014 2.409e-09 0 2.463e-09 0 2.466e-09 0.0014 2.469e-09 0 2.523e-09 0 2.526e-09 0.0014 2.529e-09 0 2.583e-09 0 2.586e-09 0.0014 2.589e-09 0 2.643e-09 0 2.646e-09 0.0014 2.649e-09 0 2.703e-09 0 2.706e-09 0.0014 2.709e-09 0 2.763e-09 0 2.766e-09 0.0014 2.769e-09 0 2.823e-09 0 2.826e-09 0.0014 2.829e-09 0 2.883e-09 0 2.886e-09 0.0014 2.889e-09 0 2.943e-09 0 2.946e-09 0.0014 2.949e-09 0 3.003e-09 0 3.006e-09 0.0014 3.009e-09 0 3.063e-09 0 3.066e-09 0.0014 3.069e-09 0 3.123e-09 0 3.126e-09 0.0014 3.129e-09 0 3.183e-09 0 3.186e-09 0.0014 3.189e-09 0 3.243e-09 0 3.246e-09 0.0014 3.249e-09 0 3.303e-09 0 3.306e-09 0.0014 3.309e-09 0 3.363e-09 0 3.366e-09 0.0014 3.369e-09 0 3.423e-09 0 3.426e-09 0.0014 3.429e-09 0 3.483e-09 0 3.486e-09 0.0014 3.489e-09 0 3.543e-09 0 3.546e-09 0.0014 3.549e-09 0 3.603e-09 0 3.606e-09 0.0014 3.609e-09 0 3.663e-09 0 3.666e-09 0.0014 3.669e-09 0 3.723e-09 0 3.726e-09 0.0014 3.729e-09 0 3.783e-09 0 3.786e-09 0.0014 3.789e-09 0 3.843e-09 0 3.846e-09 0.0014 3.849e-09 0 3.903e-09 0 3.906e-09 0.0014 3.909e-09 0 3.963e-09 0 3.966e-09 0.0014 3.969e-09 0 4.023e-09 0 4.026e-09 0.0014 4.029e-09 0 4.083e-09 0 4.086e-09 0.0014 4.089e-09 0 4.143e-09 0 4.146e-09 0.0014 4.149e-09 0 4.203e-09 0 4.206e-09 0.0014 4.209e-09 0 4.263e-09 0 4.266e-09 0.0014 4.269e-09 0 4.323e-09 0 4.326e-09 0.0014 4.329e-09 0 4.383e-09 0 4.386e-09 0.0014 4.389e-09 0 4.443e-09 0 4.446e-09 0.0014 4.449e-09 0 4.503e-09 0 4.506e-09 0.0014 4.509e-09 0 4.563e-09 0 4.566e-09 0.0014 4.569e-09 0 4.623e-09 0 4.626e-09 0.0014 4.629e-09 0 4.683e-09 0 4.686e-09 0.0014 4.689e-09 0 4.743e-09 0 4.746e-09 0.0014 4.749e-09 0 4.803e-09 0 4.806e-09 0.0014 4.809e-09 0 4.863e-09 0 4.866e-09 0.0014 4.869e-09 0 4.923e-09 0 4.926e-09 0.0014 4.929e-09 0 4.983e-09 0 4.986e-09 0.0014 4.989e-09 0 5.043e-09 0 5.046e-09 0.0014 5.049e-09 0 5.103e-09 0 5.106e-09 0.0014 5.109e-09 0 5.163e-09 0 5.166e-09 0.0014 5.169e-09 0 5.223e-09 0 5.226e-09 0.0014 5.229e-09 0 5.283e-09 0 5.286e-09 0.0014 5.289e-09 0 5.343e-09 0 5.346e-09 0.0014 5.349e-09 0 5.403e-09 0 5.406e-09 0.0014 5.409e-09 0 5.463e-09 0 5.466e-09 0.0014 5.469e-09 0 5.523e-09 0 5.526e-09 0.0014 5.529e-09 0 5.583e-09 0 5.586e-09 0.0014 5.589e-09 0 5.643e-09 0 5.646e-09 0.0014 5.649e-09 0 5.703e-09 0 5.706e-09 0.0014 5.709e-09 0 5.763e-09 0 5.766e-09 0.0014 5.769e-09 0 5.823e-09 0 5.826e-09 0.0014 5.829e-09 0 5.883e-09 0 5.886e-09 0.0014 5.889e-09 0 5.943e-09 0 5.946e-09 0.0014 5.949e-09 0 6.003e-09 0 6.006e-09 0.0014 6.009e-09 0 6.063e-09 0 6.066e-09 0.0014 6.069e-09 0 6.123e-09 0 6.126e-09 0.0014 6.129e-09 0 6.183e-09 0 6.186e-09 0.0014 6.189e-09 0 6.243e-09 0 6.246e-09 0.0014 6.249e-09 0 6.303e-09 0 6.306e-09 0.0014 6.309e-09 0 6.363e-09 0 6.366e-09 0.0014 6.369e-09 0 6.423e-09 0 6.426e-09 0.0014 6.429e-09 0 6.483e-09 0 6.486e-09 0.0014 6.489e-09 0 6.543e-09 0 6.546e-09 0.0014 6.549e-09 0 6.603e-09 0 6.606e-09 0.0014 6.609e-09 0 6.663e-09 0 6.666e-09 0.0014 6.669e-09 0 6.723e-09 0 6.726e-09 0.0014 6.729e-09 0 6.783e-09 0 6.786e-09 0.0014 6.789e-09 0 6.843e-09 0 6.846e-09 0.0014 6.849e-09 0 6.903e-09 0 6.906e-09 0.0014 6.909e-09 0 6.963e-09 0 6.966e-09 0.0014 6.969e-09 0 7.023e-09 0 7.026e-09 0.0014 7.029e-09 0 7.083e-09 0 7.086e-09 0.0014 7.089e-09 0 7.143e-09 0 7.146e-09 0.0014 7.149e-09 0 7.203e-09 0 7.206e-09 0.0014 7.209e-09 0 7.263e-09 0 7.266e-09 0.0014 7.269e-09 0 7.323e-09 0 7.326e-09 0.0014 7.329e-09 0 7.383e-09 0 7.386e-09 0.0014 7.389e-09 0 7.443e-09 0 7.446e-09 0.0014 7.449e-09 0 7.503e-09 0 7.506e-09 0.0014 7.509e-09 0 7.563e-09 0 7.566e-09 0.0014 7.569e-09 0 7.623e-09 0 7.626e-09 0.0014 7.629e-09 0 7.683e-09 0 7.686e-09 0.0014 7.689e-09 0 7.743e-09 0 7.746e-09 0.0014 7.749e-09 0 7.803e-09 0 7.806e-09 0.0014 7.809e-09 0 7.863e-09 0 7.866e-09 0.0014 7.869e-09 0 7.923e-09 0 7.926e-09 0.0014 7.929e-09 0 7.983e-09 0 7.986e-09 0.0014 7.989e-09 0 8.043e-09 0 8.046e-09 0.0014 8.049e-09 0 8.103e-09 0 8.106e-09 0.0014 8.109e-09 0 8.163e-09 0 8.166e-09 0.0014 8.169e-09 0 8.223e-09 0 8.226e-09 0.0014 8.229e-09 0 8.283e-09 0 8.286e-09 0.0014 8.289e-09 0 8.343e-09 0 8.346e-09 0.0014 8.349e-09 0 8.403e-09 0 8.406e-09 0.0014 8.409e-09 0 8.463e-09 0 8.466e-09 0.0014 8.469e-09 0 8.523e-09 0 8.526e-09 0.0014 8.529e-09 0 8.583e-09 0 8.586e-09 0.0014 8.589e-09 0 8.643e-09 0 8.646e-09 0.0014 8.649e-09 0 8.703e-09 0 8.706e-09 0.0014 8.709e-09 0 8.763e-09 0 8.766e-09 0.0014 8.769e-09 0 8.823e-09 0 8.826e-09 0.0014 8.829e-09 0 8.883e-09 0 8.886e-09 0.0014 8.889e-09 0 8.943e-09 0 8.946e-09 0.0014 8.949e-09 0 9.003e-09 0 9.006e-09 0.0014 9.009e-09 0 9.063e-09 0 9.066e-09 0.0014 9.069e-09 0 9.123e-09 0 9.126e-09 0.0014 9.129e-09 0 9.183e-09 0 9.186e-09 0.0014 9.189e-09 0 9.243e-09 0 9.246e-09 0.0014 9.249e-09 0 9.303e-09 0 9.306e-09 0.0014 9.309e-09 0 9.363e-09 0 9.366e-09 0.0014 9.369e-09 0 9.423e-09 0 9.426e-09 0.0014 9.429e-09 0 9.483e-09 0 9.486e-09 0.0014 9.489e-09 0 9.543e-09 0 9.546e-09 0.0014 9.549e-09 0 9.603e-09 0 9.606e-09 0.0014 9.609e-09 0 9.663e-09 0 9.666e-09 0.0014 9.669e-09 0 9.723e-09 0 9.726e-09 0.0014 9.729e-09 0 9.783e-09 0 9.786e-09 0.0014 9.789e-09 0 9.843e-09 0 9.846e-09 0.0014 9.849e-09 0 9.903e-09 0 9.906e-09 0.0014 9.909e-09 0 9.963e-09 0 9.966e-09 0.0014 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0014 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0014 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0014 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0014 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0014 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0014 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0014 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0014 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0014 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0014 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0014 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0014 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0014 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0014 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0014 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0014 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0014 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0014 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0014 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0014 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0014 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0014 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0014 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0014 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0014 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0014 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0014 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0014 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0014 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0014 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0014 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0014 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0014 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0014 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0014 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0014 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0014 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0014 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0014 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0014 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0014 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0014 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0014 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0014 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0014 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0014 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0014 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0014 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0014 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0014 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0014 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0014 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0014 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0014 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0014 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0014 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0014 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0014 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0014 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0014 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0014 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0014 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0014 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0014 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0014 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0014 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0014 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0014 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0014 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0014 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0014 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0014 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0014 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0014 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0014 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0014 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0014 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0014 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0014 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0014 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0014 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0014 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0014 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0014 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0014 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0014 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0014 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0014 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0014 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0014 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0014 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0014 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0014 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0014 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0014 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0014 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0014 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0014 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0014 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0014 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0014 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0014 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0014 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0014 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0014 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0014 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0014 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0014 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0014 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0014 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0014 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0014 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0014 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0014 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0014 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0014 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0014 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0014 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0014 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0014 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0014 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0014 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0014 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0014 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0014 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0014 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0014 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0014 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0014 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0014 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0014 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0014 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0014 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0014 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0014 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0014 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0014 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0014 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0014 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0014 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0014 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0014 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0014 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0014 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0014 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0014 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0014 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0014 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0014 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0014 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0014 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0014 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0014 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0014 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0014 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0014 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0014 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0014 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0014 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0014 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0014 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0014 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0014 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0014 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0014 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0014 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0014 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0014 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0014 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0014 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0014 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0014 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0014 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0014 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0014 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0014 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0014 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0014 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0014 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0014 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0014 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0014 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0014 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0014 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0014 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0014 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0014 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0014 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0014 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0014 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0014 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0014 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0014 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0014 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0014 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0014 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0014 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0014 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0014 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0014 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0014 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0014 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0014 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0014 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0014 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0014 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0014 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0014 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0014 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0014 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0014 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0014 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0014 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0014 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0014 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0014 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0014 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0014 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0014 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0014 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0014 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0014 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0014 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0014 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0014 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0014 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0014 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0014 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0014 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0014 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0014 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0014 2.3889e-08 0)
ID11|T 0 D11  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 6.3e-11 0 6.6e-11 0.0007 6.9e-11 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 1.83e-10 0 1.86e-10 0.0007 1.89e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.03e-10 0 3.06e-10 0.0007 3.09e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.23e-10 0 4.26e-10 0.0007 4.29e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 5.43e-10 0 5.46e-10 0.0007 5.49e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 6.63e-10 0 6.66e-10 0.0007 6.69e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 7.83e-10 0 7.86e-10 0.0007 7.89e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.03e-10 0 9.06e-10 0.0007 9.09e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.023e-09 0 1.026e-09 0.0007 1.029e-09 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.143e-09 0 1.146e-09 0.0007 1.149e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.263e-09 0 1.266e-09 0.0007 1.269e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.383e-09 0 1.386e-09 0.0007 1.389e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.503e-09 0 1.506e-09 0.0007 1.509e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.623e-09 0 1.626e-09 0.0007 1.629e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.743e-09 0 1.746e-09 0.0007 1.749e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.863e-09 0 1.866e-09 0.0007 1.869e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 1.983e-09 0 1.986e-09 0.0007 1.989e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.103e-09 0 2.106e-09 0.0007 2.109e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.223e-09 0 2.226e-09 0.0007 2.229e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.343e-09 0 2.346e-09 0.0007 2.349e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.463e-09 0 2.466e-09 0.0007 2.469e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.583e-09 0 2.586e-09 0.0007 2.589e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.703e-09 0 2.706e-09 0.0007 2.709e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.823e-09 0 2.826e-09 0.0007 2.829e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 2.943e-09 0 2.946e-09 0.0007 2.949e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.183e-09 0 3.186e-09 0.0007 3.189e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.303e-09 0 3.306e-09 0.0007 3.309e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.423e-09 0 3.426e-09 0.0007 3.429e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.543e-09 0 3.546e-09 0.0007 3.549e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.663e-09 0 3.666e-09 0.0007 3.669e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.783e-09 0 3.786e-09 0.0007 3.789e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.903e-09 0 3.906e-09 0.0007 3.909e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.023e-09 0 4.026e-09 0.0007 4.029e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.143e-09 0 4.146e-09 0.0007 4.149e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.383e-09 0 4.386e-09 0.0007 4.389e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.503e-09 0 4.506e-09 0.0007 4.509e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.623e-09 0 4.626e-09 0.0007 4.629e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.743e-09 0 4.746e-09 0.0007 4.749e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.863e-09 0 4.866e-09 0.0007 4.869e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 4.983e-09 0 4.986e-09 0.0007 4.989e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.103e-09 0 5.106e-09 0.0007 5.109e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.223e-09 0 5.226e-09 0.0007 5.229e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.343e-09 0 5.346e-09 0.0007 5.349e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.583e-09 0 5.586e-09 0.0007 5.589e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.703e-09 0 5.706e-09 0.0007 5.709e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.823e-09 0 5.826e-09 0.0007 5.829e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 5.943e-09 0 5.946e-09 0.0007 5.949e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.183e-09 0 6.186e-09 0.0007 6.189e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.303e-09 0 6.306e-09 0.0007 6.309e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.423e-09 0 6.426e-09 0.0007 6.429e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.543e-09 0 6.546e-09 0.0007 6.549e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.663e-09 0 6.666e-09 0.0007 6.669e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.783e-09 0 6.786e-09 0.0007 6.789e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.903e-09 0 6.906e-09 0.0007 6.909e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.023e-09 0 7.026e-09 0.0007 7.029e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.143e-09 0 7.146e-09 0.0007 7.149e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.263e-09 0 7.266e-09 0.0007 7.269e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.383e-09 0 7.386e-09 0.0007 7.389e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.503e-09 0 7.506e-09 0.0007 7.509e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.623e-09 0 7.626e-09 0.0007 7.629e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.743e-09 0 7.746e-09 0.0007 7.749e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 7.983e-09 0 7.986e-09 0.0007 7.989e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.103e-09 0 8.106e-09 0.0007 8.109e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.223e-09 0 8.226e-09 0.0007 8.229e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.343e-09 0 8.346e-09 0.0007 8.349e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.583e-09 0 8.586e-09 0.0007 8.589e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.703e-09 0 8.706e-09 0.0007 8.709e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.823e-09 0 8.826e-09 0.0007 8.829e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 8.943e-09 0 8.946e-09 0.0007 8.949e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.183e-09 0 9.186e-09 0.0007 9.189e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.303e-09 0 9.306e-09 0.0007 9.309e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.423e-09 0 9.426e-09 0.0007 9.429e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.543e-09 0 9.546e-09 0.0007 9.549e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.663e-09 0 9.666e-09 0.0007 9.669e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.783e-09 0 9.786e-09 0.0007 9.789e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.903e-09 0 9.906e-09 0.0007 9.909e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0007 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0007 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0007 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0007 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0007 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0007 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0007 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0007 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0007 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0007 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0007 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0007 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0007 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0007 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0007 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0007 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0007 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0007 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0007 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0007 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0007 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0007 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0007 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0007 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0007 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0007 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0007 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0007 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0007 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0007 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0007 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0007 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0007 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0007 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0007 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0007 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0007 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0007 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0007 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0007 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0007 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0007 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0007 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0007 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0007 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0007 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0007 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0007 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0007 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0007 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0007 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0007 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0007 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0007 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0007 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0007 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0007 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0007 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0007 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0007 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0007 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0007 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0007 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0007 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0007 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0007 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0007 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0007 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0007 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0007 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0007 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0007 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0007 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0007 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0007 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0007 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0007 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0007 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0007 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0007 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0007 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0007 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0007 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0007 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0007 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0007 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0007 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0007 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0007 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0007 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0007 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0007 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0007 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0007 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0)
L_DFF_IP1_12|1 IP1_1_OUT_RX _DFF_IP1_12|A1  2.067833848e-12
L_DFF_IP1_12|2 _DFF_IP1_12|A1 _DFF_IP1_12|A2  4.135667696e-12
L_DFF_IP1_12|3 _DFF_IP1_12|A3 _DFF_IP1_12|A4  8.271335392e-12
L_DFF_IP1_12|T D11 _DFF_IP1_12|T1  2.067833848e-12
L_DFF_IP1_12|4 _DFF_IP1_12|T1 _DFF_IP1_12|T2  4.135667696e-12
L_DFF_IP1_12|5 _DFF_IP1_12|A4 _DFF_IP1_12|Q1  4.135667696e-12
L_DFF_IP1_12|6 _DFF_IP1_12|Q1 IP1_2_OUT  2.067833848e-12
ID12|T 0 D12  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 6.3e-11 0 6.6e-11 0.0007 6.9e-11 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 1.83e-10 0 1.86e-10 0.0007 1.89e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.03e-10 0 3.06e-10 0.0007 3.09e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.23e-10 0 4.26e-10 0.0007 4.29e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 5.43e-10 0 5.46e-10 0.0007 5.49e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 6.63e-10 0 6.66e-10 0.0007 6.69e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 7.83e-10 0 7.86e-10 0.0007 7.89e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.03e-10 0 9.06e-10 0.0007 9.09e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.023e-09 0 1.026e-09 0.0007 1.029e-09 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.143e-09 0 1.146e-09 0.0007 1.149e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.263e-09 0 1.266e-09 0.0007 1.269e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.383e-09 0 1.386e-09 0.0007 1.389e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.503e-09 0 1.506e-09 0.0007 1.509e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.623e-09 0 1.626e-09 0.0007 1.629e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.743e-09 0 1.746e-09 0.0007 1.749e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.863e-09 0 1.866e-09 0.0007 1.869e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 1.983e-09 0 1.986e-09 0.0007 1.989e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.103e-09 0 2.106e-09 0.0007 2.109e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.223e-09 0 2.226e-09 0.0007 2.229e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.343e-09 0 2.346e-09 0.0007 2.349e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.463e-09 0 2.466e-09 0.0007 2.469e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.583e-09 0 2.586e-09 0.0007 2.589e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.703e-09 0 2.706e-09 0.0007 2.709e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.823e-09 0 2.826e-09 0.0007 2.829e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 2.943e-09 0 2.946e-09 0.0007 2.949e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.183e-09 0 3.186e-09 0.0007 3.189e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.303e-09 0 3.306e-09 0.0007 3.309e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.423e-09 0 3.426e-09 0.0007 3.429e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.543e-09 0 3.546e-09 0.0007 3.549e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.663e-09 0 3.666e-09 0.0007 3.669e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.783e-09 0 3.786e-09 0.0007 3.789e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.903e-09 0 3.906e-09 0.0007 3.909e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.023e-09 0 4.026e-09 0.0007 4.029e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.143e-09 0 4.146e-09 0.0007 4.149e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.383e-09 0 4.386e-09 0.0007 4.389e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.503e-09 0 4.506e-09 0.0007 4.509e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.623e-09 0 4.626e-09 0.0007 4.629e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.743e-09 0 4.746e-09 0.0007 4.749e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.863e-09 0 4.866e-09 0.0007 4.869e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 4.983e-09 0 4.986e-09 0.0007 4.989e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.103e-09 0 5.106e-09 0.0007 5.109e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.223e-09 0 5.226e-09 0.0007 5.229e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.343e-09 0 5.346e-09 0.0007 5.349e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.583e-09 0 5.586e-09 0.0007 5.589e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.703e-09 0 5.706e-09 0.0007 5.709e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.823e-09 0 5.826e-09 0.0007 5.829e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 5.943e-09 0 5.946e-09 0.0007 5.949e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.183e-09 0 6.186e-09 0.0007 6.189e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.303e-09 0 6.306e-09 0.0007 6.309e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.423e-09 0 6.426e-09 0.0007 6.429e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.543e-09 0 6.546e-09 0.0007 6.549e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.663e-09 0 6.666e-09 0.0007 6.669e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.783e-09 0 6.786e-09 0.0007 6.789e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.903e-09 0 6.906e-09 0.0007 6.909e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.023e-09 0 7.026e-09 0.0007 7.029e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.143e-09 0 7.146e-09 0.0007 7.149e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.263e-09 0 7.266e-09 0.0007 7.269e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.383e-09 0 7.386e-09 0.0007 7.389e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.503e-09 0 7.506e-09 0.0007 7.509e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.623e-09 0 7.626e-09 0.0007 7.629e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.743e-09 0 7.746e-09 0.0007 7.749e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 7.983e-09 0 7.986e-09 0.0007 7.989e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.103e-09 0 8.106e-09 0.0007 8.109e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.223e-09 0 8.226e-09 0.0007 8.229e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.343e-09 0 8.346e-09 0.0007 8.349e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.583e-09 0 8.586e-09 0.0007 8.589e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.703e-09 0 8.706e-09 0.0007 8.709e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.823e-09 0 8.826e-09 0.0007 8.829e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 8.943e-09 0 8.946e-09 0.0007 8.949e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.183e-09 0 9.186e-09 0.0007 9.189e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.303e-09 0 9.306e-09 0.0007 9.309e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.423e-09 0 9.426e-09 0.0007 9.429e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.543e-09 0 9.546e-09 0.0007 9.549e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.663e-09 0 9.666e-09 0.0007 9.669e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.783e-09 0 9.786e-09 0.0007 9.789e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.903e-09 0 9.906e-09 0.0007 9.909e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0007 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0007 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0007 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0007 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0007 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0007 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0007 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0007 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0007 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0007 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0007 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0007 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0007 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0007 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0007 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0007 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0007 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0007 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0007 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0007 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0007 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0007 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0007 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0007 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0007 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0007 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0007 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0007 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0007 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0007 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0007 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0007 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0007 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0007 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0007 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0007 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0007 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0007 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0007 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0007 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0007 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0007 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0007 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0007 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0007 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0007 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0007 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0007 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0007 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0007 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0007 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0007 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0007 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0007 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0007 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0007 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0007 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0007 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0007 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0007 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0007 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0007 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0007 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0007 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0007 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0007 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0007 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0007 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0007 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0007 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0007 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0007 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0007 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0007 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0007 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0007 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0007 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0007 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0007 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0007 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0007 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0007 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0007 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0007 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0007 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0007 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0007 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0007 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0007 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0007 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0007 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0007 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0007 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0007 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0)
L_DFF_IP2_12|1 IP2_1_OUT_RX _DFF_IP2_12|A1  2.067833848e-12
L_DFF_IP2_12|2 _DFF_IP2_12|A1 _DFF_IP2_12|A2  4.135667696e-12
L_DFF_IP2_12|3 _DFF_IP2_12|A3 _DFF_IP2_12|A4  8.271335392e-12
L_DFF_IP2_12|T D12 _DFF_IP2_12|T1  2.067833848e-12
L_DFF_IP2_12|4 _DFF_IP2_12|T1 _DFF_IP2_12|T2  4.135667696e-12
L_DFF_IP2_12|5 _DFF_IP2_12|A4 _DFF_IP2_12|Q1  4.135667696e-12
L_DFF_IP2_12|6 _DFF_IP2_12|Q1 IP2_2_OUT  2.067833848e-12
ID13|T 0 D13  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 6.3e-11 0 6.6e-11 0.0007 6.9e-11 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 1.83e-10 0 1.86e-10 0.0007 1.89e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.03e-10 0 3.06e-10 0.0007 3.09e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.23e-10 0 4.26e-10 0.0007 4.29e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 5.43e-10 0 5.46e-10 0.0007 5.49e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 6.63e-10 0 6.66e-10 0.0007 6.69e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 7.83e-10 0 7.86e-10 0.0007 7.89e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.03e-10 0 9.06e-10 0.0007 9.09e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.023e-09 0 1.026e-09 0.0007 1.029e-09 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.143e-09 0 1.146e-09 0.0007 1.149e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.263e-09 0 1.266e-09 0.0007 1.269e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.383e-09 0 1.386e-09 0.0007 1.389e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.503e-09 0 1.506e-09 0.0007 1.509e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.623e-09 0 1.626e-09 0.0007 1.629e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.743e-09 0 1.746e-09 0.0007 1.749e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.863e-09 0 1.866e-09 0.0007 1.869e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 1.983e-09 0 1.986e-09 0.0007 1.989e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.103e-09 0 2.106e-09 0.0007 2.109e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.223e-09 0 2.226e-09 0.0007 2.229e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.343e-09 0 2.346e-09 0.0007 2.349e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.463e-09 0 2.466e-09 0.0007 2.469e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.583e-09 0 2.586e-09 0.0007 2.589e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.703e-09 0 2.706e-09 0.0007 2.709e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.823e-09 0 2.826e-09 0.0007 2.829e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 2.943e-09 0 2.946e-09 0.0007 2.949e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.183e-09 0 3.186e-09 0.0007 3.189e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.303e-09 0 3.306e-09 0.0007 3.309e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.423e-09 0 3.426e-09 0.0007 3.429e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.543e-09 0 3.546e-09 0.0007 3.549e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.663e-09 0 3.666e-09 0.0007 3.669e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.783e-09 0 3.786e-09 0.0007 3.789e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.903e-09 0 3.906e-09 0.0007 3.909e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.023e-09 0 4.026e-09 0.0007 4.029e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.143e-09 0 4.146e-09 0.0007 4.149e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.383e-09 0 4.386e-09 0.0007 4.389e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.503e-09 0 4.506e-09 0.0007 4.509e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.623e-09 0 4.626e-09 0.0007 4.629e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.743e-09 0 4.746e-09 0.0007 4.749e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.863e-09 0 4.866e-09 0.0007 4.869e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 4.983e-09 0 4.986e-09 0.0007 4.989e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.103e-09 0 5.106e-09 0.0007 5.109e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.223e-09 0 5.226e-09 0.0007 5.229e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.343e-09 0 5.346e-09 0.0007 5.349e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.583e-09 0 5.586e-09 0.0007 5.589e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.703e-09 0 5.706e-09 0.0007 5.709e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.823e-09 0 5.826e-09 0.0007 5.829e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 5.943e-09 0 5.946e-09 0.0007 5.949e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.183e-09 0 6.186e-09 0.0007 6.189e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.303e-09 0 6.306e-09 0.0007 6.309e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.423e-09 0 6.426e-09 0.0007 6.429e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.543e-09 0 6.546e-09 0.0007 6.549e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.663e-09 0 6.666e-09 0.0007 6.669e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.783e-09 0 6.786e-09 0.0007 6.789e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.903e-09 0 6.906e-09 0.0007 6.909e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.023e-09 0 7.026e-09 0.0007 7.029e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.143e-09 0 7.146e-09 0.0007 7.149e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.263e-09 0 7.266e-09 0.0007 7.269e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.383e-09 0 7.386e-09 0.0007 7.389e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.503e-09 0 7.506e-09 0.0007 7.509e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.623e-09 0 7.626e-09 0.0007 7.629e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.743e-09 0 7.746e-09 0.0007 7.749e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 7.983e-09 0 7.986e-09 0.0007 7.989e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.103e-09 0 8.106e-09 0.0007 8.109e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.223e-09 0 8.226e-09 0.0007 8.229e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.343e-09 0 8.346e-09 0.0007 8.349e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.583e-09 0 8.586e-09 0.0007 8.589e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.703e-09 0 8.706e-09 0.0007 8.709e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.823e-09 0 8.826e-09 0.0007 8.829e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 8.943e-09 0 8.946e-09 0.0007 8.949e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.183e-09 0 9.186e-09 0.0007 9.189e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.303e-09 0 9.306e-09 0.0007 9.309e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.423e-09 0 9.426e-09 0.0007 9.429e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.543e-09 0 9.546e-09 0.0007 9.549e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.663e-09 0 9.666e-09 0.0007 9.669e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.783e-09 0 9.786e-09 0.0007 9.789e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.903e-09 0 9.906e-09 0.0007 9.909e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0023e-08 0 1.0026e-08 0.0007 1.0029e-08 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0143e-08 0 1.0146e-08 0.0007 1.0149e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0383e-08 0 1.0386e-08 0.0007 1.0389e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0503e-08 0 1.0506e-08 0.0007 1.0509e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0623e-08 0 1.0626e-08 0.0007 1.0629e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0743e-08 0 1.0746e-08 0.0007 1.0749e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.0983e-08 0 1.0986e-08 0.0007 1.0989e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1103e-08 0 1.1106e-08 0.0007 1.1109e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1223e-08 0 1.1226e-08 0.0007 1.1229e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1343e-08 0 1.1346e-08 0.0007 1.1349e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1583e-08 0 1.1586e-08 0.0007 1.1589e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1703e-08 0 1.1706e-08 0.0007 1.1709e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1823e-08 0 1.1826e-08 0.0007 1.1829e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.1943e-08 0 1.1946e-08 0.0007 1.1949e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2183e-08 0 1.2186e-08 0.0007 1.2189e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2303e-08 0 1.2306e-08 0.0007 1.2309e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2423e-08 0 1.2426e-08 0.0007 1.2429e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2543e-08 0 1.2546e-08 0.0007 1.2549e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2783e-08 0 1.2786e-08 0.0007 1.2789e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2903e-08 0 1.2906e-08 0.0007 1.2909e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3023e-08 0 1.3026e-08 0.0007 1.3029e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3143e-08 0 1.3146e-08 0.0007 1.3149e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3263e-08 0 1.3266e-08 0.0007 1.3269e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3383e-08 0 1.3386e-08 0.0007 1.3389e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3503e-08 0 1.3506e-08 0.0007 1.3509e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3623e-08 0 1.3626e-08 0.0007 1.3629e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3743e-08 0 1.3746e-08 0.0007 1.3749e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.3983e-08 0 1.3986e-08 0.0007 1.3989e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4103e-08 0 1.4106e-08 0.0007 1.4109e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4223e-08 0 1.4226e-08 0.0007 1.4229e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4343e-08 0 1.4346e-08 0.0007 1.4349e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4463e-08 0 1.4466e-08 0.0007 1.4469e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4583e-08 0 1.4586e-08 0.0007 1.4589e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4703e-08 0 1.4706e-08 0.0007 1.4709e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.4943e-08 0 1.4946e-08 0.0007 1.4949e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5183e-08 0 1.5186e-08 0.0007 1.5189e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5303e-08 0 1.5306e-08 0.0007 1.5309e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5423e-08 0 1.5426e-08 0.0007 1.5429e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5543e-08 0 1.5546e-08 0.0007 1.5549e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5783e-08 0 1.5786e-08 0.0007 1.5789e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5903e-08 0 1.5906e-08 0.0007 1.5909e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6023e-08 0 1.6026e-08 0.0007 1.6029e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6143e-08 0 1.6146e-08 0.0007 1.6149e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6383e-08 0 1.6386e-08 0.0007 1.6389e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6503e-08 0 1.6506e-08 0.0007 1.6509e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6623e-08 0 1.6626e-08 0.0007 1.6629e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6743e-08 0 1.6746e-08 0.0007 1.6749e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.6983e-08 0 1.6986e-08 0.0007 1.6989e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7103e-08 0 1.7106e-08 0.0007 1.7109e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7223e-08 0 1.7226e-08 0.0007 1.7229e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7343e-08 0 1.7346e-08 0.0007 1.7349e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7583e-08 0 1.7586e-08 0.0007 1.7589e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7703e-08 0 1.7706e-08 0.0007 1.7709e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7823e-08 0 1.7826e-08 0.0007 1.7829e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.7943e-08 0 1.7946e-08 0.0007 1.7949e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8183e-08 0 1.8186e-08 0.0007 1.8189e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8303e-08 0 1.8306e-08 0.0007 1.8309e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8423e-08 0 1.8426e-08 0.0007 1.8429e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8543e-08 0 1.8546e-08 0.0007 1.8549e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8783e-08 0 1.8786e-08 0.0007 1.8789e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8903e-08 0 1.8906e-08 0.0007 1.8909e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9023e-08 0 1.9026e-08 0.0007 1.9029e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9143e-08 0 1.9146e-08 0.0007 1.9149e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9263e-08 0 1.9266e-08 0.0007 1.9269e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9383e-08 0 1.9386e-08 0.0007 1.9389e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9503e-08 0 1.9506e-08 0.0007 1.9509e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9623e-08 0 1.9626e-08 0.0007 1.9629e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9743e-08 0 1.9746e-08 0.0007 1.9749e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 1.9983e-08 0 1.9986e-08 0.0007 1.9989e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0103e-08 0 2.0106e-08 0.0007 2.0109e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0223e-08 0 2.0226e-08 0.0007 2.0229e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0343e-08 0 2.0346e-08 0.0007 2.0349e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0583e-08 0 2.0586e-08 0.0007 2.0589e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0703e-08 0 2.0706e-08 0.0007 2.0709e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0823e-08 0 2.0826e-08 0.0007 2.0829e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.0943e-08 0 2.0946e-08 0.0007 2.0949e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1183e-08 0 2.1186e-08 0.0007 2.1189e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1303e-08 0 2.1306e-08 0.0007 2.1309e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1423e-08 0 2.1426e-08 0.0007 2.1429e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1543e-08 0 2.1546e-08 0.0007 2.1549e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1783e-08 0 2.1786e-08 0.0007 2.1789e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1903e-08 0 2.1906e-08 0.0007 2.1909e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2023e-08 0 2.2026e-08 0.0007 2.2029e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2383e-08 0 2.2386e-08 0.0007 2.2389e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2503e-08 0 2.2506e-08 0.0007 2.2509e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2623e-08 0 2.2626e-08 0.0007 2.2629e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2743e-08 0 2.2746e-08 0.0007 2.2749e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.2983e-08 0 2.2986e-08 0.0007 2.2989e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3103e-08 0 2.3106e-08 0.0007 2.3109e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3223e-08 0 2.3226e-08 0.0007 2.3229e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3343e-08 0 2.3346e-08 0.0007 2.3349e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3583e-08 0 2.3586e-08 0.0007 2.3589e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3703e-08 0 2.3706e-08 0.0007 2.3709e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3823e-08 0 2.3826e-08 0.0007 2.3829e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0)
L_DFF_IP3_12|1 IP3_1_OUT_RX _DFF_IP3_12|A1  2.067833848e-12
L_DFF_IP3_12|2 _DFF_IP3_12|A1 _DFF_IP3_12|A2  4.135667696e-12
L_DFF_IP3_12|3 _DFF_IP3_12|A3 _DFF_IP3_12|A4  8.271335392e-12
L_DFF_IP3_12|T D13 _DFF_IP3_12|T1  2.067833848e-12
L_DFF_IP3_12|4 _DFF_IP3_12|T1 _DFF_IP3_12|T2  4.135667696e-12
L_DFF_IP3_12|5 _DFF_IP3_12|A4 _DFF_IP3_12|Q1  4.135667696e-12
L_DFF_IP3_12|6 _DFF_IP3_12|Q1 IP3_2_OUT  2.067833848e-12
IT12|T 0 T12  PWL(0 0 0 0 3e-12 0.0007 6e-12 0 6e-11 0 6.3e-11 0.0007 6.6e-11 0 1.2e-10 0 1.23e-10 0.0007 1.26e-10 0 1.8e-10 0 1.83e-10 0.0007 1.86e-10 0 2.4e-10 0 2.43e-10 0.0007 2.46e-10 0 3e-10 0 3.03e-10 0.0007 3.06e-10 0 3.6e-10 0 3.63e-10 0.0007 3.66e-10 0 4.2e-10 0 4.23e-10 0.0007 4.26e-10 0 4.8e-10 0 4.83e-10 0.0007 4.86e-10 0 5.4e-10 0 5.43e-10 0.0007 5.46e-10 0 6e-10 0 6.03e-10 0.0007 6.06e-10 0 6.6e-10 0 6.63e-10 0.0007 6.66e-10 0 7.2e-10 0 7.23e-10 0.0007 7.26e-10 0 7.8e-10 0 7.83e-10 0.0007 7.86e-10 0 8.4e-10 0 8.43e-10 0.0007 8.46e-10 0 9e-10 0 9.03e-10 0.0007 9.06e-10 0 9.6e-10 0 9.63e-10 0.0007 9.66e-10 0 1.02e-09 0 1.023e-09 0.0007 1.026e-09 0 1.08e-09 0 1.083e-09 0.0007 1.086e-09 0 1.14e-09 0 1.143e-09 0.0007 1.146e-09 0 1.2e-09 0 1.203e-09 0.0007 1.206e-09 0 1.26e-09 0 1.263e-09 0.0007 1.266e-09 0 1.32e-09 0 1.323e-09 0.0007 1.326e-09 0 1.38e-09 0 1.383e-09 0.0007 1.386e-09 0 1.44e-09 0 1.443e-09 0.0007 1.446e-09 0 1.5e-09 0 1.503e-09 0.0007 1.506e-09 0 1.56e-09 0 1.563e-09 0.0007 1.566e-09 0 1.62e-09 0 1.623e-09 0.0007 1.626e-09 0 1.68e-09 0 1.683e-09 0.0007 1.686e-09 0 1.74e-09 0 1.743e-09 0.0007 1.746e-09 0 1.8e-09 0 1.803e-09 0.0007 1.806e-09 0 1.86e-09 0 1.863e-09 0.0007 1.866e-09 0 1.92e-09 0 1.923e-09 0.0007 1.926e-09 0 1.98e-09 0 1.983e-09 0.0007 1.986e-09 0 2.04e-09 0 2.043e-09 0.0007 2.046e-09 0 2.1e-09 0 2.103e-09 0.0007 2.106e-09 0 2.16e-09 0 2.163e-09 0.0007 2.166e-09 0 2.22e-09 0 2.223e-09 0.0007 2.226e-09 0 2.28e-09 0 2.283e-09 0.0007 2.286e-09 0 2.34e-09 0 2.343e-09 0.0007 2.346e-09 0 2.4e-09 0 2.403e-09 0.0007 2.406e-09 0 2.46e-09 0 2.463e-09 0.0007 2.466e-09 0 2.52e-09 0 2.523e-09 0.0007 2.526e-09 0 2.58e-09 0 2.583e-09 0.0007 2.586e-09 0 2.64e-09 0 2.643e-09 0.0007 2.646e-09 0 2.7e-09 0 2.703e-09 0.0007 2.706e-09 0 2.76e-09 0 2.763e-09 0.0007 2.766e-09 0 2.82e-09 0 2.823e-09 0.0007 2.826e-09 0 2.88e-09 0 2.883e-09 0.0007 2.886e-09 0 2.94e-09 0 2.943e-09 0.0007 2.946e-09 0 3e-09 0 3.003e-09 0.0007 3.006e-09 0 3.06e-09 0 3.063e-09 0.0007 3.066e-09 0 3.12e-09 0 3.123e-09 0.0007 3.126e-09 0 3.18e-09 0 3.183e-09 0.0007 3.186e-09 0 3.24e-09 0 3.243e-09 0.0007 3.246e-09 0 3.3e-09 0 3.303e-09 0.0007 3.306e-09 0 3.36e-09 0 3.363e-09 0.0007 3.366e-09 0 3.42e-09 0 3.423e-09 0.0007 3.426e-09 0 3.48e-09 0 3.483e-09 0.0007 3.486e-09 0 3.54e-09 0 3.543e-09 0.0007 3.546e-09 0 3.6e-09 0 3.603e-09 0.0007 3.606e-09 0 3.66e-09 0 3.663e-09 0.0007 3.666e-09 0 3.72e-09 0 3.723e-09 0.0007 3.726e-09 0 3.78e-09 0 3.783e-09 0.0007 3.786e-09 0 3.84e-09 0 3.843e-09 0.0007 3.846e-09 0 3.9e-09 0 3.903e-09 0.0007 3.906e-09 0 3.96e-09 0 3.963e-09 0.0007 3.966e-09 0 4.02e-09 0 4.023e-09 0.0007 4.026e-09 0 4.08e-09 0 4.083e-09 0.0007 4.086e-09 0 4.14e-09 0 4.143e-09 0.0007 4.146e-09 0 4.2e-09 0 4.203e-09 0.0007 4.206e-09 0 4.26e-09 0 4.263e-09 0.0007 4.266e-09 0 4.32e-09 0 4.323e-09 0.0007 4.326e-09 0 4.38e-09 0 4.383e-09 0.0007 4.386e-09 0 4.44e-09 0 4.443e-09 0.0007 4.446e-09 0 4.5e-09 0 4.503e-09 0.0007 4.506e-09 0 4.56e-09 0 4.563e-09 0.0007 4.566e-09 0 4.62e-09 0 4.623e-09 0.0007 4.626e-09 0 4.68e-09 0 4.683e-09 0.0007 4.686e-09 0 4.74e-09 0 4.743e-09 0.0007 4.746e-09 0 4.8e-09 0 4.803e-09 0.0007 4.806e-09 0 4.86e-09 0 4.863e-09 0.0007 4.866e-09 0 4.92e-09 0 4.923e-09 0.0007 4.926e-09 0 4.98e-09 0 4.983e-09 0.0007 4.986e-09 0 5.04e-09 0 5.043e-09 0.0007 5.046e-09 0 5.1e-09 0 5.103e-09 0.0007 5.106e-09 0 5.16e-09 0 5.163e-09 0.0007 5.166e-09 0 5.22e-09 0 5.223e-09 0.0007 5.226e-09 0 5.28e-09 0 5.283e-09 0.0007 5.286e-09 0 5.34e-09 0 5.343e-09 0.0007 5.346e-09 0 5.4e-09 0 5.403e-09 0.0007 5.406e-09 0 5.46e-09 0 5.463e-09 0.0007 5.466e-09 0 5.52e-09 0 5.523e-09 0.0007 5.526e-09 0 5.58e-09 0 5.583e-09 0.0007 5.586e-09 0 5.64e-09 0 5.643e-09 0.0007 5.646e-09 0 5.7e-09 0 5.703e-09 0.0007 5.706e-09 0 5.76e-09 0 5.763e-09 0.0007 5.766e-09 0 5.82e-09 0 5.823e-09 0.0007 5.826e-09 0 5.88e-09 0 5.883e-09 0.0007 5.886e-09 0 5.94e-09 0 5.943e-09 0.0007 5.946e-09 0 6e-09 0 6.003e-09 0.0007 6.006e-09 0 6.06e-09 0 6.063e-09 0.0007 6.066e-09 0 6.12e-09 0 6.123e-09 0.0007 6.126e-09 0 6.18e-09 0 6.183e-09 0.0007 6.186e-09 0 6.24e-09 0 6.243e-09 0.0007 6.246e-09 0 6.3e-09 0 6.303e-09 0.0007 6.306e-09 0 6.36e-09 0 6.363e-09 0.0007 6.366e-09 0 6.42e-09 0 6.423e-09 0.0007 6.426e-09 0 6.48e-09 0 6.483e-09 0.0007 6.486e-09 0 6.54e-09 0 6.543e-09 0.0007 6.546e-09 0 6.6e-09 0 6.603e-09 0.0007 6.606e-09 0 6.66e-09 0 6.663e-09 0.0007 6.666e-09 0 6.72e-09 0 6.723e-09 0.0007 6.726e-09 0 6.78e-09 0 6.783e-09 0.0007 6.786e-09 0 6.84e-09 0 6.843e-09 0.0007 6.846e-09 0 6.9e-09 0 6.903e-09 0.0007 6.906e-09 0 6.96e-09 0 6.963e-09 0.0007 6.966e-09 0 7.02e-09 0 7.023e-09 0.0007 7.026e-09 0 7.08e-09 0 7.083e-09 0.0007 7.086e-09 0 7.14e-09 0 7.143e-09 0.0007 7.146e-09 0 7.2e-09 0 7.203e-09 0.0007 7.206e-09 0 7.26e-09 0 7.263e-09 0.0007 7.266e-09 0 7.32e-09 0 7.323e-09 0.0007 7.326e-09 0 7.38e-09 0 7.383e-09 0.0007 7.386e-09 0 7.44e-09 0 7.443e-09 0.0007 7.446e-09 0 7.5e-09 0 7.503e-09 0.0007 7.506e-09 0 7.56e-09 0 7.563e-09 0.0007 7.566e-09 0 7.62e-09 0 7.623e-09 0.0007 7.626e-09 0 7.68e-09 0 7.683e-09 0.0007 7.686e-09 0 7.74e-09 0 7.743e-09 0.0007 7.746e-09 0 7.8e-09 0 7.803e-09 0.0007 7.806e-09 0 7.86e-09 0 7.863e-09 0.0007 7.866e-09 0 7.92e-09 0 7.923e-09 0.0007 7.926e-09 0 7.98e-09 0 7.983e-09 0.0007 7.986e-09 0 8.04e-09 0 8.043e-09 0.0007 8.046e-09 0 8.1e-09 0 8.103e-09 0.0007 8.106e-09 0 8.16e-09 0 8.163e-09 0.0007 8.166e-09 0 8.22e-09 0 8.223e-09 0.0007 8.226e-09 0 8.28e-09 0 8.283e-09 0.0007 8.286e-09 0 8.34e-09 0 8.343e-09 0.0007 8.346e-09 0 8.4e-09 0 8.403e-09 0.0007 8.406e-09 0 8.46e-09 0 8.463e-09 0.0007 8.466e-09 0 8.52e-09 0 8.523e-09 0.0007 8.526e-09 0 8.58e-09 0 8.583e-09 0.0007 8.586e-09 0 8.64e-09 0 8.643e-09 0.0007 8.646e-09 0 8.7e-09 0 8.703e-09 0.0007 8.706e-09 0 8.76e-09 0 8.763e-09 0.0007 8.766e-09 0 8.82e-09 0 8.823e-09 0.0007 8.826e-09 0 8.88e-09 0 8.883e-09 0.0007 8.886e-09 0 8.94e-09 0 8.943e-09 0.0007 8.946e-09 0 9e-09 0 9.003e-09 0.0007 9.006e-09 0 9.06e-09 0 9.063e-09 0.0007 9.066e-09 0 9.12e-09 0 9.123e-09 0.0007 9.126e-09 0 9.18e-09 0 9.183e-09 0.0007 9.186e-09 0 9.24e-09 0 9.243e-09 0.0007 9.246e-09 0 9.3e-09 0 9.303e-09 0.0007 9.306e-09 0 9.36e-09 0 9.363e-09 0.0007 9.366e-09 0 9.42e-09 0 9.423e-09 0.0007 9.426e-09 0 9.48e-09 0 9.483e-09 0.0007 9.486e-09 0 9.54e-09 0 9.543e-09 0.0007 9.546e-09 0 9.6e-09 0 9.603e-09 0.0007 9.606e-09 0 9.66e-09 0 9.663e-09 0.0007 9.666e-09 0 9.72e-09 0 9.723e-09 0.0007 9.726e-09 0 9.78e-09 0 9.783e-09 0.0007 9.786e-09 0 9.84e-09 0 9.843e-09 0.0007 9.846e-09 0 9.9e-09 0 9.903e-09 0.0007 9.906e-09 0 9.96e-09 0 9.963e-09 0.0007 9.966e-09 0 1.002e-08 0 1.0023e-08 0.0007 1.0026e-08 0 1.008e-08 0 1.0083e-08 0.0007 1.0086e-08 0 1.014e-08 0 1.0143e-08 0.0007 1.0146e-08 0 1.02e-08 0 1.0203e-08 0.0007 1.0206e-08 0 1.026e-08 0 1.0263e-08 0.0007 1.0266e-08 0 1.032e-08 0 1.0323e-08 0.0007 1.0326e-08 0 1.038e-08 0 1.0383e-08 0.0007 1.0386e-08 0 1.044e-08 0 1.0443e-08 0.0007 1.0446e-08 0 1.05e-08 0 1.0503e-08 0.0007 1.0506e-08 0 1.056e-08 0 1.0563e-08 0.0007 1.0566e-08 0 1.062e-08 0 1.0623e-08 0.0007 1.0626e-08 0 1.068e-08 0 1.0683e-08 0.0007 1.0686e-08 0 1.074e-08 0 1.0743e-08 0.0007 1.0746e-08 0 1.08e-08 0 1.0803e-08 0.0007 1.0806e-08 0 1.086e-08 0 1.0863e-08 0.0007 1.0866e-08 0 1.092e-08 0 1.0923e-08 0.0007 1.0926e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.104e-08 0 1.1043e-08 0.0007 1.1046e-08 0 1.11e-08 0 1.1103e-08 0.0007 1.1106e-08 0 1.116e-08 0 1.1163e-08 0.0007 1.1166e-08 0 1.122e-08 0 1.1223e-08 0.0007 1.1226e-08 0 1.128e-08 0 1.1283e-08 0.0007 1.1286e-08 0 1.134e-08 0 1.1343e-08 0.0007 1.1346e-08 0 1.14e-08 0 1.1403e-08 0.0007 1.1406e-08 0 1.146e-08 0 1.1463e-08 0.0007 1.1466e-08 0 1.152e-08 0 1.1523e-08 0.0007 1.1526e-08 0 1.158e-08 0 1.1583e-08 0.0007 1.1586e-08 0 1.164e-08 0 1.1643e-08 0.0007 1.1646e-08 0 1.17e-08 0 1.1703e-08 0.0007 1.1706e-08 0 1.176e-08 0 1.1763e-08 0.0007 1.1766e-08 0 1.182e-08 0 1.1823e-08 0.0007 1.1826e-08 0 1.188e-08 0 1.1883e-08 0.0007 1.1886e-08 0 1.194e-08 0 1.1943e-08 0.0007 1.1946e-08 0 1.2e-08 0 1.2003e-08 0.0007 1.2006e-08 0 1.206e-08 0 1.2063e-08 0.0007 1.2066e-08 0 1.212e-08 0 1.2123e-08 0.0007 1.2126e-08 0 1.218e-08 0 1.2183e-08 0.0007 1.2186e-08 0 1.224e-08 0 1.2243e-08 0.0007 1.2246e-08 0 1.23e-08 0 1.2303e-08 0.0007 1.2306e-08 0 1.236e-08 0 1.2363e-08 0.0007 1.2366e-08 0 1.242e-08 0 1.2423e-08 0.0007 1.2426e-08 0 1.248e-08 0 1.2483e-08 0.0007 1.2486e-08 0 1.254e-08 0 1.2543e-08 0.0007 1.2546e-08 0 1.26e-08 0 1.2603e-08 0.0007 1.2606e-08 0 1.266e-08 0 1.2663e-08 0.0007 1.2666e-08 0 1.272e-08 0 1.2723e-08 0.0007 1.2726e-08 0 1.278e-08 0 1.2783e-08 0.0007 1.2786e-08 0 1.284e-08 0 1.2843e-08 0.0007 1.2846e-08 0 1.29e-08 0 1.2903e-08 0.0007 1.2906e-08 0 1.296e-08 0 1.2963e-08 0.0007 1.2966e-08 0 1.302e-08 0 1.3023e-08 0.0007 1.3026e-08 0 1.308e-08 0 1.3083e-08 0.0007 1.3086e-08 0 1.314e-08 0 1.3143e-08 0.0007 1.3146e-08 0 1.32e-08 0 1.3203e-08 0.0007 1.3206e-08 0 1.326e-08 0 1.3263e-08 0.0007 1.3266e-08 0 1.332e-08 0 1.3323e-08 0.0007 1.3326e-08 0 1.338e-08 0 1.3383e-08 0.0007 1.3386e-08 0 1.344e-08 0 1.3443e-08 0.0007 1.3446e-08 0 1.35e-08 0 1.3503e-08 0.0007 1.3506e-08 0 1.356e-08 0 1.3563e-08 0.0007 1.3566e-08 0 1.362e-08 0 1.3623e-08 0.0007 1.3626e-08 0 1.368e-08 0 1.3683e-08 0.0007 1.3686e-08 0 1.374e-08 0 1.3743e-08 0.0007 1.3746e-08 0 1.38e-08 0 1.3803e-08 0.0007 1.3806e-08 0 1.386e-08 0 1.3863e-08 0.0007 1.3866e-08 0 1.392e-08 0 1.3923e-08 0.0007 1.3926e-08 0 1.398e-08 0 1.3983e-08 0.0007 1.3986e-08 0 1.404e-08 0 1.4043e-08 0.0007 1.4046e-08 0 1.41e-08 0 1.4103e-08 0.0007 1.4106e-08 0 1.416e-08 0 1.4163e-08 0.0007 1.4166e-08 0 1.422e-08 0 1.4223e-08 0.0007 1.4226e-08 0 1.428e-08 0 1.4283e-08 0.0007 1.4286e-08 0 1.434e-08 0 1.4343e-08 0.0007 1.4346e-08 0 1.44e-08 0 1.4403e-08 0.0007 1.4406e-08 0 1.446e-08 0 1.4463e-08 0.0007 1.4466e-08 0 1.452e-08 0 1.4523e-08 0.0007 1.4526e-08 0 1.458e-08 0 1.4583e-08 0.0007 1.4586e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.47e-08 0 1.4703e-08 0.0007 1.4706e-08 0 1.476e-08 0 1.4763e-08 0.0007 1.4766e-08 0 1.482e-08 0 1.4823e-08 0.0007 1.4826e-08 0 1.488e-08 0 1.4883e-08 0.0007 1.4886e-08 0 1.494e-08 0 1.4943e-08 0.0007 1.4946e-08 0 1.5e-08 0 1.5003e-08 0.0007 1.5006e-08 0 1.506e-08 0 1.5063e-08 0.0007 1.5066e-08 0 1.512e-08 0 1.5123e-08 0.0007 1.5126e-08 0 1.518e-08 0 1.5183e-08 0.0007 1.5186e-08 0 1.524e-08 0 1.5243e-08 0.0007 1.5246e-08 0 1.53e-08 0 1.5303e-08 0.0007 1.5306e-08 0 1.536e-08 0 1.5363e-08 0.0007 1.5366e-08 0 1.542e-08 0 1.5423e-08 0.0007 1.5426e-08 0 1.548e-08 0 1.5483e-08 0.0007 1.5486e-08 0 1.554e-08 0 1.5543e-08 0.0007 1.5546e-08 0 1.56e-08 0 1.5603e-08 0.0007 1.5606e-08 0 1.566e-08 0 1.5663e-08 0.0007 1.5666e-08 0 1.572e-08 0 1.5723e-08 0.0007 1.5726e-08 0 1.578e-08 0 1.5783e-08 0.0007 1.5786e-08 0 1.584e-08 0 1.5843e-08 0.0007 1.5846e-08 0 1.59e-08 0 1.5903e-08 0.0007 1.5906e-08 0 1.596e-08 0 1.5963e-08 0.0007 1.5966e-08 0 1.602e-08 0 1.6023e-08 0.0007 1.6026e-08 0 1.608e-08 0 1.6083e-08 0.0007 1.6086e-08 0 1.614e-08 0 1.6143e-08 0.0007 1.6146e-08 0 1.62e-08 0 1.6203e-08 0.0007 1.6206e-08 0 1.626e-08 0 1.6263e-08 0.0007 1.6266e-08 0 1.632e-08 0 1.6323e-08 0.0007 1.6326e-08 0 1.638e-08 0 1.6383e-08 0.0007 1.6386e-08 0 1.644e-08 0 1.6443e-08 0.0007 1.6446e-08 0 1.65e-08 0 1.6503e-08 0.0007 1.6506e-08 0 1.656e-08 0 1.6563e-08 0.0007 1.6566e-08 0 1.662e-08 0 1.6623e-08 0.0007 1.6626e-08 0 1.668e-08 0 1.6683e-08 0.0007 1.6686e-08 0 1.674e-08 0 1.6743e-08 0.0007 1.6746e-08 0 1.68e-08 0 1.6803e-08 0.0007 1.6806e-08 0 1.686e-08 0 1.6863e-08 0.0007 1.6866e-08 0 1.692e-08 0 1.6923e-08 0.0007 1.6926e-08 0 1.698e-08 0 1.6983e-08 0.0007 1.6986e-08 0 1.704e-08 0 1.7043e-08 0.0007 1.7046e-08 0 1.71e-08 0 1.7103e-08 0.0007 1.7106e-08 0 1.716e-08 0 1.7163e-08 0.0007 1.7166e-08 0 1.722e-08 0 1.7223e-08 0.0007 1.7226e-08 0 1.728e-08 0 1.7283e-08 0.0007 1.7286e-08 0 1.734e-08 0 1.7343e-08 0.0007 1.7346e-08 0 1.74e-08 0 1.7403e-08 0.0007 1.7406e-08 0 1.746e-08 0 1.7463e-08 0.0007 1.7466e-08 0 1.752e-08 0 1.7523e-08 0.0007 1.7526e-08 0 1.758e-08 0 1.7583e-08 0.0007 1.7586e-08 0 1.764e-08 0 1.7643e-08 0.0007 1.7646e-08 0 1.77e-08 0 1.7703e-08 0.0007 1.7706e-08 0 1.776e-08 0 1.7763e-08 0.0007 1.7766e-08 0 1.782e-08 0 1.7823e-08 0.0007 1.7826e-08 0 1.788e-08 0 1.7883e-08 0.0007 1.7886e-08 0 1.794e-08 0 1.7943e-08 0.0007 1.7946e-08 0 1.8e-08 0 1.8003e-08 0.0007 1.8006e-08 0 1.806e-08 0 1.8063e-08 0.0007 1.8066e-08 0 1.812e-08 0 1.8123e-08 0.0007 1.8126e-08 0 1.818e-08 0 1.8183e-08 0.0007 1.8186e-08 0 1.824e-08 0 1.8243e-08 0.0007 1.8246e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.836e-08 0 1.8363e-08 0.0007 1.8366e-08 0 1.842e-08 0 1.8423e-08 0.0007 1.8426e-08 0 1.848e-08 0 1.8483e-08 0.0007 1.8486e-08 0 1.854e-08 0 1.8543e-08 0.0007 1.8546e-08 0 1.86e-08 0 1.8603e-08 0.0007 1.8606e-08 0 1.866e-08 0 1.8663e-08 0.0007 1.8666e-08 0 1.872e-08 0 1.8723e-08 0.0007 1.8726e-08 0 1.878e-08 0 1.8783e-08 0.0007 1.8786e-08 0 1.884e-08 0 1.8843e-08 0.0007 1.8846e-08 0 1.89e-08 0 1.8903e-08 0.0007 1.8906e-08 0 1.896e-08 0 1.8963e-08 0.0007 1.8966e-08 0 1.902e-08 0 1.9023e-08 0.0007 1.9026e-08 0 1.908e-08 0 1.9083e-08 0.0007 1.9086e-08 0 1.914e-08 0 1.9143e-08 0.0007 1.9146e-08 0 1.92e-08 0 1.9203e-08 0.0007 1.9206e-08 0 1.926e-08 0 1.9263e-08 0.0007 1.9266e-08 0 1.932e-08 0 1.9323e-08 0.0007 1.9326e-08 0 1.938e-08 0 1.9383e-08 0.0007 1.9386e-08 0 1.944e-08 0 1.9443e-08 0.0007 1.9446e-08 0 1.95e-08 0 1.9503e-08 0.0007 1.9506e-08 0 1.956e-08 0 1.9563e-08 0.0007 1.9566e-08 0 1.962e-08 0 1.9623e-08 0.0007 1.9626e-08 0 1.968e-08 0 1.9683e-08 0.0007 1.9686e-08 0 1.974e-08 0 1.9743e-08 0.0007 1.9746e-08 0 1.98e-08 0 1.9803e-08 0.0007 1.9806e-08 0 1.986e-08 0 1.9863e-08 0.0007 1.9866e-08 0 1.992e-08 0 1.9923e-08 0.0007 1.9926e-08 0 1.998e-08 0 1.9983e-08 0.0007 1.9986e-08 0 2.004e-08 0 2.0043e-08 0.0007 2.0046e-08 0 2.01e-08 0 2.0103e-08 0.0007 2.0106e-08 0 2.016e-08 0 2.0163e-08 0.0007 2.0166e-08 0 2.022e-08 0 2.0223e-08 0.0007 2.0226e-08 0 2.028e-08 0 2.0283e-08 0.0007 2.0286e-08 0 2.034e-08 0 2.0343e-08 0.0007 2.0346e-08 0 2.04e-08 0 2.0403e-08 0.0007 2.0406e-08 0 2.046e-08 0 2.0463e-08 0.0007 2.0466e-08 0 2.052e-08 0 2.0523e-08 0.0007 2.0526e-08 0 2.058e-08 0 2.0583e-08 0.0007 2.0586e-08 0 2.064e-08 0 2.0643e-08 0.0007 2.0646e-08 0 2.07e-08 0 2.0703e-08 0.0007 2.0706e-08 0 2.076e-08 0 2.0763e-08 0.0007 2.0766e-08 0 2.082e-08 0 2.0823e-08 0.0007 2.0826e-08 0 2.088e-08 0 2.0883e-08 0.0007 2.0886e-08 0 2.094e-08 0 2.0943e-08 0.0007 2.0946e-08 0 2.1e-08 0 2.1003e-08 0.0007 2.1006e-08 0 2.106e-08 0 2.1063e-08 0.0007 2.1066e-08 0 2.112e-08 0 2.1123e-08 0.0007 2.1126e-08 0 2.118e-08 0 2.1183e-08 0.0007 2.1186e-08 0 2.124e-08 0 2.1243e-08 0.0007 2.1246e-08 0 2.13e-08 0 2.1303e-08 0.0007 2.1306e-08 0 2.136e-08 0 2.1363e-08 0.0007 2.1366e-08 0 2.142e-08 0 2.1423e-08 0.0007 2.1426e-08 0 2.148e-08 0 2.1483e-08 0.0007 2.1486e-08 0 2.154e-08 0 2.1543e-08 0.0007 2.1546e-08 0 2.16e-08 0 2.1603e-08 0.0007 2.1606e-08 0 2.166e-08 0 2.1663e-08 0.0007 2.1666e-08 0 2.172e-08 0 2.1723e-08 0.0007 2.1726e-08 0 2.178e-08 0 2.1783e-08 0.0007 2.1786e-08 0 2.184e-08 0 2.1843e-08 0.0007 2.1846e-08 0 2.19e-08 0 2.1903e-08 0.0007 2.1906e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.202e-08 0 2.2023e-08 0.0007 2.2026e-08 0 2.208e-08 0 2.2083e-08 0.0007 2.2086e-08 0 2.214e-08 0 2.2143e-08 0.0007 2.2146e-08 0 2.22e-08 0 2.2203e-08 0.0007 2.2206e-08 0 2.226e-08 0 2.2263e-08 0.0007 2.2266e-08 0 2.232e-08 0 2.2323e-08 0.0007 2.2326e-08 0 2.238e-08 0 2.2383e-08 0.0007 2.2386e-08 0 2.244e-08 0 2.2443e-08 0.0007 2.2446e-08 0 2.25e-08 0 2.2503e-08 0.0007 2.2506e-08 0 2.256e-08 0 2.2563e-08 0.0007 2.2566e-08 0 2.262e-08 0 2.2623e-08 0.0007 2.2626e-08 0 2.268e-08 0 2.2683e-08 0.0007 2.2686e-08 0 2.274e-08 0 2.2743e-08 0.0007 2.2746e-08 0 2.28e-08 0 2.2803e-08 0.0007 2.2806e-08 0 2.286e-08 0 2.2863e-08 0.0007 2.2866e-08 0 2.292e-08 0 2.2923e-08 0.0007 2.2926e-08 0 2.298e-08 0 2.2983e-08 0.0007 2.2986e-08 0 2.304e-08 0 2.3043e-08 0.0007 2.3046e-08 0 2.31e-08 0 2.3103e-08 0.0007 2.3106e-08 0 2.316e-08 0 2.3163e-08 0.0007 2.3166e-08 0 2.322e-08 0 2.3223e-08 0.0007 2.3226e-08 0 2.328e-08 0 2.3283e-08 0.0007 2.3286e-08 0 2.334e-08 0 2.3343e-08 0.0007 2.3346e-08 0 2.34e-08 0 2.3403e-08 0.0007 2.3406e-08 0 2.346e-08 0 2.3463e-08 0.0007 2.3466e-08 0 2.352e-08 0 2.3523e-08 0.0007 2.3526e-08 0 2.358e-08 0 2.3583e-08 0.0007 2.3586e-08 0 2.364e-08 0 2.3643e-08 0.0007 2.3646e-08 0 2.37e-08 0 2.3703e-08 0.0007 2.3706e-08 0 2.376e-08 0 2.3763e-08 0.0007 2.3766e-08 0 2.382e-08 0 2.3823e-08 0.0007 2.3826e-08 0 2.388e-08 0 2.3883e-08 0.0007 2.3886e-08 0)
L_S0|1 P0_2_RX _S0|A1  2.067833848e-12
L_S0|2 _S0|A1 _S0|A2  4.135667696e-12
L_S0|3 _S0|A3 _S0|A4  8.271335392e-12
L_S0|T T12 _S0|T1  2.067833848e-12
L_S0|4 _S0|T1 _S0|T2  4.135667696e-12
L_S0|5 _S0|A4 _S0|Q1  4.135667696e-12
L_S0|6 _S0|Q1 S0  2.067833848e-12
IT13|T 0 T13  PWL(0 0 0 0 3e-12 0.0007 6e-12 0 6e-11 0 6.3e-11 0.0007 6.6e-11 0 1.2e-10 0 1.23e-10 0.0007 1.26e-10 0 1.8e-10 0 1.83e-10 0.0007 1.86e-10 0 2.4e-10 0 2.43e-10 0.0007 2.46e-10 0 3e-10 0 3.03e-10 0.0007 3.06e-10 0 3.6e-10 0 3.63e-10 0.0007 3.66e-10 0 4.2e-10 0 4.23e-10 0.0007 4.26e-10 0 4.8e-10 0 4.83e-10 0.0007 4.86e-10 0 5.4e-10 0 5.43e-10 0.0007 5.46e-10 0 6e-10 0 6.03e-10 0.0007 6.06e-10 0 6.6e-10 0 6.63e-10 0.0007 6.66e-10 0 7.2e-10 0 7.23e-10 0.0007 7.26e-10 0 7.8e-10 0 7.83e-10 0.0007 7.86e-10 0 8.4e-10 0 8.43e-10 0.0007 8.46e-10 0 9e-10 0 9.03e-10 0.0007 9.06e-10 0 9.6e-10 0 9.63e-10 0.0007 9.66e-10 0 1.02e-09 0 1.023e-09 0.0007 1.026e-09 0 1.08e-09 0 1.083e-09 0.0007 1.086e-09 0 1.14e-09 0 1.143e-09 0.0007 1.146e-09 0 1.2e-09 0 1.203e-09 0.0007 1.206e-09 0 1.26e-09 0 1.263e-09 0.0007 1.266e-09 0 1.32e-09 0 1.323e-09 0.0007 1.326e-09 0 1.38e-09 0 1.383e-09 0.0007 1.386e-09 0 1.44e-09 0 1.443e-09 0.0007 1.446e-09 0 1.5e-09 0 1.503e-09 0.0007 1.506e-09 0 1.56e-09 0 1.563e-09 0.0007 1.566e-09 0 1.62e-09 0 1.623e-09 0.0007 1.626e-09 0 1.68e-09 0 1.683e-09 0.0007 1.686e-09 0 1.74e-09 0 1.743e-09 0.0007 1.746e-09 0 1.8e-09 0 1.803e-09 0.0007 1.806e-09 0 1.86e-09 0 1.863e-09 0.0007 1.866e-09 0 1.92e-09 0 1.923e-09 0.0007 1.926e-09 0 1.98e-09 0 1.983e-09 0.0007 1.986e-09 0 2.04e-09 0 2.043e-09 0.0007 2.046e-09 0 2.1e-09 0 2.103e-09 0.0007 2.106e-09 0 2.16e-09 0 2.163e-09 0.0007 2.166e-09 0 2.22e-09 0 2.223e-09 0.0007 2.226e-09 0 2.28e-09 0 2.283e-09 0.0007 2.286e-09 0 2.34e-09 0 2.343e-09 0.0007 2.346e-09 0 2.4e-09 0 2.403e-09 0.0007 2.406e-09 0 2.46e-09 0 2.463e-09 0.0007 2.466e-09 0 2.52e-09 0 2.523e-09 0.0007 2.526e-09 0 2.58e-09 0 2.583e-09 0.0007 2.586e-09 0 2.64e-09 0 2.643e-09 0.0007 2.646e-09 0 2.7e-09 0 2.703e-09 0.0007 2.706e-09 0 2.76e-09 0 2.763e-09 0.0007 2.766e-09 0 2.82e-09 0 2.823e-09 0.0007 2.826e-09 0 2.88e-09 0 2.883e-09 0.0007 2.886e-09 0 2.94e-09 0 2.943e-09 0.0007 2.946e-09 0 3e-09 0 3.003e-09 0.0007 3.006e-09 0 3.06e-09 0 3.063e-09 0.0007 3.066e-09 0 3.12e-09 0 3.123e-09 0.0007 3.126e-09 0 3.18e-09 0 3.183e-09 0.0007 3.186e-09 0 3.24e-09 0 3.243e-09 0.0007 3.246e-09 0 3.3e-09 0 3.303e-09 0.0007 3.306e-09 0 3.36e-09 0 3.363e-09 0.0007 3.366e-09 0 3.42e-09 0 3.423e-09 0.0007 3.426e-09 0 3.48e-09 0 3.483e-09 0.0007 3.486e-09 0 3.54e-09 0 3.543e-09 0.0007 3.546e-09 0 3.6e-09 0 3.603e-09 0.0007 3.606e-09 0 3.66e-09 0 3.663e-09 0.0007 3.666e-09 0 3.72e-09 0 3.723e-09 0.0007 3.726e-09 0 3.78e-09 0 3.783e-09 0.0007 3.786e-09 0 3.84e-09 0 3.843e-09 0.0007 3.846e-09 0 3.9e-09 0 3.903e-09 0.0007 3.906e-09 0 3.96e-09 0 3.963e-09 0.0007 3.966e-09 0 4.02e-09 0 4.023e-09 0.0007 4.026e-09 0 4.08e-09 0 4.083e-09 0.0007 4.086e-09 0 4.14e-09 0 4.143e-09 0.0007 4.146e-09 0 4.2e-09 0 4.203e-09 0.0007 4.206e-09 0 4.26e-09 0 4.263e-09 0.0007 4.266e-09 0 4.32e-09 0 4.323e-09 0.0007 4.326e-09 0 4.38e-09 0 4.383e-09 0.0007 4.386e-09 0 4.44e-09 0 4.443e-09 0.0007 4.446e-09 0 4.5e-09 0 4.503e-09 0.0007 4.506e-09 0 4.56e-09 0 4.563e-09 0.0007 4.566e-09 0 4.62e-09 0 4.623e-09 0.0007 4.626e-09 0 4.68e-09 0 4.683e-09 0.0007 4.686e-09 0 4.74e-09 0 4.743e-09 0.0007 4.746e-09 0 4.8e-09 0 4.803e-09 0.0007 4.806e-09 0 4.86e-09 0 4.863e-09 0.0007 4.866e-09 0 4.92e-09 0 4.923e-09 0.0007 4.926e-09 0 4.98e-09 0 4.983e-09 0.0007 4.986e-09 0 5.04e-09 0 5.043e-09 0.0007 5.046e-09 0 5.1e-09 0 5.103e-09 0.0007 5.106e-09 0 5.16e-09 0 5.163e-09 0.0007 5.166e-09 0 5.22e-09 0 5.223e-09 0.0007 5.226e-09 0 5.28e-09 0 5.283e-09 0.0007 5.286e-09 0 5.34e-09 0 5.343e-09 0.0007 5.346e-09 0 5.4e-09 0 5.403e-09 0.0007 5.406e-09 0 5.46e-09 0 5.463e-09 0.0007 5.466e-09 0 5.52e-09 0 5.523e-09 0.0007 5.526e-09 0 5.58e-09 0 5.583e-09 0.0007 5.586e-09 0 5.64e-09 0 5.643e-09 0.0007 5.646e-09 0 5.7e-09 0 5.703e-09 0.0007 5.706e-09 0 5.76e-09 0 5.763e-09 0.0007 5.766e-09 0 5.82e-09 0 5.823e-09 0.0007 5.826e-09 0 5.88e-09 0 5.883e-09 0.0007 5.886e-09 0 5.94e-09 0 5.943e-09 0.0007 5.946e-09 0 6e-09 0 6.003e-09 0.0007 6.006e-09 0 6.06e-09 0 6.063e-09 0.0007 6.066e-09 0 6.12e-09 0 6.123e-09 0.0007 6.126e-09 0 6.18e-09 0 6.183e-09 0.0007 6.186e-09 0 6.24e-09 0 6.243e-09 0.0007 6.246e-09 0 6.3e-09 0 6.303e-09 0.0007 6.306e-09 0 6.36e-09 0 6.363e-09 0.0007 6.366e-09 0 6.42e-09 0 6.423e-09 0.0007 6.426e-09 0 6.48e-09 0 6.483e-09 0.0007 6.486e-09 0 6.54e-09 0 6.543e-09 0.0007 6.546e-09 0 6.6e-09 0 6.603e-09 0.0007 6.606e-09 0 6.66e-09 0 6.663e-09 0.0007 6.666e-09 0 6.72e-09 0 6.723e-09 0.0007 6.726e-09 0 6.78e-09 0 6.783e-09 0.0007 6.786e-09 0 6.84e-09 0 6.843e-09 0.0007 6.846e-09 0 6.9e-09 0 6.903e-09 0.0007 6.906e-09 0 6.96e-09 0 6.963e-09 0.0007 6.966e-09 0 7.02e-09 0 7.023e-09 0.0007 7.026e-09 0 7.08e-09 0 7.083e-09 0.0007 7.086e-09 0 7.14e-09 0 7.143e-09 0.0007 7.146e-09 0 7.2e-09 0 7.203e-09 0.0007 7.206e-09 0 7.26e-09 0 7.263e-09 0.0007 7.266e-09 0 7.32e-09 0 7.323e-09 0.0007 7.326e-09 0 7.38e-09 0 7.383e-09 0.0007 7.386e-09 0 7.44e-09 0 7.443e-09 0.0007 7.446e-09 0 7.5e-09 0 7.503e-09 0.0007 7.506e-09 0 7.56e-09 0 7.563e-09 0.0007 7.566e-09 0 7.62e-09 0 7.623e-09 0.0007 7.626e-09 0 7.68e-09 0 7.683e-09 0.0007 7.686e-09 0 7.74e-09 0 7.743e-09 0.0007 7.746e-09 0 7.8e-09 0 7.803e-09 0.0007 7.806e-09 0 7.86e-09 0 7.863e-09 0.0007 7.866e-09 0 7.92e-09 0 7.923e-09 0.0007 7.926e-09 0 7.98e-09 0 7.983e-09 0.0007 7.986e-09 0 8.04e-09 0 8.043e-09 0.0007 8.046e-09 0 8.1e-09 0 8.103e-09 0.0007 8.106e-09 0 8.16e-09 0 8.163e-09 0.0007 8.166e-09 0 8.22e-09 0 8.223e-09 0.0007 8.226e-09 0 8.28e-09 0 8.283e-09 0.0007 8.286e-09 0 8.34e-09 0 8.343e-09 0.0007 8.346e-09 0 8.4e-09 0 8.403e-09 0.0007 8.406e-09 0 8.46e-09 0 8.463e-09 0.0007 8.466e-09 0 8.52e-09 0 8.523e-09 0.0007 8.526e-09 0 8.58e-09 0 8.583e-09 0.0007 8.586e-09 0 8.64e-09 0 8.643e-09 0.0007 8.646e-09 0 8.7e-09 0 8.703e-09 0.0007 8.706e-09 0 8.76e-09 0 8.763e-09 0.0007 8.766e-09 0 8.82e-09 0 8.823e-09 0.0007 8.826e-09 0 8.88e-09 0 8.883e-09 0.0007 8.886e-09 0 8.94e-09 0 8.943e-09 0.0007 8.946e-09 0 9e-09 0 9.003e-09 0.0007 9.006e-09 0 9.06e-09 0 9.063e-09 0.0007 9.066e-09 0 9.12e-09 0 9.123e-09 0.0007 9.126e-09 0 9.18e-09 0 9.183e-09 0.0007 9.186e-09 0 9.24e-09 0 9.243e-09 0.0007 9.246e-09 0 9.3e-09 0 9.303e-09 0.0007 9.306e-09 0 9.36e-09 0 9.363e-09 0.0007 9.366e-09 0 9.42e-09 0 9.423e-09 0.0007 9.426e-09 0 9.48e-09 0 9.483e-09 0.0007 9.486e-09 0 9.54e-09 0 9.543e-09 0.0007 9.546e-09 0 9.6e-09 0 9.603e-09 0.0007 9.606e-09 0 9.66e-09 0 9.663e-09 0.0007 9.666e-09 0 9.72e-09 0 9.723e-09 0.0007 9.726e-09 0 9.78e-09 0 9.783e-09 0.0007 9.786e-09 0 9.84e-09 0 9.843e-09 0.0007 9.846e-09 0 9.9e-09 0 9.903e-09 0.0007 9.906e-09 0 9.96e-09 0 9.963e-09 0.0007 9.966e-09 0 1.002e-08 0 1.0023e-08 0.0007 1.0026e-08 0 1.008e-08 0 1.0083e-08 0.0007 1.0086e-08 0 1.014e-08 0 1.0143e-08 0.0007 1.0146e-08 0 1.02e-08 0 1.0203e-08 0.0007 1.0206e-08 0 1.026e-08 0 1.0263e-08 0.0007 1.0266e-08 0 1.032e-08 0 1.0323e-08 0.0007 1.0326e-08 0 1.038e-08 0 1.0383e-08 0.0007 1.0386e-08 0 1.044e-08 0 1.0443e-08 0.0007 1.0446e-08 0 1.05e-08 0 1.0503e-08 0.0007 1.0506e-08 0 1.056e-08 0 1.0563e-08 0.0007 1.0566e-08 0 1.062e-08 0 1.0623e-08 0.0007 1.0626e-08 0 1.068e-08 0 1.0683e-08 0.0007 1.0686e-08 0 1.074e-08 0 1.0743e-08 0.0007 1.0746e-08 0 1.08e-08 0 1.0803e-08 0.0007 1.0806e-08 0 1.086e-08 0 1.0863e-08 0.0007 1.0866e-08 0 1.092e-08 0 1.0923e-08 0.0007 1.0926e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.104e-08 0 1.1043e-08 0.0007 1.1046e-08 0 1.11e-08 0 1.1103e-08 0.0007 1.1106e-08 0 1.116e-08 0 1.1163e-08 0.0007 1.1166e-08 0 1.122e-08 0 1.1223e-08 0.0007 1.1226e-08 0 1.128e-08 0 1.1283e-08 0.0007 1.1286e-08 0 1.134e-08 0 1.1343e-08 0.0007 1.1346e-08 0 1.14e-08 0 1.1403e-08 0.0007 1.1406e-08 0 1.146e-08 0 1.1463e-08 0.0007 1.1466e-08 0 1.152e-08 0 1.1523e-08 0.0007 1.1526e-08 0 1.158e-08 0 1.1583e-08 0.0007 1.1586e-08 0 1.164e-08 0 1.1643e-08 0.0007 1.1646e-08 0 1.17e-08 0 1.1703e-08 0.0007 1.1706e-08 0 1.176e-08 0 1.1763e-08 0.0007 1.1766e-08 0 1.182e-08 0 1.1823e-08 0.0007 1.1826e-08 0 1.188e-08 0 1.1883e-08 0.0007 1.1886e-08 0 1.194e-08 0 1.1943e-08 0.0007 1.1946e-08 0 1.2e-08 0 1.2003e-08 0.0007 1.2006e-08 0 1.206e-08 0 1.2063e-08 0.0007 1.2066e-08 0 1.212e-08 0 1.2123e-08 0.0007 1.2126e-08 0 1.218e-08 0 1.2183e-08 0.0007 1.2186e-08 0 1.224e-08 0 1.2243e-08 0.0007 1.2246e-08 0 1.23e-08 0 1.2303e-08 0.0007 1.2306e-08 0 1.236e-08 0 1.2363e-08 0.0007 1.2366e-08 0 1.242e-08 0 1.2423e-08 0.0007 1.2426e-08 0 1.248e-08 0 1.2483e-08 0.0007 1.2486e-08 0 1.254e-08 0 1.2543e-08 0.0007 1.2546e-08 0 1.26e-08 0 1.2603e-08 0.0007 1.2606e-08 0 1.266e-08 0 1.2663e-08 0.0007 1.2666e-08 0 1.272e-08 0 1.2723e-08 0.0007 1.2726e-08 0 1.278e-08 0 1.2783e-08 0.0007 1.2786e-08 0 1.284e-08 0 1.2843e-08 0.0007 1.2846e-08 0 1.29e-08 0 1.2903e-08 0.0007 1.2906e-08 0 1.296e-08 0 1.2963e-08 0.0007 1.2966e-08 0 1.302e-08 0 1.3023e-08 0.0007 1.3026e-08 0 1.308e-08 0 1.3083e-08 0.0007 1.3086e-08 0 1.314e-08 0 1.3143e-08 0.0007 1.3146e-08 0 1.32e-08 0 1.3203e-08 0.0007 1.3206e-08 0 1.326e-08 0 1.3263e-08 0.0007 1.3266e-08 0 1.332e-08 0 1.3323e-08 0.0007 1.3326e-08 0 1.338e-08 0 1.3383e-08 0.0007 1.3386e-08 0 1.344e-08 0 1.3443e-08 0.0007 1.3446e-08 0 1.35e-08 0 1.3503e-08 0.0007 1.3506e-08 0 1.356e-08 0 1.3563e-08 0.0007 1.3566e-08 0 1.362e-08 0 1.3623e-08 0.0007 1.3626e-08 0 1.368e-08 0 1.3683e-08 0.0007 1.3686e-08 0 1.374e-08 0 1.3743e-08 0.0007 1.3746e-08 0 1.38e-08 0 1.3803e-08 0.0007 1.3806e-08 0 1.386e-08 0 1.3863e-08 0.0007 1.3866e-08 0 1.392e-08 0 1.3923e-08 0.0007 1.3926e-08 0 1.398e-08 0 1.3983e-08 0.0007 1.3986e-08 0 1.404e-08 0 1.4043e-08 0.0007 1.4046e-08 0 1.41e-08 0 1.4103e-08 0.0007 1.4106e-08 0 1.416e-08 0 1.4163e-08 0.0007 1.4166e-08 0 1.422e-08 0 1.4223e-08 0.0007 1.4226e-08 0 1.428e-08 0 1.4283e-08 0.0007 1.4286e-08 0 1.434e-08 0 1.4343e-08 0.0007 1.4346e-08 0 1.44e-08 0 1.4403e-08 0.0007 1.4406e-08 0 1.446e-08 0 1.4463e-08 0.0007 1.4466e-08 0 1.452e-08 0 1.4523e-08 0.0007 1.4526e-08 0 1.458e-08 0 1.4583e-08 0.0007 1.4586e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.47e-08 0 1.4703e-08 0.0007 1.4706e-08 0 1.476e-08 0 1.4763e-08 0.0007 1.4766e-08 0 1.482e-08 0 1.4823e-08 0.0007 1.4826e-08 0 1.488e-08 0 1.4883e-08 0.0007 1.4886e-08 0 1.494e-08 0 1.4943e-08 0.0007 1.4946e-08 0 1.5e-08 0 1.5003e-08 0.0007 1.5006e-08 0 1.506e-08 0 1.5063e-08 0.0007 1.5066e-08 0 1.512e-08 0 1.5123e-08 0.0007 1.5126e-08 0 1.518e-08 0 1.5183e-08 0.0007 1.5186e-08 0 1.524e-08 0 1.5243e-08 0.0007 1.5246e-08 0 1.53e-08 0 1.5303e-08 0.0007 1.5306e-08 0 1.536e-08 0 1.5363e-08 0.0007 1.5366e-08 0 1.542e-08 0 1.5423e-08 0.0007 1.5426e-08 0 1.548e-08 0 1.5483e-08 0.0007 1.5486e-08 0 1.554e-08 0 1.5543e-08 0.0007 1.5546e-08 0 1.56e-08 0 1.5603e-08 0.0007 1.5606e-08 0 1.566e-08 0 1.5663e-08 0.0007 1.5666e-08 0 1.572e-08 0 1.5723e-08 0.0007 1.5726e-08 0 1.578e-08 0 1.5783e-08 0.0007 1.5786e-08 0 1.584e-08 0 1.5843e-08 0.0007 1.5846e-08 0 1.59e-08 0 1.5903e-08 0.0007 1.5906e-08 0 1.596e-08 0 1.5963e-08 0.0007 1.5966e-08 0 1.602e-08 0 1.6023e-08 0.0007 1.6026e-08 0 1.608e-08 0 1.6083e-08 0.0007 1.6086e-08 0 1.614e-08 0 1.6143e-08 0.0007 1.6146e-08 0 1.62e-08 0 1.6203e-08 0.0007 1.6206e-08 0 1.626e-08 0 1.6263e-08 0.0007 1.6266e-08 0 1.632e-08 0 1.6323e-08 0.0007 1.6326e-08 0 1.638e-08 0 1.6383e-08 0.0007 1.6386e-08 0 1.644e-08 0 1.6443e-08 0.0007 1.6446e-08 0 1.65e-08 0 1.6503e-08 0.0007 1.6506e-08 0 1.656e-08 0 1.6563e-08 0.0007 1.6566e-08 0 1.662e-08 0 1.6623e-08 0.0007 1.6626e-08 0 1.668e-08 0 1.6683e-08 0.0007 1.6686e-08 0 1.674e-08 0 1.6743e-08 0.0007 1.6746e-08 0 1.68e-08 0 1.6803e-08 0.0007 1.6806e-08 0 1.686e-08 0 1.6863e-08 0.0007 1.6866e-08 0 1.692e-08 0 1.6923e-08 0.0007 1.6926e-08 0 1.698e-08 0 1.6983e-08 0.0007 1.6986e-08 0 1.704e-08 0 1.7043e-08 0.0007 1.7046e-08 0 1.71e-08 0 1.7103e-08 0.0007 1.7106e-08 0 1.716e-08 0 1.7163e-08 0.0007 1.7166e-08 0 1.722e-08 0 1.7223e-08 0.0007 1.7226e-08 0 1.728e-08 0 1.7283e-08 0.0007 1.7286e-08 0 1.734e-08 0 1.7343e-08 0.0007 1.7346e-08 0 1.74e-08 0 1.7403e-08 0.0007 1.7406e-08 0 1.746e-08 0 1.7463e-08 0.0007 1.7466e-08 0 1.752e-08 0 1.7523e-08 0.0007 1.7526e-08 0 1.758e-08 0 1.7583e-08 0.0007 1.7586e-08 0 1.764e-08 0 1.7643e-08 0.0007 1.7646e-08 0 1.77e-08 0 1.7703e-08 0.0007 1.7706e-08 0 1.776e-08 0 1.7763e-08 0.0007 1.7766e-08 0 1.782e-08 0 1.7823e-08 0.0007 1.7826e-08 0 1.788e-08 0 1.7883e-08 0.0007 1.7886e-08 0 1.794e-08 0 1.7943e-08 0.0007 1.7946e-08 0 1.8e-08 0 1.8003e-08 0.0007 1.8006e-08 0 1.806e-08 0 1.8063e-08 0.0007 1.8066e-08 0 1.812e-08 0 1.8123e-08 0.0007 1.8126e-08 0 1.818e-08 0 1.8183e-08 0.0007 1.8186e-08 0 1.824e-08 0 1.8243e-08 0.0007 1.8246e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.836e-08 0 1.8363e-08 0.0007 1.8366e-08 0 1.842e-08 0 1.8423e-08 0.0007 1.8426e-08 0 1.848e-08 0 1.8483e-08 0.0007 1.8486e-08 0 1.854e-08 0 1.8543e-08 0.0007 1.8546e-08 0 1.86e-08 0 1.8603e-08 0.0007 1.8606e-08 0 1.866e-08 0 1.8663e-08 0.0007 1.8666e-08 0 1.872e-08 0 1.8723e-08 0.0007 1.8726e-08 0 1.878e-08 0 1.8783e-08 0.0007 1.8786e-08 0 1.884e-08 0 1.8843e-08 0.0007 1.8846e-08 0 1.89e-08 0 1.8903e-08 0.0007 1.8906e-08 0 1.896e-08 0 1.8963e-08 0.0007 1.8966e-08 0 1.902e-08 0 1.9023e-08 0.0007 1.9026e-08 0 1.908e-08 0 1.9083e-08 0.0007 1.9086e-08 0 1.914e-08 0 1.9143e-08 0.0007 1.9146e-08 0 1.92e-08 0 1.9203e-08 0.0007 1.9206e-08 0 1.926e-08 0 1.9263e-08 0.0007 1.9266e-08 0 1.932e-08 0 1.9323e-08 0.0007 1.9326e-08 0 1.938e-08 0 1.9383e-08 0.0007 1.9386e-08 0 1.944e-08 0 1.9443e-08 0.0007 1.9446e-08 0 1.95e-08 0 1.9503e-08 0.0007 1.9506e-08 0 1.956e-08 0 1.9563e-08 0.0007 1.9566e-08 0 1.962e-08 0 1.9623e-08 0.0007 1.9626e-08 0 1.968e-08 0 1.9683e-08 0.0007 1.9686e-08 0 1.974e-08 0 1.9743e-08 0.0007 1.9746e-08 0 1.98e-08 0 1.9803e-08 0.0007 1.9806e-08 0 1.986e-08 0 1.9863e-08 0.0007 1.9866e-08 0 1.992e-08 0 1.9923e-08 0.0007 1.9926e-08 0 1.998e-08 0 1.9983e-08 0.0007 1.9986e-08 0 2.004e-08 0 2.0043e-08 0.0007 2.0046e-08 0 2.01e-08 0 2.0103e-08 0.0007 2.0106e-08 0 2.016e-08 0 2.0163e-08 0.0007 2.0166e-08 0 2.022e-08 0 2.0223e-08 0.0007 2.0226e-08 0 2.028e-08 0 2.0283e-08 0.0007 2.0286e-08 0 2.034e-08 0 2.0343e-08 0.0007 2.0346e-08 0 2.04e-08 0 2.0403e-08 0.0007 2.0406e-08 0 2.046e-08 0 2.0463e-08 0.0007 2.0466e-08 0 2.052e-08 0 2.0523e-08 0.0007 2.0526e-08 0 2.058e-08 0 2.0583e-08 0.0007 2.0586e-08 0 2.064e-08 0 2.0643e-08 0.0007 2.0646e-08 0 2.07e-08 0 2.0703e-08 0.0007 2.0706e-08 0 2.076e-08 0 2.0763e-08 0.0007 2.0766e-08 0 2.082e-08 0 2.0823e-08 0.0007 2.0826e-08 0 2.088e-08 0 2.0883e-08 0.0007 2.0886e-08 0 2.094e-08 0 2.0943e-08 0.0007 2.0946e-08 0 2.1e-08 0 2.1003e-08 0.0007 2.1006e-08 0 2.106e-08 0 2.1063e-08 0.0007 2.1066e-08 0 2.112e-08 0 2.1123e-08 0.0007 2.1126e-08 0 2.118e-08 0 2.1183e-08 0.0007 2.1186e-08 0 2.124e-08 0 2.1243e-08 0.0007 2.1246e-08 0 2.13e-08 0 2.1303e-08 0.0007 2.1306e-08 0 2.136e-08 0 2.1363e-08 0.0007 2.1366e-08 0 2.142e-08 0 2.1423e-08 0.0007 2.1426e-08 0 2.148e-08 0 2.1483e-08 0.0007 2.1486e-08 0 2.154e-08 0 2.1543e-08 0.0007 2.1546e-08 0 2.16e-08 0 2.1603e-08 0.0007 2.1606e-08 0 2.166e-08 0 2.1663e-08 0.0007 2.1666e-08 0 2.172e-08 0 2.1723e-08 0.0007 2.1726e-08 0 2.178e-08 0 2.1783e-08 0.0007 2.1786e-08 0 2.184e-08 0 2.1843e-08 0.0007 2.1846e-08 0 2.19e-08 0 2.1903e-08 0.0007 2.1906e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.202e-08 0 2.2023e-08 0.0007 2.2026e-08 0 2.208e-08 0 2.2083e-08 0.0007 2.2086e-08 0 2.214e-08 0 2.2143e-08 0.0007 2.2146e-08 0 2.22e-08 0 2.2203e-08 0.0007 2.2206e-08 0 2.226e-08 0 2.2263e-08 0.0007 2.2266e-08 0 2.232e-08 0 2.2323e-08 0.0007 2.2326e-08 0 2.238e-08 0 2.2383e-08 0.0007 2.2386e-08 0 2.244e-08 0 2.2443e-08 0.0007 2.2446e-08 0 2.25e-08 0 2.2503e-08 0.0007 2.2506e-08 0 2.256e-08 0 2.2563e-08 0.0007 2.2566e-08 0 2.262e-08 0 2.2623e-08 0.0007 2.2626e-08 0 2.268e-08 0 2.2683e-08 0.0007 2.2686e-08 0 2.274e-08 0 2.2743e-08 0.0007 2.2746e-08 0 2.28e-08 0 2.2803e-08 0.0007 2.2806e-08 0 2.286e-08 0 2.2863e-08 0.0007 2.2866e-08 0 2.292e-08 0 2.2923e-08 0.0007 2.2926e-08 0 2.298e-08 0 2.2983e-08 0.0007 2.2986e-08 0 2.304e-08 0 2.3043e-08 0.0007 2.3046e-08 0 2.31e-08 0 2.3103e-08 0.0007 2.3106e-08 0 2.316e-08 0 2.3163e-08 0.0007 2.3166e-08 0 2.322e-08 0 2.3223e-08 0.0007 2.3226e-08 0 2.328e-08 0 2.3283e-08 0.0007 2.3286e-08 0 2.334e-08 0 2.3343e-08 0.0007 2.3346e-08 0 2.34e-08 0 2.3403e-08 0.0007 2.3406e-08 0 2.346e-08 0 2.3463e-08 0.0007 2.3466e-08 0 2.352e-08 0 2.3523e-08 0.0007 2.3526e-08 0 2.358e-08 0 2.3583e-08 0.0007 2.3586e-08 0 2.364e-08 0 2.3643e-08 0.0007 2.3646e-08 0 2.37e-08 0 2.3703e-08 0.0007 2.3706e-08 0 2.376e-08 0 2.3763e-08 0.0007 2.3766e-08 0 2.382e-08 0 2.3823e-08 0.0007 2.3826e-08 0 2.388e-08 0 2.3883e-08 0.0007 2.3886e-08 0)
L_S1|A1 G0_2_RX _S1|A1  2.067833848e-12
L_S1|A2 _S1|A1 _S1|A2  4.135667696e-12
L_S1|A3 _S1|A3 _S1|AB  8.271335392e-12
L_S1|B1 IP1_2_OUT_RX _S1|B1  2.067833848e-12
L_S1|B2 _S1|B1 _S1|B2  4.135667696e-12
L_S1|B3 _S1|B3 _S1|AB  8.271335392e-12
L_S1|T1 T13 _S1|T1  2.067833848e-12
L_S1|T2 _S1|T1 _S1|T2  4.135667696e-12
L_S1|Q2 _S1|ABTQ _S1|Q1  4.135667696e-12
L_S1|Q1 _S1|Q1 S1  2.067833848e-12
IT14|T 0 T14  PWL(0 0 0 0 3e-12 0.0007 6e-12 0 6e-11 0 6.3e-11 0.0007 6.6e-11 0 1.2e-10 0 1.23e-10 0.0007 1.26e-10 0 1.8e-10 0 1.83e-10 0.0007 1.86e-10 0 2.4e-10 0 2.43e-10 0.0007 2.46e-10 0 3e-10 0 3.03e-10 0.0007 3.06e-10 0 3.6e-10 0 3.63e-10 0.0007 3.66e-10 0 4.2e-10 0 4.23e-10 0.0007 4.26e-10 0 4.8e-10 0 4.83e-10 0.0007 4.86e-10 0 5.4e-10 0 5.43e-10 0.0007 5.46e-10 0 6e-10 0 6.03e-10 0.0007 6.06e-10 0 6.6e-10 0 6.63e-10 0.0007 6.66e-10 0 7.2e-10 0 7.23e-10 0.0007 7.26e-10 0 7.8e-10 0 7.83e-10 0.0007 7.86e-10 0 8.4e-10 0 8.43e-10 0.0007 8.46e-10 0 9e-10 0 9.03e-10 0.0007 9.06e-10 0 9.6e-10 0 9.63e-10 0.0007 9.66e-10 0 1.02e-09 0 1.023e-09 0.0007 1.026e-09 0 1.08e-09 0 1.083e-09 0.0007 1.086e-09 0 1.14e-09 0 1.143e-09 0.0007 1.146e-09 0 1.2e-09 0 1.203e-09 0.0007 1.206e-09 0 1.26e-09 0 1.263e-09 0.0007 1.266e-09 0 1.32e-09 0 1.323e-09 0.0007 1.326e-09 0 1.38e-09 0 1.383e-09 0.0007 1.386e-09 0 1.44e-09 0 1.443e-09 0.0007 1.446e-09 0 1.5e-09 0 1.503e-09 0.0007 1.506e-09 0 1.56e-09 0 1.563e-09 0.0007 1.566e-09 0 1.62e-09 0 1.623e-09 0.0007 1.626e-09 0 1.68e-09 0 1.683e-09 0.0007 1.686e-09 0 1.74e-09 0 1.743e-09 0.0007 1.746e-09 0 1.8e-09 0 1.803e-09 0.0007 1.806e-09 0 1.86e-09 0 1.863e-09 0.0007 1.866e-09 0 1.92e-09 0 1.923e-09 0.0007 1.926e-09 0 1.98e-09 0 1.983e-09 0.0007 1.986e-09 0 2.04e-09 0 2.043e-09 0.0007 2.046e-09 0 2.1e-09 0 2.103e-09 0.0007 2.106e-09 0 2.16e-09 0 2.163e-09 0.0007 2.166e-09 0 2.22e-09 0 2.223e-09 0.0007 2.226e-09 0 2.28e-09 0 2.283e-09 0.0007 2.286e-09 0 2.34e-09 0 2.343e-09 0.0007 2.346e-09 0 2.4e-09 0 2.403e-09 0.0007 2.406e-09 0 2.46e-09 0 2.463e-09 0.0007 2.466e-09 0 2.52e-09 0 2.523e-09 0.0007 2.526e-09 0 2.58e-09 0 2.583e-09 0.0007 2.586e-09 0 2.64e-09 0 2.643e-09 0.0007 2.646e-09 0 2.7e-09 0 2.703e-09 0.0007 2.706e-09 0 2.76e-09 0 2.763e-09 0.0007 2.766e-09 0 2.82e-09 0 2.823e-09 0.0007 2.826e-09 0 2.88e-09 0 2.883e-09 0.0007 2.886e-09 0 2.94e-09 0 2.943e-09 0.0007 2.946e-09 0 3e-09 0 3.003e-09 0.0007 3.006e-09 0 3.06e-09 0 3.063e-09 0.0007 3.066e-09 0 3.12e-09 0 3.123e-09 0.0007 3.126e-09 0 3.18e-09 0 3.183e-09 0.0007 3.186e-09 0 3.24e-09 0 3.243e-09 0.0007 3.246e-09 0 3.3e-09 0 3.303e-09 0.0007 3.306e-09 0 3.36e-09 0 3.363e-09 0.0007 3.366e-09 0 3.42e-09 0 3.423e-09 0.0007 3.426e-09 0 3.48e-09 0 3.483e-09 0.0007 3.486e-09 0 3.54e-09 0 3.543e-09 0.0007 3.546e-09 0 3.6e-09 0 3.603e-09 0.0007 3.606e-09 0 3.66e-09 0 3.663e-09 0.0007 3.666e-09 0 3.72e-09 0 3.723e-09 0.0007 3.726e-09 0 3.78e-09 0 3.783e-09 0.0007 3.786e-09 0 3.84e-09 0 3.843e-09 0.0007 3.846e-09 0 3.9e-09 0 3.903e-09 0.0007 3.906e-09 0 3.96e-09 0 3.963e-09 0.0007 3.966e-09 0 4.02e-09 0 4.023e-09 0.0007 4.026e-09 0 4.08e-09 0 4.083e-09 0.0007 4.086e-09 0 4.14e-09 0 4.143e-09 0.0007 4.146e-09 0 4.2e-09 0 4.203e-09 0.0007 4.206e-09 0 4.26e-09 0 4.263e-09 0.0007 4.266e-09 0 4.32e-09 0 4.323e-09 0.0007 4.326e-09 0 4.38e-09 0 4.383e-09 0.0007 4.386e-09 0 4.44e-09 0 4.443e-09 0.0007 4.446e-09 0 4.5e-09 0 4.503e-09 0.0007 4.506e-09 0 4.56e-09 0 4.563e-09 0.0007 4.566e-09 0 4.62e-09 0 4.623e-09 0.0007 4.626e-09 0 4.68e-09 0 4.683e-09 0.0007 4.686e-09 0 4.74e-09 0 4.743e-09 0.0007 4.746e-09 0 4.8e-09 0 4.803e-09 0.0007 4.806e-09 0 4.86e-09 0 4.863e-09 0.0007 4.866e-09 0 4.92e-09 0 4.923e-09 0.0007 4.926e-09 0 4.98e-09 0 4.983e-09 0.0007 4.986e-09 0 5.04e-09 0 5.043e-09 0.0007 5.046e-09 0 5.1e-09 0 5.103e-09 0.0007 5.106e-09 0 5.16e-09 0 5.163e-09 0.0007 5.166e-09 0 5.22e-09 0 5.223e-09 0.0007 5.226e-09 0 5.28e-09 0 5.283e-09 0.0007 5.286e-09 0 5.34e-09 0 5.343e-09 0.0007 5.346e-09 0 5.4e-09 0 5.403e-09 0.0007 5.406e-09 0 5.46e-09 0 5.463e-09 0.0007 5.466e-09 0 5.52e-09 0 5.523e-09 0.0007 5.526e-09 0 5.58e-09 0 5.583e-09 0.0007 5.586e-09 0 5.64e-09 0 5.643e-09 0.0007 5.646e-09 0 5.7e-09 0 5.703e-09 0.0007 5.706e-09 0 5.76e-09 0 5.763e-09 0.0007 5.766e-09 0 5.82e-09 0 5.823e-09 0.0007 5.826e-09 0 5.88e-09 0 5.883e-09 0.0007 5.886e-09 0 5.94e-09 0 5.943e-09 0.0007 5.946e-09 0 6e-09 0 6.003e-09 0.0007 6.006e-09 0 6.06e-09 0 6.063e-09 0.0007 6.066e-09 0 6.12e-09 0 6.123e-09 0.0007 6.126e-09 0 6.18e-09 0 6.183e-09 0.0007 6.186e-09 0 6.24e-09 0 6.243e-09 0.0007 6.246e-09 0 6.3e-09 0 6.303e-09 0.0007 6.306e-09 0 6.36e-09 0 6.363e-09 0.0007 6.366e-09 0 6.42e-09 0 6.423e-09 0.0007 6.426e-09 0 6.48e-09 0 6.483e-09 0.0007 6.486e-09 0 6.54e-09 0 6.543e-09 0.0007 6.546e-09 0 6.6e-09 0 6.603e-09 0.0007 6.606e-09 0 6.66e-09 0 6.663e-09 0.0007 6.666e-09 0 6.72e-09 0 6.723e-09 0.0007 6.726e-09 0 6.78e-09 0 6.783e-09 0.0007 6.786e-09 0 6.84e-09 0 6.843e-09 0.0007 6.846e-09 0 6.9e-09 0 6.903e-09 0.0007 6.906e-09 0 6.96e-09 0 6.963e-09 0.0007 6.966e-09 0 7.02e-09 0 7.023e-09 0.0007 7.026e-09 0 7.08e-09 0 7.083e-09 0.0007 7.086e-09 0 7.14e-09 0 7.143e-09 0.0007 7.146e-09 0 7.2e-09 0 7.203e-09 0.0007 7.206e-09 0 7.26e-09 0 7.263e-09 0.0007 7.266e-09 0 7.32e-09 0 7.323e-09 0.0007 7.326e-09 0 7.38e-09 0 7.383e-09 0.0007 7.386e-09 0 7.44e-09 0 7.443e-09 0.0007 7.446e-09 0 7.5e-09 0 7.503e-09 0.0007 7.506e-09 0 7.56e-09 0 7.563e-09 0.0007 7.566e-09 0 7.62e-09 0 7.623e-09 0.0007 7.626e-09 0 7.68e-09 0 7.683e-09 0.0007 7.686e-09 0 7.74e-09 0 7.743e-09 0.0007 7.746e-09 0 7.8e-09 0 7.803e-09 0.0007 7.806e-09 0 7.86e-09 0 7.863e-09 0.0007 7.866e-09 0 7.92e-09 0 7.923e-09 0.0007 7.926e-09 0 7.98e-09 0 7.983e-09 0.0007 7.986e-09 0 8.04e-09 0 8.043e-09 0.0007 8.046e-09 0 8.1e-09 0 8.103e-09 0.0007 8.106e-09 0 8.16e-09 0 8.163e-09 0.0007 8.166e-09 0 8.22e-09 0 8.223e-09 0.0007 8.226e-09 0 8.28e-09 0 8.283e-09 0.0007 8.286e-09 0 8.34e-09 0 8.343e-09 0.0007 8.346e-09 0 8.4e-09 0 8.403e-09 0.0007 8.406e-09 0 8.46e-09 0 8.463e-09 0.0007 8.466e-09 0 8.52e-09 0 8.523e-09 0.0007 8.526e-09 0 8.58e-09 0 8.583e-09 0.0007 8.586e-09 0 8.64e-09 0 8.643e-09 0.0007 8.646e-09 0 8.7e-09 0 8.703e-09 0.0007 8.706e-09 0 8.76e-09 0 8.763e-09 0.0007 8.766e-09 0 8.82e-09 0 8.823e-09 0.0007 8.826e-09 0 8.88e-09 0 8.883e-09 0.0007 8.886e-09 0 8.94e-09 0 8.943e-09 0.0007 8.946e-09 0 9e-09 0 9.003e-09 0.0007 9.006e-09 0 9.06e-09 0 9.063e-09 0.0007 9.066e-09 0 9.12e-09 0 9.123e-09 0.0007 9.126e-09 0 9.18e-09 0 9.183e-09 0.0007 9.186e-09 0 9.24e-09 0 9.243e-09 0.0007 9.246e-09 0 9.3e-09 0 9.303e-09 0.0007 9.306e-09 0 9.36e-09 0 9.363e-09 0.0007 9.366e-09 0 9.42e-09 0 9.423e-09 0.0007 9.426e-09 0 9.48e-09 0 9.483e-09 0.0007 9.486e-09 0 9.54e-09 0 9.543e-09 0.0007 9.546e-09 0 9.6e-09 0 9.603e-09 0.0007 9.606e-09 0 9.66e-09 0 9.663e-09 0.0007 9.666e-09 0 9.72e-09 0 9.723e-09 0.0007 9.726e-09 0 9.78e-09 0 9.783e-09 0.0007 9.786e-09 0 9.84e-09 0 9.843e-09 0.0007 9.846e-09 0 9.9e-09 0 9.903e-09 0.0007 9.906e-09 0 9.96e-09 0 9.963e-09 0.0007 9.966e-09 0 1.002e-08 0 1.0023e-08 0.0007 1.0026e-08 0 1.008e-08 0 1.0083e-08 0.0007 1.0086e-08 0 1.014e-08 0 1.0143e-08 0.0007 1.0146e-08 0 1.02e-08 0 1.0203e-08 0.0007 1.0206e-08 0 1.026e-08 0 1.0263e-08 0.0007 1.0266e-08 0 1.032e-08 0 1.0323e-08 0.0007 1.0326e-08 0 1.038e-08 0 1.0383e-08 0.0007 1.0386e-08 0 1.044e-08 0 1.0443e-08 0.0007 1.0446e-08 0 1.05e-08 0 1.0503e-08 0.0007 1.0506e-08 0 1.056e-08 0 1.0563e-08 0.0007 1.0566e-08 0 1.062e-08 0 1.0623e-08 0.0007 1.0626e-08 0 1.068e-08 0 1.0683e-08 0.0007 1.0686e-08 0 1.074e-08 0 1.0743e-08 0.0007 1.0746e-08 0 1.08e-08 0 1.0803e-08 0.0007 1.0806e-08 0 1.086e-08 0 1.0863e-08 0.0007 1.0866e-08 0 1.092e-08 0 1.0923e-08 0.0007 1.0926e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.104e-08 0 1.1043e-08 0.0007 1.1046e-08 0 1.11e-08 0 1.1103e-08 0.0007 1.1106e-08 0 1.116e-08 0 1.1163e-08 0.0007 1.1166e-08 0 1.122e-08 0 1.1223e-08 0.0007 1.1226e-08 0 1.128e-08 0 1.1283e-08 0.0007 1.1286e-08 0 1.134e-08 0 1.1343e-08 0.0007 1.1346e-08 0 1.14e-08 0 1.1403e-08 0.0007 1.1406e-08 0 1.146e-08 0 1.1463e-08 0.0007 1.1466e-08 0 1.152e-08 0 1.1523e-08 0.0007 1.1526e-08 0 1.158e-08 0 1.1583e-08 0.0007 1.1586e-08 0 1.164e-08 0 1.1643e-08 0.0007 1.1646e-08 0 1.17e-08 0 1.1703e-08 0.0007 1.1706e-08 0 1.176e-08 0 1.1763e-08 0.0007 1.1766e-08 0 1.182e-08 0 1.1823e-08 0.0007 1.1826e-08 0 1.188e-08 0 1.1883e-08 0.0007 1.1886e-08 0 1.194e-08 0 1.1943e-08 0.0007 1.1946e-08 0 1.2e-08 0 1.2003e-08 0.0007 1.2006e-08 0 1.206e-08 0 1.2063e-08 0.0007 1.2066e-08 0 1.212e-08 0 1.2123e-08 0.0007 1.2126e-08 0 1.218e-08 0 1.2183e-08 0.0007 1.2186e-08 0 1.224e-08 0 1.2243e-08 0.0007 1.2246e-08 0 1.23e-08 0 1.2303e-08 0.0007 1.2306e-08 0 1.236e-08 0 1.2363e-08 0.0007 1.2366e-08 0 1.242e-08 0 1.2423e-08 0.0007 1.2426e-08 0 1.248e-08 0 1.2483e-08 0.0007 1.2486e-08 0 1.254e-08 0 1.2543e-08 0.0007 1.2546e-08 0 1.26e-08 0 1.2603e-08 0.0007 1.2606e-08 0 1.266e-08 0 1.2663e-08 0.0007 1.2666e-08 0 1.272e-08 0 1.2723e-08 0.0007 1.2726e-08 0 1.278e-08 0 1.2783e-08 0.0007 1.2786e-08 0 1.284e-08 0 1.2843e-08 0.0007 1.2846e-08 0 1.29e-08 0 1.2903e-08 0.0007 1.2906e-08 0 1.296e-08 0 1.2963e-08 0.0007 1.2966e-08 0 1.302e-08 0 1.3023e-08 0.0007 1.3026e-08 0 1.308e-08 0 1.3083e-08 0.0007 1.3086e-08 0 1.314e-08 0 1.3143e-08 0.0007 1.3146e-08 0 1.32e-08 0 1.3203e-08 0.0007 1.3206e-08 0 1.326e-08 0 1.3263e-08 0.0007 1.3266e-08 0 1.332e-08 0 1.3323e-08 0.0007 1.3326e-08 0 1.338e-08 0 1.3383e-08 0.0007 1.3386e-08 0 1.344e-08 0 1.3443e-08 0.0007 1.3446e-08 0 1.35e-08 0 1.3503e-08 0.0007 1.3506e-08 0 1.356e-08 0 1.3563e-08 0.0007 1.3566e-08 0 1.362e-08 0 1.3623e-08 0.0007 1.3626e-08 0 1.368e-08 0 1.3683e-08 0.0007 1.3686e-08 0 1.374e-08 0 1.3743e-08 0.0007 1.3746e-08 0 1.38e-08 0 1.3803e-08 0.0007 1.3806e-08 0 1.386e-08 0 1.3863e-08 0.0007 1.3866e-08 0 1.392e-08 0 1.3923e-08 0.0007 1.3926e-08 0 1.398e-08 0 1.3983e-08 0.0007 1.3986e-08 0 1.404e-08 0 1.4043e-08 0.0007 1.4046e-08 0 1.41e-08 0 1.4103e-08 0.0007 1.4106e-08 0 1.416e-08 0 1.4163e-08 0.0007 1.4166e-08 0 1.422e-08 0 1.4223e-08 0.0007 1.4226e-08 0 1.428e-08 0 1.4283e-08 0.0007 1.4286e-08 0 1.434e-08 0 1.4343e-08 0.0007 1.4346e-08 0 1.44e-08 0 1.4403e-08 0.0007 1.4406e-08 0 1.446e-08 0 1.4463e-08 0.0007 1.4466e-08 0 1.452e-08 0 1.4523e-08 0.0007 1.4526e-08 0 1.458e-08 0 1.4583e-08 0.0007 1.4586e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.47e-08 0 1.4703e-08 0.0007 1.4706e-08 0 1.476e-08 0 1.4763e-08 0.0007 1.4766e-08 0 1.482e-08 0 1.4823e-08 0.0007 1.4826e-08 0 1.488e-08 0 1.4883e-08 0.0007 1.4886e-08 0 1.494e-08 0 1.4943e-08 0.0007 1.4946e-08 0 1.5e-08 0 1.5003e-08 0.0007 1.5006e-08 0 1.506e-08 0 1.5063e-08 0.0007 1.5066e-08 0 1.512e-08 0 1.5123e-08 0.0007 1.5126e-08 0 1.518e-08 0 1.5183e-08 0.0007 1.5186e-08 0 1.524e-08 0 1.5243e-08 0.0007 1.5246e-08 0 1.53e-08 0 1.5303e-08 0.0007 1.5306e-08 0 1.536e-08 0 1.5363e-08 0.0007 1.5366e-08 0 1.542e-08 0 1.5423e-08 0.0007 1.5426e-08 0 1.548e-08 0 1.5483e-08 0.0007 1.5486e-08 0 1.554e-08 0 1.5543e-08 0.0007 1.5546e-08 0 1.56e-08 0 1.5603e-08 0.0007 1.5606e-08 0 1.566e-08 0 1.5663e-08 0.0007 1.5666e-08 0 1.572e-08 0 1.5723e-08 0.0007 1.5726e-08 0 1.578e-08 0 1.5783e-08 0.0007 1.5786e-08 0 1.584e-08 0 1.5843e-08 0.0007 1.5846e-08 0 1.59e-08 0 1.5903e-08 0.0007 1.5906e-08 0 1.596e-08 0 1.5963e-08 0.0007 1.5966e-08 0 1.602e-08 0 1.6023e-08 0.0007 1.6026e-08 0 1.608e-08 0 1.6083e-08 0.0007 1.6086e-08 0 1.614e-08 0 1.6143e-08 0.0007 1.6146e-08 0 1.62e-08 0 1.6203e-08 0.0007 1.6206e-08 0 1.626e-08 0 1.6263e-08 0.0007 1.6266e-08 0 1.632e-08 0 1.6323e-08 0.0007 1.6326e-08 0 1.638e-08 0 1.6383e-08 0.0007 1.6386e-08 0 1.644e-08 0 1.6443e-08 0.0007 1.6446e-08 0 1.65e-08 0 1.6503e-08 0.0007 1.6506e-08 0 1.656e-08 0 1.6563e-08 0.0007 1.6566e-08 0 1.662e-08 0 1.6623e-08 0.0007 1.6626e-08 0 1.668e-08 0 1.6683e-08 0.0007 1.6686e-08 0 1.674e-08 0 1.6743e-08 0.0007 1.6746e-08 0 1.68e-08 0 1.6803e-08 0.0007 1.6806e-08 0 1.686e-08 0 1.6863e-08 0.0007 1.6866e-08 0 1.692e-08 0 1.6923e-08 0.0007 1.6926e-08 0 1.698e-08 0 1.6983e-08 0.0007 1.6986e-08 0 1.704e-08 0 1.7043e-08 0.0007 1.7046e-08 0 1.71e-08 0 1.7103e-08 0.0007 1.7106e-08 0 1.716e-08 0 1.7163e-08 0.0007 1.7166e-08 0 1.722e-08 0 1.7223e-08 0.0007 1.7226e-08 0 1.728e-08 0 1.7283e-08 0.0007 1.7286e-08 0 1.734e-08 0 1.7343e-08 0.0007 1.7346e-08 0 1.74e-08 0 1.7403e-08 0.0007 1.7406e-08 0 1.746e-08 0 1.7463e-08 0.0007 1.7466e-08 0 1.752e-08 0 1.7523e-08 0.0007 1.7526e-08 0 1.758e-08 0 1.7583e-08 0.0007 1.7586e-08 0 1.764e-08 0 1.7643e-08 0.0007 1.7646e-08 0 1.77e-08 0 1.7703e-08 0.0007 1.7706e-08 0 1.776e-08 0 1.7763e-08 0.0007 1.7766e-08 0 1.782e-08 0 1.7823e-08 0.0007 1.7826e-08 0 1.788e-08 0 1.7883e-08 0.0007 1.7886e-08 0 1.794e-08 0 1.7943e-08 0.0007 1.7946e-08 0 1.8e-08 0 1.8003e-08 0.0007 1.8006e-08 0 1.806e-08 0 1.8063e-08 0.0007 1.8066e-08 0 1.812e-08 0 1.8123e-08 0.0007 1.8126e-08 0 1.818e-08 0 1.8183e-08 0.0007 1.8186e-08 0 1.824e-08 0 1.8243e-08 0.0007 1.8246e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.836e-08 0 1.8363e-08 0.0007 1.8366e-08 0 1.842e-08 0 1.8423e-08 0.0007 1.8426e-08 0 1.848e-08 0 1.8483e-08 0.0007 1.8486e-08 0 1.854e-08 0 1.8543e-08 0.0007 1.8546e-08 0 1.86e-08 0 1.8603e-08 0.0007 1.8606e-08 0 1.866e-08 0 1.8663e-08 0.0007 1.8666e-08 0 1.872e-08 0 1.8723e-08 0.0007 1.8726e-08 0 1.878e-08 0 1.8783e-08 0.0007 1.8786e-08 0 1.884e-08 0 1.8843e-08 0.0007 1.8846e-08 0 1.89e-08 0 1.8903e-08 0.0007 1.8906e-08 0 1.896e-08 0 1.8963e-08 0.0007 1.8966e-08 0 1.902e-08 0 1.9023e-08 0.0007 1.9026e-08 0 1.908e-08 0 1.9083e-08 0.0007 1.9086e-08 0 1.914e-08 0 1.9143e-08 0.0007 1.9146e-08 0 1.92e-08 0 1.9203e-08 0.0007 1.9206e-08 0 1.926e-08 0 1.9263e-08 0.0007 1.9266e-08 0 1.932e-08 0 1.9323e-08 0.0007 1.9326e-08 0 1.938e-08 0 1.9383e-08 0.0007 1.9386e-08 0 1.944e-08 0 1.9443e-08 0.0007 1.9446e-08 0 1.95e-08 0 1.9503e-08 0.0007 1.9506e-08 0 1.956e-08 0 1.9563e-08 0.0007 1.9566e-08 0 1.962e-08 0 1.9623e-08 0.0007 1.9626e-08 0 1.968e-08 0 1.9683e-08 0.0007 1.9686e-08 0 1.974e-08 0 1.9743e-08 0.0007 1.9746e-08 0 1.98e-08 0 1.9803e-08 0.0007 1.9806e-08 0 1.986e-08 0 1.9863e-08 0.0007 1.9866e-08 0 1.992e-08 0 1.9923e-08 0.0007 1.9926e-08 0 1.998e-08 0 1.9983e-08 0.0007 1.9986e-08 0 2.004e-08 0 2.0043e-08 0.0007 2.0046e-08 0 2.01e-08 0 2.0103e-08 0.0007 2.0106e-08 0 2.016e-08 0 2.0163e-08 0.0007 2.0166e-08 0 2.022e-08 0 2.0223e-08 0.0007 2.0226e-08 0 2.028e-08 0 2.0283e-08 0.0007 2.0286e-08 0 2.034e-08 0 2.0343e-08 0.0007 2.0346e-08 0 2.04e-08 0 2.0403e-08 0.0007 2.0406e-08 0 2.046e-08 0 2.0463e-08 0.0007 2.0466e-08 0 2.052e-08 0 2.0523e-08 0.0007 2.0526e-08 0 2.058e-08 0 2.0583e-08 0.0007 2.0586e-08 0 2.064e-08 0 2.0643e-08 0.0007 2.0646e-08 0 2.07e-08 0 2.0703e-08 0.0007 2.0706e-08 0 2.076e-08 0 2.0763e-08 0.0007 2.0766e-08 0 2.082e-08 0 2.0823e-08 0.0007 2.0826e-08 0 2.088e-08 0 2.0883e-08 0.0007 2.0886e-08 0 2.094e-08 0 2.0943e-08 0.0007 2.0946e-08 0 2.1e-08 0 2.1003e-08 0.0007 2.1006e-08 0 2.106e-08 0 2.1063e-08 0.0007 2.1066e-08 0 2.112e-08 0 2.1123e-08 0.0007 2.1126e-08 0 2.118e-08 0 2.1183e-08 0.0007 2.1186e-08 0 2.124e-08 0 2.1243e-08 0.0007 2.1246e-08 0 2.13e-08 0 2.1303e-08 0.0007 2.1306e-08 0 2.136e-08 0 2.1363e-08 0.0007 2.1366e-08 0 2.142e-08 0 2.1423e-08 0.0007 2.1426e-08 0 2.148e-08 0 2.1483e-08 0.0007 2.1486e-08 0 2.154e-08 0 2.1543e-08 0.0007 2.1546e-08 0 2.16e-08 0 2.1603e-08 0.0007 2.1606e-08 0 2.166e-08 0 2.1663e-08 0.0007 2.1666e-08 0 2.172e-08 0 2.1723e-08 0.0007 2.1726e-08 0 2.178e-08 0 2.1783e-08 0.0007 2.1786e-08 0 2.184e-08 0 2.1843e-08 0.0007 2.1846e-08 0 2.19e-08 0 2.1903e-08 0.0007 2.1906e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.202e-08 0 2.2023e-08 0.0007 2.2026e-08 0 2.208e-08 0 2.2083e-08 0.0007 2.2086e-08 0 2.214e-08 0 2.2143e-08 0.0007 2.2146e-08 0 2.22e-08 0 2.2203e-08 0.0007 2.2206e-08 0 2.226e-08 0 2.2263e-08 0.0007 2.2266e-08 0 2.232e-08 0 2.2323e-08 0.0007 2.2326e-08 0 2.238e-08 0 2.2383e-08 0.0007 2.2386e-08 0 2.244e-08 0 2.2443e-08 0.0007 2.2446e-08 0 2.25e-08 0 2.2503e-08 0.0007 2.2506e-08 0 2.256e-08 0 2.2563e-08 0.0007 2.2566e-08 0 2.262e-08 0 2.2623e-08 0.0007 2.2626e-08 0 2.268e-08 0 2.2683e-08 0.0007 2.2686e-08 0 2.274e-08 0 2.2743e-08 0.0007 2.2746e-08 0 2.28e-08 0 2.2803e-08 0.0007 2.2806e-08 0 2.286e-08 0 2.2863e-08 0.0007 2.2866e-08 0 2.292e-08 0 2.2923e-08 0.0007 2.2926e-08 0 2.298e-08 0 2.2983e-08 0.0007 2.2986e-08 0 2.304e-08 0 2.3043e-08 0.0007 2.3046e-08 0 2.31e-08 0 2.3103e-08 0.0007 2.3106e-08 0 2.316e-08 0 2.3163e-08 0.0007 2.3166e-08 0 2.322e-08 0 2.3223e-08 0.0007 2.3226e-08 0 2.328e-08 0 2.3283e-08 0.0007 2.3286e-08 0 2.334e-08 0 2.3343e-08 0.0007 2.3346e-08 0 2.34e-08 0 2.3403e-08 0.0007 2.3406e-08 0 2.346e-08 0 2.3463e-08 0.0007 2.3466e-08 0 2.352e-08 0 2.3523e-08 0.0007 2.3526e-08 0 2.358e-08 0 2.3583e-08 0.0007 2.3586e-08 0 2.364e-08 0 2.3643e-08 0.0007 2.3646e-08 0 2.37e-08 0 2.3703e-08 0.0007 2.3706e-08 0 2.376e-08 0 2.3763e-08 0.0007 2.3766e-08 0 2.382e-08 0 2.3823e-08 0.0007 2.3826e-08 0 2.388e-08 0 2.3883e-08 0.0007 2.3886e-08 0)
L_S2|A1 G1_2_RX _S2|A1  2.067833848e-12
L_S2|A2 _S2|A1 _S2|A2  4.135667696e-12
L_S2|A3 _S2|A3 _S2|AB  8.271335392e-12
L_S2|B1 IP2_2_OUT_RX _S2|B1  2.067833848e-12
L_S2|B2 _S2|B1 _S2|B2  4.135667696e-12
L_S2|B3 _S2|B3 _S2|AB  8.271335392e-12
L_S2|T1 T14 _S2|T1  2.067833848e-12
L_S2|T2 _S2|T1 _S2|T2  4.135667696e-12
L_S2|Q2 _S2|ABTQ _S2|Q1  4.135667696e-12
L_S2|Q1 _S2|Q1 S2  2.067833848e-12
IT15|T 0 T15  PWL(0 0 0 0 3e-12 0.0007 6e-12 0 6e-11 0 6.3e-11 0.0007 6.6e-11 0 1.2e-10 0 1.23e-10 0.0007 1.26e-10 0 1.8e-10 0 1.83e-10 0.0007 1.86e-10 0 2.4e-10 0 2.43e-10 0.0007 2.46e-10 0 3e-10 0 3.03e-10 0.0007 3.06e-10 0 3.6e-10 0 3.63e-10 0.0007 3.66e-10 0 4.2e-10 0 4.23e-10 0.0007 4.26e-10 0 4.8e-10 0 4.83e-10 0.0007 4.86e-10 0 5.4e-10 0 5.43e-10 0.0007 5.46e-10 0 6e-10 0 6.03e-10 0.0007 6.06e-10 0 6.6e-10 0 6.63e-10 0.0007 6.66e-10 0 7.2e-10 0 7.23e-10 0.0007 7.26e-10 0 7.8e-10 0 7.83e-10 0.0007 7.86e-10 0 8.4e-10 0 8.43e-10 0.0007 8.46e-10 0 9e-10 0 9.03e-10 0.0007 9.06e-10 0 9.6e-10 0 9.63e-10 0.0007 9.66e-10 0 1.02e-09 0 1.023e-09 0.0007 1.026e-09 0 1.08e-09 0 1.083e-09 0.0007 1.086e-09 0 1.14e-09 0 1.143e-09 0.0007 1.146e-09 0 1.2e-09 0 1.203e-09 0.0007 1.206e-09 0 1.26e-09 0 1.263e-09 0.0007 1.266e-09 0 1.32e-09 0 1.323e-09 0.0007 1.326e-09 0 1.38e-09 0 1.383e-09 0.0007 1.386e-09 0 1.44e-09 0 1.443e-09 0.0007 1.446e-09 0 1.5e-09 0 1.503e-09 0.0007 1.506e-09 0 1.56e-09 0 1.563e-09 0.0007 1.566e-09 0 1.62e-09 0 1.623e-09 0.0007 1.626e-09 0 1.68e-09 0 1.683e-09 0.0007 1.686e-09 0 1.74e-09 0 1.743e-09 0.0007 1.746e-09 0 1.8e-09 0 1.803e-09 0.0007 1.806e-09 0 1.86e-09 0 1.863e-09 0.0007 1.866e-09 0 1.92e-09 0 1.923e-09 0.0007 1.926e-09 0 1.98e-09 0 1.983e-09 0.0007 1.986e-09 0 2.04e-09 0 2.043e-09 0.0007 2.046e-09 0 2.1e-09 0 2.103e-09 0.0007 2.106e-09 0 2.16e-09 0 2.163e-09 0.0007 2.166e-09 0 2.22e-09 0 2.223e-09 0.0007 2.226e-09 0 2.28e-09 0 2.283e-09 0.0007 2.286e-09 0 2.34e-09 0 2.343e-09 0.0007 2.346e-09 0 2.4e-09 0 2.403e-09 0.0007 2.406e-09 0 2.46e-09 0 2.463e-09 0.0007 2.466e-09 0 2.52e-09 0 2.523e-09 0.0007 2.526e-09 0 2.58e-09 0 2.583e-09 0.0007 2.586e-09 0 2.64e-09 0 2.643e-09 0.0007 2.646e-09 0 2.7e-09 0 2.703e-09 0.0007 2.706e-09 0 2.76e-09 0 2.763e-09 0.0007 2.766e-09 0 2.82e-09 0 2.823e-09 0.0007 2.826e-09 0 2.88e-09 0 2.883e-09 0.0007 2.886e-09 0 2.94e-09 0 2.943e-09 0.0007 2.946e-09 0 3e-09 0 3.003e-09 0.0007 3.006e-09 0 3.06e-09 0 3.063e-09 0.0007 3.066e-09 0 3.12e-09 0 3.123e-09 0.0007 3.126e-09 0 3.18e-09 0 3.183e-09 0.0007 3.186e-09 0 3.24e-09 0 3.243e-09 0.0007 3.246e-09 0 3.3e-09 0 3.303e-09 0.0007 3.306e-09 0 3.36e-09 0 3.363e-09 0.0007 3.366e-09 0 3.42e-09 0 3.423e-09 0.0007 3.426e-09 0 3.48e-09 0 3.483e-09 0.0007 3.486e-09 0 3.54e-09 0 3.543e-09 0.0007 3.546e-09 0 3.6e-09 0 3.603e-09 0.0007 3.606e-09 0 3.66e-09 0 3.663e-09 0.0007 3.666e-09 0 3.72e-09 0 3.723e-09 0.0007 3.726e-09 0 3.78e-09 0 3.783e-09 0.0007 3.786e-09 0 3.84e-09 0 3.843e-09 0.0007 3.846e-09 0 3.9e-09 0 3.903e-09 0.0007 3.906e-09 0 3.96e-09 0 3.963e-09 0.0007 3.966e-09 0 4.02e-09 0 4.023e-09 0.0007 4.026e-09 0 4.08e-09 0 4.083e-09 0.0007 4.086e-09 0 4.14e-09 0 4.143e-09 0.0007 4.146e-09 0 4.2e-09 0 4.203e-09 0.0007 4.206e-09 0 4.26e-09 0 4.263e-09 0.0007 4.266e-09 0 4.32e-09 0 4.323e-09 0.0007 4.326e-09 0 4.38e-09 0 4.383e-09 0.0007 4.386e-09 0 4.44e-09 0 4.443e-09 0.0007 4.446e-09 0 4.5e-09 0 4.503e-09 0.0007 4.506e-09 0 4.56e-09 0 4.563e-09 0.0007 4.566e-09 0 4.62e-09 0 4.623e-09 0.0007 4.626e-09 0 4.68e-09 0 4.683e-09 0.0007 4.686e-09 0 4.74e-09 0 4.743e-09 0.0007 4.746e-09 0 4.8e-09 0 4.803e-09 0.0007 4.806e-09 0 4.86e-09 0 4.863e-09 0.0007 4.866e-09 0 4.92e-09 0 4.923e-09 0.0007 4.926e-09 0 4.98e-09 0 4.983e-09 0.0007 4.986e-09 0 5.04e-09 0 5.043e-09 0.0007 5.046e-09 0 5.1e-09 0 5.103e-09 0.0007 5.106e-09 0 5.16e-09 0 5.163e-09 0.0007 5.166e-09 0 5.22e-09 0 5.223e-09 0.0007 5.226e-09 0 5.28e-09 0 5.283e-09 0.0007 5.286e-09 0 5.34e-09 0 5.343e-09 0.0007 5.346e-09 0 5.4e-09 0 5.403e-09 0.0007 5.406e-09 0 5.46e-09 0 5.463e-09 0.0007 5.466e-09 0 5.52e-09 0 5.523e-09 0.0007 5.526e-09 0 5.58e-09 0 5.583e-09 0.0007 5.586e-09 0 5.64e-09 0 5.643e-09 0.0007 5.646e-09 0 5.7e-09 0 5.703e-09 0.0007 5.706e-09 0 5.76e-09 0 5.763e-09 0.0007 5.766e-09 0 5.82e-09 0 5.823e-09 0.0007 5.826e-09 0 5.88e-09 0 5.883e-09 0.0007 5.886e-09 0 5.94e-09 0 5.943e-09 0.0007 5.946e-09 0 6e-09 0 6.003e-09 0.0007 6.006e-09 0 6.06e-09 0 6.063e-09 0.0007 6.066e-09 0 6.12e-09 0 6.123e-09 0.0007 6.126e-09 0 6.18e-09 0 6.183e-09 0.0007 6.186e-09 0 6.24e-09 0 6.243e-09 0.0007 6.246e-09 0 6.3e-09 0 6.303e-09 0.0007 6.306e-09 0 6.36e-09 0 6.363e-09 0.0007 6.366e-09 0 6.42e-09 0 6.423e-09 0.0007 6.426e-09 0 6.48e-09 0 6.483e-09 0.0007 6.486e-09 0 6.54e-09 0 6.543e-09 0.0007 6.546e-09 0 6.6e-09 0 6.603e-09 0.0007 6.606e-09 0 6.66e-09 0 6.663e-09 0.0007 6.666e-09 0 6.72e-09 0 6.723e-09 0.0007 6.726e-09 0 6.78e-09 0 6.783e-09 0.0007 6.786e-09 0 6.84e-09 0 6.843e-09 0.0007 6.846e-09 0 6.9e-09 0 6.903e-09 0.0007 6.906e-09 0 6.96e-09 0 6.963e-09 0.0007 6.966e-09 0 7.02e-09 0 7.023e-09 0.0007 7.026e-09 0 7.08e-09 0 7.083e-09 0.0007 7.086e-09 0 7.14e-09 0 7.143e-09 0.0007 7.146e-09 0 7.2e-09 0 7.203e-09 0.0007 7.206e-09 0 7.26e-09 0 7.263e-09 0.0007 7.266e-09 0 7.32e-09 0 7.323e-09 0.0007 7.326e-09 0 7.38e-09 0 7.383e-09 0.0007 7.386e-09 0 7.44e-09 0 7.443e-09 0.0007 7.446e-09 0 7.5e-09 0 7.503e-09 0.0007 7.506e-09 0 7.56e-09 0 7.563e-09 0.0007 7.566e-09 0 7.62e-09 0 7.623e-09 0.0007 7.626e-09 0 7.68e-09 0 7.683e-09 0.0007 7.686e-09 0 7.74e-09 0 7.743e-09 0.0007 7.746e-09 0 7.8e-09 0 7.803e-09 0.0007 7.806e-09 0 7.86e-09 0 7.863e-09 0.0007 7.866e-09 0 7.92e-09 0 7.923e-09 0.0007 7.926e-09 0 7.98e-09 0 7.983e-09 0.0007 7.986e-09 0 8.04e-09 0 8.043e-09 0.0007 8.046e-09 0 8.1e-09 0 8.103e-09 0.0007 8.106e-09 0 8.16e-09 0 8.163e-09 0.0007 8.166e-09 0 8.22e-09 0 8.223e-09 0.0007 8.226e-09 0 8.28e-09 0 8.283e-09 0.0007 8.286e-09 0 8.34e-09 0 8.343e-09 0.0007 8.346e-09 0 8.4e-09 0 8.403e-09 0.0007 8.406e-09 0 8.46e-09 0 8.463e-09 0.0007 8.466e-09 0 8.52e-09 0 8.523e-09 0.0007 8.526e-09 0 8.58e-09 0 8.583e-09 0.0007 8.586e-09 0 8.64e-09 0 8.643e-09 0.0007 8.646e-09 0 8.7e-09 0 8.703e-09 0.0007 8.706e-09 0 8.76e-09 0 8.763e-09 0.0007 8.766e-09 0 8.82e-09 0 8.823e-09 0.0007 8.826e-09 0 8.88e-09 0 8.883e-09 0.0007 8.886e-09 0 8.94e-09 0 8.943e-09 0.0007 8.946e-09 0 9e-09 0 9.003e-09 0.0007 9.006e-09 0 9.06e-09 0 9.063e-09 0.0007 9.066e-09 0 9.12e-09 0 9.123e-09 0.0007 9.126e-09 0 9.18e-09 0 9.183e-09 0.0007 9.186e-09 0 9.24e-09 0 9.243e-09 0.0007 9.246e-09 0 9.3e-09 0 9.303e-09 0.0007 9.306e-09 0 9.36e-09 0 9.363e-09 0.0007 9.366e-09 0 9.42e-09 0 9.423e-09 0.0007 9.426e-09 0 9.48e-09 0 9.483e-09 0.0007 9.486e-09 0 9.54e-09 0 9.543e-09 0.0007 9.546e-09 0 9.6e-09 0 9.603e-09 0.0007 9.606e-09 0 9.66e-09 0 9.663e-09 0.0007 9.666e-09 0 9.72e-09 0 9.723e-09 0.0007 9.726e-09 0 9.78e-09 0 9.783e-09 0.0007 9.786e-09 0 9.84e-09 0 9.843e-09 0.0007 9.846e-09 0 9.9e-09 0 9.903e-09 0.0007 9.906e-09 0 9.96e-09 0 9.963e-09 0.0007 9.966e-09 0 1.002e-08 0 1.0023e-08 0.0007 1.0026e-08 0 1.008e-08 0 1.0083e-08 0.0007 1.0086e-08 0 1.014e-08 0 1.0143e-08 0.0007 1.0146e-08 0 1.02e-08 0 1.0203e-08 0.0007 1.0206e-08 0 1.026e-08 0 1.0263e-08 0.0007 1.0266e-08 0 1.032e-08 0 1.0323e-08 0.0007 1.0326e-08 0 1.038e-08 0 1.0383e-08 0.0007 1.0386e-08 0 1.044e-08 0 1.0443e-08 0.0007 1.0446e-08 0 1.05e-08 0 1.0503e-08 0.0007 1.0506e-08 0 1.056e-08 0 1.0563e-08 0.0007 1.0566e-08 0 1.062e-08 0 1.0623e-08 0.0007 1.0626e-08 0 1.068e-08 0 1.0683e-08 0.0007 1.0686e-08 0 1.074e-08 0 1.0743e-08 0.0007 1.0746e-08 0 1.08e-08 0 1.0803e-08 0.0007 1.0806e-08 0 1.086e-08 0 1.0863e-08 0.0007 1.0866e-08 0 1.092e-08 0 1.0923e-08 0.0007 1.0926e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.104e-08 0 1.1043e-08 0.0007 1.1046e-08 0 1.11e-08 0 1.1103e-08 0.0007 1.1106e-08 0 1.116e-08 0 1.1163e-08 0.0007 1.1166e-08 0 1.122e-08 0 1.1223e-08 0.0007 1.1226e-08 0 1.128e-08 0 1.1283e-08 0.0007 1.1286e-08 0 1.134e-08 0 1.1343e-08 0.0007 1.1346e-08 0 1.14e-08 0 1.1403e-08 0.0007 1.1406e-08 0 1.146e-08 0 1.1463e-08 0.0007 1.1466e-08 0 1.152e-08 0 1.1523e-08 0.0007 1.1526e-08 0 1.158e-08 0 1.1583e-08 0.0007 1.1586e-08 0 1.164e-08 0 1.1643e-08 0.0007 1.1646e-08 0 1.17e-08 0 1.1703e-08 0.0007 1.1706e-08 0 1.176e-08 0 1.1763e-08 0.0007 1.1766e-08 0 1.182e-08 0 1.1823e-08 0.0007 1.1826e-08 0 1.188e-08 0 1.1883e-08 0.0007 1.1886e-08 0 1.194e-08 0 1.1943e-08 0.0007 1.1946e-08 0 1.2e-08 0 1.2003e-08 0.0007 1.2006e-08 0 1.206e-08 0 1.2063e-08 0.0007 1.2066e-08 0 1.212e-08 0 1.2123e-08 0.0007 1.2126e-08 0 1.218e-08 0 1.2183e-08 0.0007 1.2186e-08 0 1.224e-08 0 1.2243e-08 0.0007 1.2246e-08 0 1.23e-08 0 1.2303e-08 0.0007 1.2306e-08 0 1.236e-08 0 1.2363e-08 0.0007 1.2366e-08 0 1.242e-08 0 1.2423e-08 0.0007 1.2426e-08 0 1.248e-08 0 1.2483e-08 0.0007 1.2486e-08 0 1.254e-08 0 1.2543e-08 0.0007 1.2546e-08 0 1.26e-08 0 1.2603e-08 0.0007 1.2606e-08 0 1.266e-08 0 1.2663e-08 0.0007 1.2666e-08 0 1.272e-08 0 1.2723e-08 0.0007 1.2726e-08 0 1.278e-08 0 1.2783e-08 0.0007 1.2786e-08 0 1.284e-08 0 1.2843e-08 0.0007 1.2846e-08 0 1.29e-08 0 1.2903e-08 0.0007 1.2906e-08 0 1.296e-08 0 1.2963e-08 0.0007 1.2966e-08 0 1.302e-08 0 1.3023e-08 0.0007 1.3026e-08 0 1.308e-08 0 1.3083e-08 0.0007 1.3086e-08 0 1.314e-08 0 1.3143e-08 0.0007 1.3146e-08 0 1.32e-08 0 1.3203e-08 0.0007 1.3206e-08 0 1.326e-08 0 1.3263e-08 0.0007 1.3266e-08 0 1.332e-08 0 1.3323e-08 0.0007 1.3326e-08 0 1.338e-08 0 1.3383e-08 0.0007 1.3386e-08 0 1.344e-08 0 1.3443e-08 0.0007 1.3446e-08 0 1.35e-08 0 1.3503e-08 0.0007 1.3506e-08 0 1.356e-08 0 1.3563e-08 0.0007 1.3566e-08 0 1.362e-08 0 1.3623e-08 0.0007 1.3626e-08 0 1.368e-08 0 1.3683e-08 0.0007 1.3686e-08 0 1.374e-08 0 1.3743e-08 0.0007 1.3746e-08 0 1.38e-08 0 1.3803e-08 0.0007 1.3806e-08 0 1.386e-08 0 1.3863e-08 0.0007 1.3866e-08 0 1.392e-08 0 1.3923e-08 0.0007 1.3926e-08 0 1.398e-08 0 1.3983e-08 0.0007 1.3986e-08 0 1.404e-08 0 1.4043e-08 0.0007 1.4046e-08 0 1.41e-08 0 1.4103e-08 0.0007 1.4106e-08 0 1.416e-08 0 1.4163e-08 0.0007 1.4166e-08 0 1.422e-08 0 1.4223e-08 0.0007 1.4226e-08 0 1.428e-08 0 1.4283e-08 0.0007 1.4286e-08 0 1.434e-08 0 1.4343e-08 0.0007 1.4346e-08 0 1.44e-08 0 1.4403e-08 0.0007 1.4406e-08 0 1.446e-08 0 1.4463e-08 0.0007 1.4466e-08 0 1.452e-08 0 1.4523e-08 0.0007 1.4526e-08 0 1.458e-08 0 1.4583e-08 0.0007 1.4586e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.47e-08 0 1.4703e-08 0.0007 1.4706e-08 0 1.476e-08 0 1.4763e-08 0.0007 1.4766e-08 0 1.482e-08 0 1.4823e-08 0.0007 1.4826e-08 0 1.488e-08 0 1.4883e-08 0.0007 1.4886e-08 0 1.494e-08 0 1.4943e-08 0.0007 1.4946e-08 0 1.5e-08 0 1.5003e-08 0.0007 1.5006e-08 0 1.506e-08 0 1.5063e-08 0.0007 1.5066e-08 0 1.512e-08 0 1.5123e-08 0.0007 1.5126e-08 0 1.518e-08 0 1.5183e-08 0.0007 1.5186e-08 0 1.524e-08 0 1.5243e-08 0.0007 1.5246e-08 0 1.53e-08 0 1.5303e-08 0.0007 1.5306e-08 0 1.536e-08 0 1.5363e-08 0.0007 1.5366e-08 0 1.542e-08 0 1.5423e-08 0.0007 1.5426e-08 0 1.548e-08 0 1.5483e-08 0.0007 1.5486e-08 0 1.554e-08 0 1.5543e-08 0.0007 1.5546e-08 0 1.56e-08 0 1.5603e-08 0.0007 1.5606e-08 0 1.566e-08 0 1.5663e-08 0.0007 1.5666e-08 0 1.572e-08 0 1.5723e-08 0.0007 1.5726e-08 0 1.578e-08 0 1.5783e-08 0.0007 1.5786e-08 0 1.584e-08 0 1.5843e-08 0.0007 1.5846e-08 0 1.59e-08 0 1.5903e-08 0.0007 1.5906e-08 0 1.596e-08 0 1.5963e-08 0.0007 1.5966e-08 0 1.602e-08 0 1.6023e-08 0.0007 1.6026e-08 0 1.608e-08 0 1.6083e-08 0.0007 1.6086e-08 0 1.614e-08 0 1.6143e-08 0.0007 1.6146e-08 0 1.62e-08 0 1.6203e-08 0.0007 1.6206e-08 0 1.626e-08 0 1.6263e-08 0.0007 1.6266e-08 0 1.632e-08 0 1.6323e-08 0.0007 1.6326e-08 0 1.638e-08 0 1.6383e-08 0.0007 1.6386e-08 0 1.644e-08 0 1.6443e-08 0.0007 1.6446e-08 0 1.65e-08 0 1.6503e-08 0.0007 1.6506e-08 0 1.656e-08 0 1.6563e-08 0.0007 1.6566e-08 0 1.662e-08 0 1.6623e-08 0.0007 1.6626e-08 0 1.668e-08 0 1.6683e-08 0.0007 1.6686e-08 0 1.674e-08 0 1.6743e-08 0.0007 1.6746e-08 0 1.68e-08 0 1.6803e-08 0.0007 1.6806e-08 0 1.686e-08 0 1.6863e-08 0.0007 1.6866e-08 0 1.692e-08 0 1.6923e-08 0.0007 1.6926e-08 0 1.698e-08 0 1.6983e-08 0.0007 1.6986e-08 0 1.704e-08 0 1.7043e-08 0.0007 1.7046e-08 0 1.71e-08 0 1.7103e-08 0.0007 1.7106e-08 0 1.716e-08 0 1.7163e-08 0.0007 1.7166e-08 0 1.722e-08 0 1.7223e-08 0.0007 1.7226e-08 0 1.728e-08 0 1.7283e-08 0.0007 1.7286e-08 0 1.734e-08 0 1.7343e-08 0.0007 1.7346e-08 0 1.74e-08 0 1.7403e-08 0.0007 1.7406e-08 0 1.746e-08 0 1.7463e-08 0.0007 1.7466e-08 0 1.752e-08 0 1.7523e-08 0.0007 1.7526e-08 0 1.758e-08 0 1.7583e-08 0.0007 1.7586e-08 0 1.764e-08 0 1.7643e-08 0.0007 1.7646e-08 0 1.77e-08 0 1.7703e-08 0.0007 1.7706e-08 0 1.776e-08 0 1.7763e-08 0.0007 1.7766e-08 0 1.782e-08 0 1.7823e-08 0.0007 1.7826e-08 0 1.788e-08 0 1.7883e-08 0.0007 1.7886e-08 0 1.794e-08 0 1.7943e-08 0.0007 1.7946e-08 0 1.8e-08 0 1.8003e-08 0.0007 1.8006e-08 0 1.806e-08 0 1.8063e-08 0.0007 1.8066e-08 0 1.812e-08 0 1.8123e-08 0.0007 1.8126e-08 0 1.818e-08 0 1.8183e-08 0.0007 1.8186e-08 0 1.824e-08 0 1.8243e-08 0.0007 1.8246e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.836e-08 0 1.8363e-08 0.0007 1.8366e-08 0 1.842e-08 0 1.8423e-08 0.0007 1.8426e-08 0 1.848e-08 0 1.8483e-08 0.0007 1.8486e-08 0 1.854e-08 0 1.8543e-08 0.0007 1.8546e-08 0 1.86e-08 0 1.8603e-08 0.0007 1.8606e-08 0 1.866e-08 0 1.8663e-08 0.0007 1.8666e-08 0 1.872e-08 0 1.8723e-08 0.0007 1.8726e-08 0 1.878e-08 0 1.8783e-08 0.0007 1.8786e-08 0 1.884e-08 0 1.8843e-08 0.0007 1.8846e-08 0 1.89e-08 0 1.8903e-08 0.0007 1.8906e-08 0 1.896e-08 0 1.8963e-08 0.0007 1.8966e-08 0 1.902e-08 0 1.9023e-08 0.0007 1.9026e-08 0 1.908e-08 0 1.9083e-08 0.0007 1.9086e-08 0 1.914e-08 0 1.9143e-08 0.0007 1.9146e-08 0 1.92e-08 0 1.9203e-08 0.0007 1.9206e-08 0 1.926e-08 0 1.9263e-08 0.0007 1.9266e-08 0 1.932e-08 0 1.9323e-08 0.0007 1.9326e-08 0 1.938e-08 0 1.9383e-08 0.0007 1.9386e-08 0 1.944e-08 0 1.9443e-08 0.0007 1.9446e-08 0 1.95e-08 0 1.9503e-08 0.0007 1.9506e-08 0 1.956e-08 0 1.9563e-08 0.0007 1.9566e-08 0 1.962e-08 0 1.9623e-08 0.0007 1.9626e-08 0 1.968e-08 0 1.9683e-08 0.0007 1.9686e-08 0 1.974e-08 0 1.9743e-08 0.0007 1.9746e-08 0 1.98e-08 0 1.9803e-08 0.0007 1.9806e-08 0 1.986e-08 0 1.9863e-08 0.0007 1.9866e-08 0 1.992e-08 0 1.9923e-08 0.0007 1.9926e-08 0 1.998e-08 0 1.9983e-08 0.0007 1.9986e-08 0 2.004e-08 0 2.0043e-08 0.0007 2.0046e-08 0 2.01e-08 0 2.0103e-08 0.0007 2.0106e-08 0 2.016e-08 0 2.0163e-08 0.0007 2.0166e-08 0 2.022e-08 0 2.0223e-08 0.0007 2.0226e-08 0 2.028e-08 0 2.0283e-08 0.0007 2.0286e-08 0 2.034e-08 0 2.0343e-08 0.0007 2.0346e-08 0 2.04e-08 0 2.0403e-08 0.0007 2.0406e-08 0 2.046e-08 0 2.0463e-08 0.0007 2.0466e-08 0 2.052e-08 0 2.0523e-08 0.0007 2.0526e-08 0 2.058e-08 0 2.0583e-08 0.0007 2.0586e-08 0 2.064e-08 0 2.0643e-08 0.0007 2.0646e-08 0 2.07e-08 0 2.0703e-08 0.0007 2.0706e-08 0 2.076e-08 0 2.0763e-08 0.0007 2.0766e-08 0 2.082e-08 0 2.0823e-08 0.0007 2.0826e-08 0 2.088e-08 0 2.0883e-08 0.0007 2.0886e-08 0 2.094e-08 0 2.0943e-08 0.0007 2.0946e-08 0 2.1e-08 0 2.1003e-08 0.0007 2.1006e-08 0 2.106e-08 0 2.1063e-08 0.0007 2.1066e-08 0 2.112e-08 0 2.1123e-08 0.0007 2.1126e-08 0 2.118e-08 0 2.1183e-08 0.0007 2.1186e-08 0 2.124e-08 0 2.1243e-08 0.0007 2.1246e-08 0 2.13e-08 0 2.1303e-08 0.0007 2.1306e-08 0 2.136e-08 0 2.1363e-08 0.0007 2.1366e-08 0 2.142e-08 0 2.1423e-08 0.0007 2.1426e-08 0 2.148e-08 0 2.1483e-08 0.0007 2.1486e-08 0 2.154e-08 0 2.1543e-08 0.0007 2.1546e-08 0 2.16e-08 0 2.1603e-08 0.0007 2.1606e-08 0 2.166e-08 0 2.1663e-08 0.0007 2.1666e-08 0 2.172e-08 0 2.1723e-08 0.0007 2.1726e-08 0 2.178e-08 0 2.1783e-08 0.0007 2.1786e-08 0 2.184e-08 0 2.1843e-08 0.0007 2.1846e-08 0 2.19e-08 0 2.1903e-08 0.0007 2.1906e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.202e-08 0 2.2023e-08 0.0007 2.2026e-08 0 2.208e-08 0 2.2083e-08 0.0007 2.2086e-08 0 2.214e-08 0 2.2143e-08 0.0007 2.2146e-08 0 2.22e-08 0 2.2203e-08 0.0007 2.2206e-08 0 2.226e-08 0 2.2263e-08 0.0007 2.2266e-08 0 2.232e-08 0 2.2323e-08 0.0007 2.2326e-08 0 2.238e-08 0 2.2383e-08 0.0007 2.2386e-08 0 2.244e-08 0 2.2443e-08 0.0007 2.2446e-08 0 2.25e-08 0 2.2503e-08 0.0007 2.2506e-08 0 2.256e-08 0 2.2563e-08 0.0007 2.2566e-08 0 2.262e-08 0 2.2623e-08 0.0007 2.2626e-08 0 2.268e-08 0 2.2683e-08 0.0007 2.2686e-08 0 2.274e-08 0 2.2743e-08 0.0007 2.2746e-08 0 2.28e-08 0 2.2803e-08 0.0007 2.2806e-08 0 2.286e-08 0 2.2863e-08 0.0007 2.2866e-08 0 2.292e-08 0 2.2923e-08 0.0007 2.2926e-08 0 2.298e-08 0 2.2983e-08 0.0007 2.2986e-08 0 2.304e-08 0 2.3043e-08 0.0007 2.3046e-08 0 2.31e-08 0 2.3103e-08 0.0007 2.3106e-08 0 2.316e-08 0 2.3163e-08 0.0007 2.3166e-08 0 2.322e-08 0 2.3223e-08 0.0007 2.3226e-08 0 2.328e-08 0 2.3283e-08 0.0007 2.3286e-08 0 2.334e-08 0 2.3343e-08 0.0007 2.3346e-08 0 2.34e-08 0 2.3403e-08 0.0007 2.3406e-08 0 2.346e-08 0 2.3463e-08 0.0007 2.3466e-08 0 2.352e-08 0 2.3523e-08 0.0007 2.3526e-08 0 2.358e-08 0 2.3583e-08 0.0007 2.3586e-08 0 2.364e-08 0 2.3643e-08 0.0007 2.3646e-08 0 2.37e-08 0 2.3703e-08 0.0007 2.3706e-08 0 2.376e-08 0 2.3763e-08 0.0007 2.3766e-08 0 2.382e-08 0 2.3823e-08 0.0007 2.3826e-08 0 2.388e-08 0 2.3883e-08 0.0007 2.3886e-08 0)
L_S3|A1 G2_2_RX _S3|A1  2.067833848e-12
L_S3|A2 _S3|A1 _S3|A2  4.135667696e-12
L_S3|A3 _S3|A3 _S3|AB  8.271335392e-12
L_S3|B1 IP3_2_OUT_RX _S3|B1  2.067833848e-12
L_S3|B2 _S3|B1 _S3|B2  4.135667696e-12
L_S3|B3 _S3|B3 _S3|AB  8.271335392e-12
L_S3|T1 T15 _S3|T1  2.067833848e-12
L_S3|T2 _S3|T1 _S3|T2  4.135667696e-12
L_S3|Q2 _S3|ABTQ _S3|Q1  4.135667696e-12
L_S3|Q1 _S3|Q1 S3  2.067833848e-12
IT16|T 0 T16  PWL(0 0 0 0 3e-12 0.0007 6e-12 0 6e-11 0 6.3e-11 0.0007 6.6e-11 0 1.2e-10 0 1.23e-10 0.0007 1.26e-10 0 1.8e-10 0 1.83e-10 0.0007 1.86e-10 0 2.4e-10 0 2.43e-10 0.0007 2.46e-10 0 3e-10 0 3.03e-10 0.0007 3.06e-10 0 3.6e-10 0 3.63e-10 0.0007 3.66e-10 0 4.2e-10 0 4.23e-10 0.0007 4.26e-10 0 4.8e-10 0 4.83e-10 0.0007 4.86e-10 0 5.4e-10 0 5.43e-10 0.0007 5.46e-10 0 6e-10 0 6.03e-10 0.0007 6.06e-10 0 6.6e-10 0 6.63e-10 0.0007 6.66e-10 0 7.2e-10 0 7.23e-10 0.0007 7.26e-10 0 7.8e-10 0 7.83e-10 0.0007 7.86e-10 0 8.4e-10 0 8.43e-10 0.0007 8.46e-10 0 9e-10 0 9.03e-10 0.0007 9.06e-10 0 9.6e-10 0 9.63e-10 0.0007 9.66e-10 0 1.02e-09 0 1.023e-09 0.0007 1.026e-09 0 1.08e-09 0 1.083e-09 0.0007 1.086e-09 0 1.14e-09 0 1.143e-09 0.0007 1.146e-09 0 1.2e-09 0 1.203e-09 0.0007 1.206e-09 0 1.26e-09 0 1.263e-09 0.0007 1.266e-09 0 1.32e-09 0 1.323e-09 0.0007 1.326e-09 0 1.38e-09 0 1.383e-09 0.0007 1.386e-09 0 1.44e-09 0 1.443e-09 0.0007 1.446e-09 0 1.5e-09 0 1.503e-09 0.0007 1.506e-09 0 1.56e-09 0 1.563e-09 0.0007 1.566e-09 0 1.62e-09 0 1.623e-09 0.0007 1.626e-09 0 1.68e-09 0 1.683e-09 0.0007 1.686e-09 0 1.74e-09 0 1.743e-09 0.0007 1.746e-09 0 1.8e-09 0 1.803e-09 0.0007 1.806e-09 0 1.86e-09 0 1.863e-09 0.0007 1.866e-09 0 1.92e-09 0 1.923e-09 0.0007 1.926e-09 0 1.98e-09 0 1.983e-09 0.0007 1.986e-09 0 2.04e-09 0 2.043e-09 0.0007 2.046e-09 0 2.1e-09 0 2.103e-09 0.0007 2.106e-09 0 2.16e-09 0 2.163e-09 0.0007 2.166e-09 0 2.22e-09 0 2.223e-09 0.0007 2.226e-09 0 2.28e-09 0 2.283e-09 0.0007 2.286e-09 0 2.34e-09 0 2.343e-09 0.0007 2.346e-09 0 2.4e-09 0 2.403e-09 0.0007 2.406e-09 0 2.46e-09 0 2.463e-09 0.0007 2.466e-09 0 2.52e-09 0 2.523e-09 0.0007 2.526e-09 0 2.58e-09 0 2.583e-09 0.0007 2.586e-09 0 2.64e-09 0 2.643e-09 0.0007 2.646e-09 0 2.7e-09 0 2.703e-09 0.0007 2.706e-09 0 2.76e-09 0 2.763e-09 0.0007 2.766e-09 0 2.82e-09 0 2.823e-09 0.0007 2.826e-09 0 2.88e-09 0 2.883e-09 0.0007 2.886e-09 0 2.94e-09 0 2.943e-09 0.0007 2.946e-09 0 3e-09 0 3.003e-09 0.0007 3.006e-09 0 3.06e-09 0 3.063e-09 0.0007 3.066e-09 0 3.12e-09 0 3.123e-09 0.0007 3.126e-09 0 3.18e-09 0 3.183e-09 0.0007 3.186e-09 0 3.24e-09 0 3.243e-09 0.0007 3.246e-09 0 3.3e-09 0 3.303e-09 0.0007 3.306e-09 0 3.36e-09 0 3.363e-09 0.0007 3.366e-09 0 3.42e-09 0 3.423e-09 0.0007 3.426e-09 0 3.48e-09 0 3.483e-09 0.0007 3.486e-09 0 3.54e-09 0 3.543e-09 0.0007 3.546e-09 0 3.6e-09 0 3.603e-09 0.0007 3.606e-09 0 3.66e-09 0 3.663e-09 0.0007 3.666e-09 0 3.72e-09 0 3.723e-09 0.0007 3.726e-09 0 3.78e-09 0 3.783e-09 0.0007 3.786e-09 0 3.84e-09 0 3.843e-09 0.0007 3.846e-09 0 3.9e-09 0 3.903e-09 0.0007 3.906e-09 0 3.96e-09 0 3.963e-09 0.0007 3.966e-09 0 4.02e-09 0 4.023e-09 0.0007 4.026e-09 0 4.08e-09 0 4.083e-09 0.0007 4.086e-09 0 4.14e-09 0 4.143e-09 0.0007 4.146e-09 0 4.2e-09 0 4.203e-09 0.0007 4.206e-09 0 4.26e-09 0 4.263e-09 0.0007 4.266e-09 0 4.32e-09 0 4.323e-09 0.0007 4.326e-09 0 4.38e-09 0 4.383e-09 0.0007 4.386e-09 0 4.44e-09 0 4.443e-09 0.0007 4.446e-09 0 4.5e-09 0 4.503e-09 0.0007 4.506e-09 0 4.56e-09 0 4.563e-09 0.0007 4.566e-09 0 4.62e-09 0 4.623e-09 0.0007 4.626e-09 0 4.68e-09 0 4.683e-09 0.0007 4.686e-09 0 4.74e-09 0 4.743e-09 0.0007 4.746e-09 0 4.8e-09 0 4.803e-09 0.0007 4.806e-09 0 4.86e-09 0 4.863e-09 0.0007 4.866e-09 0 4.92e-09 0 4.923e-09 0.0007 4.926e-09 0 4.98e-09 0 4.983e-09 0.0007 4.986e-09 0 5.04e-09 0 5.043e-09 0.0007 5.046e-09 0 5.1e-09 0 5.103e-09 0.0007 5.106e-09 0 5.16e-09 0 5.163e-09 0.0007 5.166e-09 0 5.22e-09 0 5.223e-09 0.0007 5.226e-09 0 5.28e-09 0 5.283e-09 0.0007 5.286e-09 0 5.34e-09 0 5.343e-09 0.0007 5.346e-09 0 5.4e-09 0 5.403e-09 0.0007 5.406e-09 0 5.46e-09 0 5.463e-09 0.0007 5.466e-09 0 5.52e-09 0 5.523e-09 0.0007 5.526e-09 0 5.58e-09 0 5.583e-09 0.0007 5.586e-09 0 5.64e-09 0 5.643e-09 0.0007 5.646e-09 0 5.7e-09 0 5.703e-09 0.0007 5.706e-09 0 5.76e-09 0 5.763e-09 0.0007 5.766e-09 0 5.82e-09 0 5.823e-09 0.0007 5.826e-09 0 5.88e-09 0 5.883e-09 0.0007 5.886e-09 0 5.94e-09 0 5.943e-09 0.0007 5.946e-09 0 6e-09 0 6.003e-09 0.0007 6.006e-09 0 6.06e-09 0 6.063e-09 0.0007 6.066e-09 0 6.12e-09 0 6.123e-09 0.0007 6.126e-09 0 6.18e-09 0 6.183e-09 0.0007 6.186e-09 0 6.24e-09 0 6.243e-09 0.0007 6.246e-09 0 6.3e-09 0 6.303e-09 0.0007 6.306e-09 0 6.36e-09 0 6.363e-09 0.0007 6.366e-09 0 6.42e-09 0 6.423e-09 0.0007 6.426e-09 0 6.48e-09 0 6.483e-09 0.0007 6.486e-09 0 6.54e-09 0 6.543e-09 0.0007 6.546e-09 0 6.6e-09 0 6.603e-09 0.0007 6.606e-09 0 6.66e-09 0 6.663e-09 0.0007 6.666e-09 0 6.72e-09 0 6.723e-09 0.0007 6.726e-09 0 6.78e-09 0 6.783e-09 0.0007 6.786e-09 0 6.84e-09 0 6.843e-09 0.0007 6.846e-09 0 6.9e-09 0 6.903e-09 0.0007 6.906e-09 0 6.96e-09 0 6.963e-09 0.0007 6.966e-09 0 7.02e-09 0 7.023e-09 0.0007 7.026e-09 0 7.08e-09 0 7.083e-09 0.0007 7.086e-09 0 7.14e-09 0 7.143e-09 0.0007 7.146e-09 0 7.2e-09 0 7.203e-09 0.0007 7.206e-09 0 7.26e-09 0 7.263e-09 0.0007 7.266e-09 0 7.32e-09 0 7.323e-09 0.0007 7.326e-09 0 7.38e-09 0 7.383e-09 0.0007 7.386e-09 0 7.44e-09 0 7.443e-09 0.0007 7.446e-09 0 7.5e-09 0 7.503e-09 0.0007 7.506e-09 0 7.56e-09 0 7.563e-09 0.0007 7.566e-09 0 7.62e-09 0 7.623e-09 0.0007 7.626e-09 0 7.68e-09 0 7.683e-09 0.0007 7.686e-09 0 7.74e-09 0 7.743e-09 0.0007 7.746e-09 0 7.8e-09 0 7.803e-09 0.0007 7.806e-09 0 7.86e-09 0 7.863e-09 0.0007 7.866e-09 0 7.92e-09 0 7.923e-09 0.0007 7.926e-09 0 7.98e-09 0 7.983e-09 0.0007 7.986e-09 0 8.04e-09 0 8.043e-09 0.0007 8.046e-09 0 8.1e-09 0 8.103e-09 0.0007 8.106e-09 0 8.16e-09 0 8.163e-09 0.0007 8.166e-09 0 8.22e-09 0 8.223e-09 0.0007 8.226e-09 0 8.28e-09 0 8.283e-09 0.0007 8.286e-09 0 8.34e-09 0 8.343e-09 0.0007 8.346e-09 0 8.4e-09 0 8.403e-09 0.0007 8.406e-09 0 8.46e-09 0 8.463e-09 0.0007 8.466e-09 0 8.52e-09 0 8.523e-09 0.0007 8.526e-09 0 8.58e-09 0 8.583e-09 0.0007 8.586e-09 0 8.64e-09 0 8.643e-09 0.0007 8.646e-09 0 8.7e-09 0 8.703e-09 0.0007 8.706e-09 0 8.76e-09 0 8.763e-09 0.0007 8.766e-09 0 8.82e-09 0 8.823e-09 0.0007 8.826e-09 0 8.88e-09 0 8.883e-09 0.0007 8.886e-09 0 8.94e-09 0 8.943e-09 0.0007 8.946e-09 0 9e-09 0 9.003e-09 0.0007 9.006e-09 0 9.06e-09 0 9.063e-09 0.0007 9.066e-09 0 9.12e-09 0 9.123e-09 0.0007 9.126e-09 0 9.18e-09 0 9.183e-09 0.0007 9.186e-09 0 9.24e-09 0 9.243e-09 0.0007 9.246e-09 0 9.3e-09 0 9.303e-09 0.0007 9.306e-09 0 9.36e-09 0 9.363e-09 0.0007 9.366e-09 0 9.42e-09 0 9.423e-09 0.0007 9.426e-09 0 9.48e-09 0 9.483e-09 0.0007 9.486e-09 0 9.54e-09 0 9.543e-09 0.0007 9.546e-09 0 9.6e-09 0 9.603e-09 0.0007 9.606e-09 0 9.66e-09 0 9.663e-09 0.0007 9.666e-09 0 9.72e-09 0 9.723e-09 0.0007 9.726e-09 0 9.78e-09 0 9.783e-09 0.0007 9.786e-09 0 9.84e-09 0 9.843e-09 0.0007 9.846e-09 0 9.9e-09 0 9.903e-09 0.0007 9.906e-09 0 9.96e-09 0 9.963e-09 0.0007 9.966e-09 0 1.002e-08 0 1.0023e-08 0.0007 1.0026e-08 0 1.008e-08 0 1.0083e-08 0.0007 1.0086e-08 0 1.014e-08 0 1.0143e-08 0.0007 1.0146e-08 0 1.02e-08 0 1.0203e-08 0.0007 1.0206e-08 0 1.026e-08 0 1.0263e-08 0.0007 1.0266e-08 0 1.032e-08 0 1.0323e-08 0.0007 1.0326e-08 0 1.038e-08 0 1.0383e-08 0.0007 1.0386e-08 0 1.044e-08 0 1.0443e-08 0.0007 1.0446e-08 0 1.05e-08 0 1.0503e-08 0.0007 1.0506e-08 0 1.056e-08 0 1.0563e-08 0.0007 1.0566e-08 0 1.062e-08 0 1.0623e-08 0.0007 1.0626e-08 0 1.068e-08 0 1.0683e-08 0.0007 1.0686e-08 0 1.074e-08 0 1.0743e-08 0.0007 1.0746e-08 0 1.08e-08 0 1.0803e-08 0.0007 1.0806e-08 0 1.086e-08 0 1.0863e-08 0.0007 1.0866e-08 0 1.092e-08 0 1.0923e-08 0.0007 1.0926e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.104e-08 0 1.1043e-08 0.0007 1.1046e-08 0 1.11e-08 0 1.1103e-08 0.0007 1.1106e-08 0 1.116e-08 0 1.1163e-08 0.0007 1.1166e-08 0 1.122e-08 0 1.1223e-08 0.0007 1.1226e-08 0 1.128e-08 0 1.1283e-08 0.0007 1.1286e-08 0 1.134e-08 0 1.1343e-08 0.0007 1.1346e-08 0 1.14e-08 0 1.1403e-08 0.0007 1.1406e-08 0 1.146e-08 0 1.1463e-08 0.0007 1.1466e-08 0 1.152e-08 0 1.1523e-08 0.0007 1.1526e-08 0 1.158e-08 0 1.1583e-08 0.0007 1.1586e-08 0 1.164e-08 0 1.1643e-08 0.0007 1.1646e-08 0 1.17e-08 0 1.1703e-08 0.0007 1.1706e-08 0 1.176e-08 0 1.1763e-08 0.0007 1.1766e-08 0 1.182e-08 0 1.1823e-08 0.0007 1.1826e-08 0 1.188e-08 0 1.1883e-08 0.0007 1.1886e-08 0 1.194e-08 0 1.1943e-08 0.0007 1.1946e-08 0 1.2e-08 0 1.2003e-08 0.0007 1.2006e-08 0 1.206e-08 0 1.2063e-08 0.0007 1.2066e-08 0 1.212e-08 0 1.2123e-08 0.0007 1.2126e-08 0 1.218e-08 0 1.2183e-08 0.0007 1.2186e-08 0 1.224e-08 0 1.2243e-08 0.0007 1.2246e-08 0 1.23e-08 0 1.2303e-08 0.0007 1.2306e-08 0 1.236e-08 0 1.2363e-08 0.0007 1.2366e-08 0 1.242e-08 0 1.2423e-08 0.0007 1.2426e-08 0 1.248e-08 0 1.2483e-08 0.0007 1.2486e-08 0 1.254e-08 0 1.2543e-08 0.0007 1.2546e-08 0 1.26e-08 0 1.2603e-08 0.0007 1.2606e-08 0 1.266e-08 0 1.2663e-08 0.0007 1.2666e-08 0 1.272e-08 0 1.2723e-08 0.0007 1.2726e-08 0 1.278e-08 0 1.2783e-08 0.0007 1.2786e-08 0 1.284e-08 0 1.2843e-08 0.0007 1.2846e-08 0 1.29e-08 0 1.2903e-08 0.0007 1.2906e-08 0 1.296e-08 0 1.2963e-08 0.0007 1.2966e-08 0 1.302e-08 0 1.3023e-08 0.0007 1.3026e-08 0 1.308e-08 0 1.3083e-08 0.0007 1.3086e-08 0 1.314e-08 0 1.3143e-08 0.0007 1.3146e-08 0 1.32e-08 0 1.3203e-08 0.0007 1.3206e-08 0 1.326e-08 0 1.3263e-08 0.0007 1.3266e-08 0 1.332e-08 0 1.3323e-08 0.0007 1.3326e-08 0 1.338e-08 0 1.3383e-08 0.0007 1.3386e-08 0 1.344e-08 0 1.3443e-08 0.0007 1.3446e-08 0 1.35e-08 0 1.3503e-08 0.0007 1.3506e-08 0 1.356e-08 0 1.3563e-08 0.0007 1.3566e-08 0 1.362e-08 0 1.3623e-08 0.0007 1.3626e-08 0 1.368e-08 0 1.3683e-08 0.0007 1.3686e-08 0 1.374e-08 0 1.3743e-08 0.0007 1.3746e-08 0 1.38e-08 0 1.3803e-08 0.0007 1.3806e-08 0 1.386e-08 0 1.3863e-08 0.0007 1.3866e-08 0 1.392e-08 0 1.3923e-08 0.0007 1.3926e-08 0 1.398e-08 0 1.3983e-08 0.0007 1.3986e-08 0 1.404e-08 0 1.4043e-08 0.0007 1.4046e-08 0 1.41e-08 0 1.4103e-08 0.0007 1.4106e-08 0 1.416e-08 0 1.4163e-08 0.0007 1.4166e-08 0 1.422e-08 0 1.4223e-08 0.0007 1.4226e-08 0 1.428e-08 0 1.4283e-08 0.0007 1.4286e-08 0 1.434e-08 0 1.4343e-08 0.0007 1.4346e-08 0 1.44e-08 0 1.4403e-08 0.0007 1.4406e-08 0 1.446e-08 0 1.4463e-08 0.0007 1.4466e-08 0 1.452e-08 0 1.4523e-08 0.0007 1.4526e-08 0 1.458e-08 0 1.4583e-08 0.0007 1.4586e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.47e-08 0 1.4703e-08 0.0007 1.4706e-08 0 1.476e-08 0 1.4763e-08 0.0007 1.4766e-08 0 1.482e-08 0 1.4823e-08 0.0007 1.4826e-08 0 1.488e-08 0 1.4883e-08 0.0007 1.4886e-08 0 1.494e-08 0 1.4943e-08 0.0007 1.4946e-08 0 1.5e-08 0 1.5003e-08 0.0007 1.5006e-08 0 1.506e-08 0 1.5063e-08 0.0007 1.5066e-08 0 1.512e-08 0 1.5123e-08 0.0007 1.5126e-08 0 1.518e-08 0 1.5183e-08 0.0007 1.5186e-08 0 1.524e-08 0 1.5243e-08 0.0007 1.5246e-08 0 1.53e-08 0 1.5303e-08 0.0007 1.5306e-08 0 1.536e-08 0 1.5363e-08 0.0007 1.5366e-08 0 1.542e-08 0 1.5423e-08 0.0007 1.5426e-08 0 1.548e-08 0 1.5483e-08 0.0007 1.5486e-08 0 1.554e-08 0 1.5543e-08 0.0007 1.5546e-08 0 1.56e-08 0 1.5603e-08 0.0007 1.5606e-08 0 1.566e-08 0 1.5663e-08 0.0007 1.5666e-08 0 1.572e-08 0 1.5723e-08 0.0007 1.5726e-08 0 1.578e-08 0 1.5783e-08 0.0007 1.5786e-08 0 1.584e-08 0 1.5843e-08 0.0007 1.5846e-08 0 1.59e-08 0 1.5903e-08 0.0007 1.5906e-08 0 1.596e-08 0 1.5963e-08 0.0007 1.5966e-08 0 1.602e-08 0 1.6023e-08 0.0007 1.6026e-08 0 1.608e-08 0 1.6083e-08 0.0007 1.6086e-08 0 1.614e-08 0 1.6143e-08 0.0007 1.6146e-08 0 1.62e-08 0 1.6203e-08 0.0007 1.6206e-08 0 1.626e-08 0 1.6263e-08 0.0007 1.6266e-08 0 1.632e-08 0 1.6323e-08 0.0007 1.6326e-08 0 1.638e-08 0 1.6383e-08 0.0007 1.6386e-08 0 1.644e-08 0 1.6443e-08 0.0007 1.6446e-08 0 1.65e-08 0 1.6503e-08 0.0007 1.6506e-08 0 1.656e-08 0 1.6563e-08 0.0007 1.6566e-08 0 1.662e-08 0 1.6623e-08 0.0007 1.6626e-08 0 1.668e-08 0 1.6683e-08 0.0007 1.6686e-08 0 1.674e-08 0 1.6743e-08 0.0007 1.6746e-08 0 1.68e-08 0 1.6803e-08 0.0007 1.6806e-08 0 1.686e-08 0 1.6863e-08 0.0007 1.6866e-08 0 1.692e-08 0 1.6923e-08 0.0007 1.6926e-08 0 1.698e-08 0 1.6983e-08 0.0007 1.6986e-08 0 1.704e-08 0 1.7043e-08 0.0007 1.7046e-08 0 1.71e-08 0 1.7103e-08 0.0007 1.7106e-08 0 1.716e-08 0 1.7163e-08 0.0007 1.7166e-08 0 1.722e-08 0 1.7223e-08 0.0007 1.7226e-08 0 1.728e-08 0 1.7283e-08 0.0007 1.7286e-08 0 1.734e-08 0 1.7343e-08 0.0007 1.7346e-08 0 1.74e-08 0 1.7403e-08 0.0007 1.7406e-08 0 1.746e-08 0 1.7463e-08 0.0007 1.7466e-08 0 1.752e-08 0 1.7523e-08 0.0007 1.7526e-08 0 1.758e-08 0 1.7583e-08 0.0007 1.7586e-08 0 1.764e-08 0 1.7643e-08 0.0007 1.7646e-08 0 1.77e-08 0 1.7703e-08 0.0007 1.7706e-08 0 1.776e-08 0 1.7763e-08 0.0007 1.7766e-08 0 1.782e-08 0 1.7823e-08 0.0007 1.7826e-08 0 1.788e-08 0 1.7883e-08 0.0007 1.7886e-08 0 1.794e-08 0 1.7943e-08 0.0007 1.7946e-08 0 1.8e-08 0 1.8003e-08 0.0007 1.8006e-08 0 1.806e-08 0 1.8063e-08 0.0007 1.8066e-08 0 1.812e-08 0 1.8123e-08 0.0007 1.8126e-08 0 1.818e-08 0 1.8183e-08 0.0007 1.8186e-08 0 1.824e-08 0 1.8243e-08 0.0007 1.8246e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.836e-08 0 1.8363e-08 0.0007 1.8366e-08 0 1.842e-08 0 1.8423e-08 0.0007 1.8426e-08 0 1.848e-08 0 1.8483e-08 0.0007 1.8486e-08 0 1.854e-08 0 1.8543e-08 0.0007 1.8546e-08 0 1.86e-08 0 1.8603e-08 0.0007 1.8606e-08 0 1.866e-08 0 1.8663e-08 0.0007 1.8666e-08 0 1.872e-08 0 1.8723e-08 0.0007 1.8726e-08 0 1.878e-08 0 1.8783e-08 0.0007 1.8786e-08 0 1.884e-08 0 1.8843e-08 0.0007 1.8846e-08 0 1.89e-08 0 1.8903e-08 0.0007 1.8906e-08 0 1.896e-08 0 1.8963e-08 0.0007 1.8966e-08 0 1.902e-08 0 1.9023e-08 0.0007 1.9026e-08 0 1.908e-08 0 1.9083e-08 0.0007 1.9086e-08 0 1.914e-08 0 1.9143e-08 0.0007 1.9146e-08 0 1.92e-08 0 1.9203e-08 0.0007 1.9206e-08 0 1.926e-08 0 1.9263e-08 0.0007 1.9266e-08 0 1.932e-08 0 1.9323e-08 0.0007 1.9326e-08 0 1.938e-08 0 1.9383e-08 0.0007 1.9386e-08 0 1.944e-08 0 1.9443e-08 0.0007 1.9446e-08 0 1.95e-08 0 1.9503e-08 0.0007 1.9506e-08 0 1.956e-08 0 1.9563e-08 0.0007 1.9566e-08 0 1.962e-08 0 1.9623e-08 0.0007 1.9626e-08 0 1.968e-08 0 1.9683e-08 0.0007 1.9686e-08 0 1.974e-08 0 1.9743e-08 0.0007 1.9746e-08 0 1.98e-08 0 1.9803e-08 0.0007 1.9806e-08 0 1.986e-08 0 1.9863e-08 0.0007 1.9866e-08 0 1.992e-08 0 1.9923e-08 0.0007 1.9926e-08 0 1.998e-08 0 1.9983e-08 0.0007 1.9986e-08 0 2.004e-08 0 2.0043e-08 0.0007 2.0046e-08 0 2.01e-08 0 2.0103e-08 0.0007 2.0106e-08 0 2.016e-08 0 2.0163e-08 0.0007 2.0166e-08 0 2.022e-08 0 2.0223e-08 0.0007 2.0226e-08 0 2.028e-08 0 2.0283e-08 0.0007 2.0286e-08 0 2.034e-08 0 2.0343e-08 0.0007 2.0346e-08 0 2.04e-08 0 2.0403e-08 0.0007 2.0406e-08 0 2.046e-08 0 2.0463e-08 0.0007 2.0466e-08 0 2.052e-08 0 2.0523e-08 0.0007 2.0526e-08 0 2.058e-08 0 2.0583e-08 0.0007 2.0586e-08 0 2.064e-08 0 2.0643e-08 0.0007 2.0646e-08 0 2.07e-08 0 2.0703e-08 0.0007 2.0706e-08 0 2.076e-08 0 2.0763e-08 0.0007 2.0766e-08 0 2.082e-08 0 2.0823e-08 0.0007 2.0826e-08 0 2.088e-08 0 2.0883e-08 0.0007 2.0886e-08 0 2.094e-08 0 2.0943e-08 0.0007 2.0946e-08 0 2.1e-08 0 2.1003e-08 0.0007 2.1006e-08 0 2.106e-08 0 2.1063e-08 0.0007 2.1066e-08 0 2.112e-08 0 2.1123e-08 0.0007 2.1126e-08 0 2.118e-08 0 2.1183e-08 0.0007 2.1186e-08 0 2.124e-08 0 2.1243e-08 0.0007 2.1246e-08 0 2.13e-08 0 2.1303e-08 0.0007 2.1306e-08 0 2.136e-08 0 2.1363e-08 0.0007 2.1366e-08 0 2.142e-08 0 2.1423e-08 0.0007 2.1426e-08 0 2.148e-08 0 2.1483e-08 0.0007 2.1486e-08 0 2.154e-08 0 2.1543e-08 0.0007 2.1546e-08 0 2.16e-08 0 2.1603e-08 0.0007 2.1606e-08 0 2.166e-08 0 2.1663e-08 0.0007 2.1666e-08 0 2.172e-08 0 2.1723e-08 0.0007 2.1726e-08 0 2.178e-08 0 2.1783e-08 0.0007 2.1786e-08 0 2.184e-08 0 2.1843e-08 0.0007 2.1846e-08 0 2.19e-08 0 2.1903e-08 0.0007 2.1906e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.202e-08 0 2.2023e-08 0.0007 2.2026e-08 0 2.208e-08 0 2.2083e-08 0.0007 2.2086e-08 0 2.214e-08 0 2.2143e-08 0.0007 2.2146e-08 0 2.22e-08 0 2.2203e-08 0.0007 2.2206e-08 0 2.226e-08 0 2.2263e-08 0.0007 2.2266e-08 0 2.232e-08 0 2.2323e-08 0.0007 2.2326e-08 0 2.238e-08 0 2.2383e-08 0.0007 2.2386e-08 0 2.244e-08 0 2.2443e-08 0.0007 2.2446e-08 0 2.25e-08 0 2.2503e-08 0.0007 2.2506e-08 0 2.256e-08 0 2.2563e-08 0.0007 2.2566e-08 0 2.262e-08 0 2.2623e-08 0.0007 2.2626e-08 0 2.268e-08 0 2.2683e-08 0.0007 2.2686e-08 0 2.274e-08 0 2.2743e-08 0.0007 2.2746e-08 0 2.28e-08 0 2.2803e-08 0.0007 2.2806e-08 0 2.286e-08 0 2.2863e-08 0.0007 2.2866e-08 0 2.292e-08 0 2.2923e-08 0.0007 2.2926e-08 0 2.298e-08 0 2.2983e-08 0.0007 2.2986e-08 0 2.304e-08 0 2.3043e-08 0.0007 2.3046e-08 0 2.31e-08 0 2.3103e-08 0.0007 2.3106e-08 0 2.316e-08 0 2.3163e-08 0.0007 2.3166e-08 0 2.322e-08 0 2.3223e-08 0.0007 2.3226e-08 0 2.328e-08 0 2.3283e-08 0.0007 2.3286e-08 0 2.334e-08 0 2.3343e-08 0.0007 2.3346e-08 0 2.34e-08 0 2.3403e-08 0.0007 2.3406e-08 0 2.346e-08 0 2.3463e-08 0.0007 2.3466e-08 0 2.352e-08 0 2.3523e-08 0.0007 2.3526e-08 0 2.358e-08 0 2.3583e-08 0.0007 2.3586e-08 0 2.364e-08 0 2.3643e-08 0.0007 2.3646e-08 0 2.37e-08 0 2.3703e-08 0.0007 2.3706e-08 0 2.376e-08 0 2.3763e-08 0.0007 2.3766e-08 0 2.382e-08 0 2.3823e-08 0.0007 2.3826e-08 0 2.388e-08 0 2.3883e-08 0.0007 2.3886e-08 0)
L_S4|1 G3_2_RX _S4|A1  2.067833848e-12
L_S4|2 _S4|A1 _S4|A2  4.135667696e-12
L_S4|3 _S4|A3 _S4|A4  8.271335392e-12
L_S4|T T16 _S4|T1  2.067833848e-12
L_S4|4 _S4|T1 _S4|T2  4.135667696e-12
L_S4|5 _S4|A4 _S4|Q1  4.135667696e-12
L_S4|6 _S4|Q1 S4  2.067833848e-12
B_PTL_A0|_TX|1 _PTL_A0|_TX|1 _PTL_A0|_TX|2 JJMIT AREA=2.5
B_PTL_A0|_TX|2 _PTL_A0|_TX|4 _PTL_A0|_TX|5 JJMIT AREA=2.5
I_PTL_A0|_TX|B1 0 _PTL_A0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A0|_TX|B2 0 _PTL_A0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|3  1.684e-12
L_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|6  3.596e-12
L_PTL_A0|_TX|1 A0_TX _PTL_A0|_TX|1  2.063e-12
L_PTL_A0|_TX|2 _PTL_A0|_TX|1 _PTL_A0|_TX|4  4.123e-12
L_PTL_A0|_TX|3 _PTL_A0|_TX|4 _PTL_A0|_TX|7  2.193e-12
R_PTL_A0|_TX|D _PTL_A0|_TX|7 _PTL_A0|A_PTL  1.36
L_PTL_A0|_TX|P1 _PTL_A0|_TX|2 0  5.254e-13
L_PTL_A0|_TX|P2 _PTL_A0|_TX|5 0  5.141e-13
R_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|101  2.7439617672
R_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|104  2.7439617672
L_PTL_A0|_TX|RB1 _PTL_A0|_TX|101 0  1.550338398468e-12
L_PTL_A0|_TX|RB2 _PTL_A0|_TX|104 0  1.550338398468e-12
B_PTL_A0|_RX|1 _PTL_A0|_RX|1 _PTL_A0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A0|_RX|2 _PTL_A0|_RX|4 _PTL_A0|_RX|5 JJMIT AREA=2.0
B_PTL_A0|_RX|3 _PTL_A0|_RX|7 _PTL_A0|_RX|8 JJMIT AREA=2.5
I_PTL_A0|_RX|B1 0 _PTL_A0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|3  2.777e-12
I_PTL_A0|_RX|B2 0 _PTL_A0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|6  2.685e-12
I_PTL_A0|_RX|B3 0 _PTL_A0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|9  2.764e-12
L_PTL_A0|_RX|1 _PTL_A0|A_PTL _PTL_A0|_RX|1  1.346e-12
L_PTL_A0|_RX|2 _PTL_A0|_RX|1 _PTL_A0|_RX|4  6.348e-12
L_PTL_A0|_RX|3 _PTL_A0|_RX|4 _PTL_A0|_RX|7  5.197e-12
L_PTL_A0|_RX|4 _PTL_A0|_RX|7 A0_RX  2.058e-12
L_PTL_A0|_RX|P1 _PTL_A0|_RX|2 0  4.795e-13
L_PTL_A0|_RX|P2 _PTL_A0|_RX|5 0  5.431e-13
L_PTL_A0|_RX|P3 _PTL_A0|_RX|8 0  5.339e-13
R_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|101  4.225701121488
R_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|104  3.429952209
R_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|107  2.7439617672
L_PTL_A0|_RX|RB1 _PTL_A0|_RX|101 0  2.38752113364072e-12
L_PTL_A0|_RX|RB2 _PTL_A0|_RX|104 0  1.937922998085e-12
L_PTL_A0|_RX|RB3 _PTL_A0|_RX|107 0  1.550338398468e-12
B_PTL_B0|_TX|1 _PTL_B0|_TX|1 _PTL_B0|_TX|2 JJMIT AREA=2.5
B_PTL_B0|_TX|2 _PTL_B0|_TX|4 _PTL_B0|_TX|5 JJMIT AREA=2.5
I_PTL_B0|_TX|B1 0 _PTL_B0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B0|_TX|B2 0 _PTL_B0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|3  1.684e-12
L_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|6  3.596e-12
L_PTL_B0|_TX|1 B0_TX _PTL_B0|_TX|1  2.063e-12
L_PTL_B0|_TX|2 _PTL_B0|_TX|1 _PTL_B0|_TX|4  4.123e-12
L_PTL_B0|_TX|3 _PTL_B0|_TX|4 _PTL_B0|_TX|7  2.193e-12
R_PTL_B0|_TX|D _PTL_B0|_TX|7 _PTL_B0|A_PTL  1.36
L_PTL_B0|_TX|P1 _PTL_B0|_TX|2 0  5.254e-13
L_PTL_B0|_TX|P2 _PTL_B0|_TX|5 0  5.141e-13
R_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|101  2.7439617672
R_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|104  2.7439617672
L_PTL_B0|_TX|RB1 _PTL_B0|_TX|101 0  1.550338398468e-12
L_PTL_B0|_TX|RB2 _PTL_B0|_TX|104 0  1.550338398468e-12
B_PTL_B0|_RX|1 _PTL_B0|_RX|1 _PTL_B0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B0|_RX|2 _PTL_B0|_RX|4 _PTL_B0|_RX|5 JJMIT AREA=2.0
B_PTL_B0|_RX|3 _PTL_B0|_RX|7 _PTL_B0|_RX|8 JJMIT AREA=2.5
I_PTL_B0|_RX|B1 0 _PTL_B0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|3  2.777e-12
I_PTL_B0|_RX|B2 0 _PTL_B0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|6  2.685e-12
I_PTL_B0|_RX|B3 0 _PTL_B0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|9  2.764e-12
L_PTL_B0|_RX|1 _PTL_B0|A_PTL _PTL_B0|_RX|1  1.346e-12
L_PTL_B0|_RX|2 _PTL_B0|_RX|1 _PTL_B0|_RX|4  6.348e-12
L_PTL_B0|_RX|3 _PTL_B0|_RX|4 _PTL_B0|_RX|7  5.197e-12
L_PTL_B0|_RX|4 _PTL_B0|_RX|7 B0_RX  2.058e-12
L_PTL_B0|_RX|P1 _PTL_B0|_RX|2 0  4.795e-13
L_PTL_B0|_RX|P2 _PTL_B0|_RX|5 0  5.431e-13
L_PTL_B0|_RX|P3 _PTL_B0|_RX|8 0  5.339e-13
R_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|101  4.225701121488
R_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|104  3.429952209
R_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|107  2.7439617672
L_PTL_B0|_RX|RB1 _PTL_B0|_RX|101 0  2.38752113364072e-12
L_PTL_B0|_RX|RB2 _PTL_B0|_RX|104 0  1.937922998085e-12
L_PTL_B0|_RX|RB3 _PTL_B0|_RX|107 0  1.550338398468e-12
B_PTL_A1|_TX|1 _PTL_A1|_TX|1 _PTL_A1|_TX|2 JJMIT AREA=2.5
B_PTL_A1|_TX|2 _PTL_A1|_TX|4 _PTL_A1|_TX|5 JJMIT AREA=2.5
I_PTL_A1|_TX|B1 0 _PTL_A1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A1|_TX|B2 0 _PTL_A1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|3  1.684e-12
L_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|6  3.596e-12
L_PTL_A1|_TX|1 A1_TX _PTL_A1|_TX|1  2.063e-12
L_PTL_A1|_TX|2 _PTL_A1|_TX|1 _PTL_A1|_TX|4  4.123e-12
L_PTL_A1|_TX|3 _PTL_A1|_TX|4 _PTL_A1|_TX|7  2.193e-12
R_PTL_A1|_TX|D _PTL_A1|_TX|7 _PTL_A1|A_PTL  1.36
L_PTL_A1|_TX|P1 _PTL_A1|_TX|2 0  5.254e-13
L_PTL_A1|_TX|P2 _PTL_A1|_TX|5 0  5.141e-13
R_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|101  2.7439617672
R_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|104  2.7439617672
L_PTL_A1|_TX|RB1 _PTL_A1|_TX|101 0  1.550338398468e-12
L_PTL_A1|_TX|RB2 _PTL_A1|_TX|104 0  1.550338398468e-12
B_PTL_A1|_RX|1 _PTL_A1|_RX|1 _PTL_A1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A1|_RX|2 _PTL_A1|_RX|4 _PTL_A1|_RX|5 JJMIT AREA=2.0
B_PTL_A1|_RX|3 _PTL_A1|_RX|7 _PTL_A1|_RX|8 JJMIT AREA=2.5
I_PTL_A1|_RX|B1 0 _PTL_A1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|3  2.777e-12
I_PTL_A1|_RX|B2 0 _PTL_A1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|6  2.685e-12
I_PTL_A1|_RX|B3 0 _PTL_A1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|9  2.764e-12
L_PTL_A1|_RX|1 _PTL_A1|A_PTL _PTL_A1|_RX|1  1.346e-12
L_PTL_A1|_RX|2 _PTL_A1|_RX|1 _PTL_A1|_RX|4  6.348e-12
L_PTL_A1|_RX|3 _PTL_A1|_RX|4 _PTL_A1|_RX|7  5.197e-12
L_PTL_A1|_RX|4 _PTL_A1|_RX|7 A1_RX  2.058e-12
L_PTL_A1|_RX|P1 _PTL_A1|_RX|2 0  4.795e-13
L_PTL_A1|_RX|P2 _PTL_A1|_RX|5 0  5.431e-13
L_PTL_A1|_RX|P3 _PTL_A1|_RX|8 0  5.339e-13
R_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|101  4.225701121488
R_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|104  3.429952209
R_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|107  2.7439617672
L_PTL_A1|_RX|RB1 _PTL_A1|_RX|101 0  2.38752113364072e-12
L_PTL_A1|_RX|RB2 _PTL_A1|_RX|104 0  1.937922998085e-12
L_PTL_A1|_RX|RB3 _PTL_A1|_RX|107 0  1.550338398468e-12
B_PTL_B1|_TX|1 _PTL_B1|_TX|1 _PTL_B1|_TX|2 JJMIT AREA=2.5
B_PTL_B1|_TX|2 _PTL_B1|_TX|4 _PTL_B1|_TX|5 JJMIT AREA=2.5
I_PTL_B1|_TX|B1 0 _PTL_B1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B1|_TX|B2 0 _PTL_B1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|3  1.684e-12
L_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|6  3.596e-12
L_PTL_B1|_TX|1 B1_TX _PTL_B1|_TX|1  2.063e-12
L_PTL_B1|_TX|2 _PTL_B1|_TX|1 _PTL_B1|_TX|4  4.123e-12
L_PTL_B1|_TX|3 _PTL_B1|_TX|4 _PTL_B1|_TX|7  2.193e-12
R_PTL_B1|_TX|D _PTL_B1|_TX|7 _PTL_B1|A_PTL  1.36
L_PTL_B1|_TX|P1 _PTL_B1|_TX|2 0  5.254e-13
L_PTL_B1|_TX|P2 _PTL_B1|_TX|5 0  5.141e-13
R_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|101  2.7439617672
R_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|104  2.7439617672
L_PTL_B1|_TX|RB1 _PTL_B1|_TX|101 0  1.550338398468e-12
L_PTL_B1|_TX|RB2 _PTL_B1|_TX|104 0  1.550338398468e-12
B_PTL_B1|_RX|1 _PTL_B1|_RX|1 _PTL_B1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B1|_RX|2 _PTL_B1|_RX|4 _PTL_B1|_RX|5 JJMIT AREA=2.0
B_PTL_B1|_RX|3 _PTL_B1|_RX|7 _PTL_B1|_RX|8 JJMIT AREA=2.5
I_PTL_B1|_RX|B1 0 _PTL_B1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|3  2.777e-12
I_PTL_B1|_RX|B2 0 _PTL_B1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|6  2.685e-12
I_PTL_B1|_RX|B3 0 _PTL_B1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|9  2.764e-12
L_PTL_B1|_RX|1 _PTL_B1|A_PTL _PTL_B1|_RX|1  1.346e-12
L_PTL_B1|_RX|2 _PTL_B1|_RX|1 _PTL_B1|_RX|4  6.348e-12
L_PTL_B1|_RX|3 _PTL_B1|_RX|4 _PTL_B1|_RX|7  5.197e-12
L_PTL_B1|_RX|4 _PTL_B1|_RX|7 B1_RX  2.058e-12
L_PTL_B1|_RX|P1 _PTL_B1|_RX|2 0  4.795e-13
L_PTL_B1|_RX|P2 _PTL_B1|_RX|5 0  5.431e-13
L_PTL_B1|_RX|P3 _PTL_B1|_RX|8 0  5.339e-13
R_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|101  4.225701121488
R_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|104  3.429952209
R_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|107  2.7439617672
L_PTL_B1|_RX|RB1 _PTL_B1|_RX|101 0  2.38752113364072e-12
L_PTL_B1|_RX|RB2 _PTL_B1|_RX|104 0  1.937922998085e-12
L_PTL_B1|_RX|RB3 _PTL_B1|_RX|107 0  1.550338398468e-12
B_PTL_A2|_TX|1 _PTL_A2|_TX|1 _PTL_A2|_TX|2 JJMIT AREA=2.5
B_PTL_A2|_TX|2 _PTL_A2|_TX|4 _PTL_A2|_TX|5 JJMIT AREA=2.5
I_PTL_A2|_TX|B1 0 _PTL_A2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A2|_TX|B2 0 _PTL_A2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|3  1.684e-12
L_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|6  3.596e-12
L_PTL_A2|_TX|1 A2_TX _PTL_A2|_TX|1  2.063e-12
L_PTL_A2|_TX|2 _PTL_A2|_TX|1 _PTL_A2|_TX|4  4.123e-12
L_PTL_A2|_TX|3 _PTL_A2|_TX|4 _PTL_A2|_TX|7  2.193e-12
R_PTL_A2|_TX|D _PTL_A2|_TX|7 _PTL_A2|A_PTL  1.36
L_PTL_A2|_TX|P1 _PTL_A2|_TX|2 0  5.254e-13
L_PTL_A2|_TX|P2 _PTL_A2|_TX|5 0  5.141e-13
R_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|101  2.7439617672
R_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|104  2.7439617672
L_PTL_A2|_TX|RB1 _PTL_A2|_TX|101 0  1.550338398468e-12
L_PTL_A2|_TX|RB2 _PTL_A2|_TX|104 0  1.550338398468e-12
B_PTL_A2|_RX|1 _PTL_A2|_RX|1 _PTL_A2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A2|_RX|2 _PTL_A2|_RX|4 _PTL_A2|_RX|5 JJMIT AREA=2.0
B_PTL_A2|_RX|3 _PTL_A2|_RX|7 _PTL_A2|_RX|8 JJMIT AREA=2.5
I_PTL_A2|_RX|B1 0 _PTL_A2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|3  2.777e-12
I_PTL_A2|_RX|B2 0 _PTL_A2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|6  2.685e-12
I_PTL_A2|_RX|B3 0 _PTL_A2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|9  2.764e-12
L_PTL_A2|_RX|1 _PTL_A2|A_PTL _PTL_A2|_RX|1  1.346e-12
L_PTL_A2|_RX|2 _PTL_A2|_RX|1 _PTL_A2|_RX|4  6.348e-12
L_PTL_A2|_RX|3 _PTL_A2|_RX|4 _PTL_A2|_RX|7  5.197e-12
L_PTL_A2|_RX|4 _PTL_A2|_RX|7 A2_RX  2.058e-12
L_PTL_A2|_RX|P1 _PTL_A2|_RX|2 0  4.795e-13
L_PTL_A2|_RX|P2 _PTL_A2|_RX|5 0  5.431e-13
L_PTL_A2|_RX|P3 _PTL_A2|_RX|8 0  5.339e-13
R_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|101  4.225701121488
R_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|104  3.429952209
R_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|107  2.7439617672
L_PTL_A2|_RX|RB1 _PTL_A2|_RX|101 0  2.38752113364072e-12
L_PTL_A2|_RX|RB2 _PTL_A2|_RX|104 0  1.937922998085e-12
L_PTL_A2|_RX|RB3 _PTL_A2|_RX|107 0  1.550338398468e-12
B_PTL_B2|_TX|1 _PTL_B2|_TX|1 _PTL_B2|_TX|2 JJMIT AREA=2.5
B_PTL_B2|_TX|2 _PTL_B2|_TX|4 _PTL_B2|_TX|5 JJMIT AREA=2.5
I_PTL_B2|_TX|B1 0 _PTL_B2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B2|_TX|B2 0 _PTL_B2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|3  1.684e-12
L_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|6  3.596e-12
L_PTL_B2|_TX|1 B2_TX _PTL_B2|_TX|1  2.063e-12
L_PTL_B2|_TX|2 _PTL_B2|_TX|1 _PTL_B2|_TX|4  4.123e-12
L_PTL_B2|_TX|3 _PTL_B2|_TX|4 _PTL_B2|_TX|7  2.193e-12
R_PTL_B2|_TX|D _PTL_B2|_TX|7 _PTL_B2|A_PTL  1.36
L_PTL_B2|_TX|P1 _PTL_B2|_TX|2 0  5.254e-13
L_PTL_B2|_TX|P2 _PTL_B2|_TX|5 0  5.141e-13
R_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|101  2.7439617672
R_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|104  2.7439617672
L_PTL_B2|_TX|RB1 _PTL_B2|_TX|101 0  1.550338398468e-12
L_PTL_B2|_TX|RB2 _PTL_B2|_TX|104 0  1.550338398468e-12
B_PTL_B2|_RX|1 _PTL_B2|_RX|1 _PTL_B2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B2|_RX|2 _PTL_B2|_RX|4 _PTL_B2|_RX|5 JJMIT AREA=2.0
B_PTL_B2|_RX|3 _PTL_B2|_RX|7 _PTL_B2|_RX|8 JJMIT AREA=2.5
I_PTL_B2|_RX|B1 0 _PTL_B2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|3  2.777e-12
I_PTL_B2|_RX|B2 0 _PTL_B2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|6  2.685e-12
I_PTL_B2|_RX|B3 0 _PTL_B2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|9  2.764e-12
L_PTL_B2|_RX|1 _PTL_B2|A_PTL _PTL_B2|_RX|1  1.346e-12
L_PTL_B2|_RX|2 _PTL_B2|_RX|1 _PTL_B2|_RX|4  6.348e-12
L_PTL_B2|_RX|3 _PTL_B2|_RX|4 _PTL_B2|_RX|7  5.197e-12
L_PTL_B2|_RX|4 _PTL_B2|_RX|7 B2_RX  2.058e-12
L_PTL_B2|_RX|P1 _PTL_B2|_RX|2 0  4.795e-13
L_PTL_B2|_RX|P2 _PTL_B2|_RX|5 0  5.431e-13
L_PTL_B2|_RX|P3 _PTL_B2|_RX|8 0  5.339e-13
R_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|101  4.225701121488
R_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|104  3.429952209
R_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|107  2.7439617672
L_PTL_B2|_RX|RB1 _PTL_B2|_RX|101 0  2.38752113364072e-12
L_PTL_B2|_RX|RB2 _PTL_B2|_RX|104 0  1.937922998085e-12
L_PTL_B2|_RX|RB3 _PTL_B2|_RX|107 0  1.550338398468e-12
B_PTL_A3|_TX|1 _PTL_A3|_TX|1 _PTL_A3|_TX|2 JJMIT AREA=2.5
B_PTL_A3|_TX|2 _PTL_A3|_TX|4 _PTL_A3|_TX|5 JJMIT AREA=2.5
I_PTL_A3|_TX|B1 0 _PTL_A3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A3|_TX|B2 0 _PTL_A3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|3  1.684e-12
L_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|6  3.596e-12
L_PTL_A3|_TX|1 A3_TX _PTL_A3|_TX|1  2.063e-12
L_PTL_A3|_TX|2 _PTL_A3|_TX|1 _PTL_A3|_TX|4  4.123e-12
L_PTL_A3|_TX|3 _PTL_A3|_TX|4 _PTL_A3|_TX|7  2.193e-12
R_PTL_A3|_TX|D _PTL_A3|_TX|7 _PTL_A3|A_PTL  1.36
L_PTL_A3|_TX|P1 _PTL_A3|_TX|2 0  5.254e-13
L_PTL_A3|_TX|P2 _PTL_A3|_TX|5 0  5.141e-13
R_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|101  2.7439617672
R_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|104  2.7439617672
L_PTL_A3|_TX|RB1 _PTL_A3|_TX|101 0  1.550338398468e-12
L_PTL_A3|_TX|RB2 _PTL_A3|_TX|104 0  1.550338398468e-12
B_PTL_A3|_RX|1 _PTL_A3|_RX|1 _PTL_A3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A3|_RX|2 _PTL_A3|_RX|4 _PTL_A3|_RX|5 JJMIT AREA=2.0
B_PTL_A3|_RX|3 _PTL_A3|_RX|7 _PTL_A3|_RX|8 JJMIT AREA=2.5
I_PTL_A3|_RX|B1 0 _PTL_A3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|3  2.777e-12
I_PTL_A3|_RX|B2 0 _PTL_A3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|6  2.685e-12
I_PTL_A3|_RX|B3 0 _PTL_A3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|9  2.764e-12
L_PTL_A3|_RX|1 _PTL_A3|A_PTL _PTL_A3|_RX|1  1.346e-12
L_PTL_A3|_RX|2 _PTL_A3|_RX|1 _PTL_A3|_RX|4  6.348e-12
L_PTL_A3|_RX|3 _PTL_A3|_RX|4 _PTL_A3|_RX|7  5.197e-12
L_PTL_A3|_RX|4 _PTL_A3|_RX|7 A3_RX  2.058e-12
L_PTL_A3|_RX|P1 _PTL_A3|_RX|2 0  4.795e-13
L_PTL_A3|_RX|P2 _PTL_A3|_RX|5 0  5.431e-13
L_PTL_A3|_RX|P3 _PTL_A3|_RX|8 0  5.339e-13
R_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|101  4.225701121488
R_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|104  3.429952209
R_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|107  2.7439617672
L_PTL_A3|_RX|RB1 _PTL_A3|_RX|101 0  2.38752113364072e-12
L_PTL_A3|_RX|RB2 _PTL_A3|_RX|104 0  1.937922998085e-12
L_PTL_A3|_RX|RB3 _PTL_A3|_RX|107 0  1.550338398468e-12
B_PTL_B3|_TX|1 _PTL_B3|_TX|1 _PTL_B3|_TX|2 JJMIT AREA=2.5
B_PTL_B3|_TX|2 _PTL_B3|_TX|4 _PTL_B3|_TX|5 JJMIT AREA=2.5
I_PTL_B3|_TX|B1 0 _PTL_B3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B3|_TX|B2 0 _PTL_B3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|3  1.684e-12
L_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|6  3.596e-12
L_PTL_B3|_TX|1 B3_TX _PTL_B3|_TX|1  2.063e-12
L_PTL_B3|_TX|2 _PTL_B3|_TX|1 _PTL_B3|_TX|4  4.123e-12
L_PTL_B3|_TX|3 _PTL_B3|_TX|4 _PTL_B3|_TX|7  2.193e-12
R_PTL_B3|_TX|D _PTL_B3|_TX|7 _PTL_B3|A_PTL  1.36
L_PTL_B3|_TX|P1 _PTL_B3|_TX|2 0  5.254e-13
L_PTL_B3|_TX|P2 _PTL_B3|_TX|5 0  5.141e-13
R_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|101  2.7439617672
R_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|104  2.7439617672
L_PTL_B3|_TX|RB1 _PTL_B3|_TX|101 0  1.550338398468e-12
L_PTL_B3|_TX|RB2 _PTL_B3|_TX|104 0  1.550338398468e-12
B_PTL_B3|_RX|1 _PTL_B3|_RX|1 _PTL_B3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B3|_RX|2 _PTL_B3|_RX|4 _PTL_B3|_RX|5 JJMIT AREA=2.0
B_PTL_B3|_RX|3 _PTL_B3|_RX|7 _PTL_B3|_RX|8 JJMIT AREA=2.5
I_PTL_B3|_RX|B1 0 _PTL_B3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|3  2.777e-12
I_PTL_B3|_RX|B2 0 _PTL_B3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|6  2.685e-12
I_PTL_B3|_RX|B3 0 _PTL_B3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|9  2.764e-12
L_PTL_B3|_RX|1 _PTL_B3|A_PTL _PTL_B3|_RX|1  1.346e-12
L_PTL_B3|_RX|2 _PTL_B3|_RX|1 _PTL_B3|_RX|4  6.348e-12
L_PTL_B3|_RX|3 _PTL_B3|_RX|4 _PTL_B3|_RX|7  5.197e-12
L_PTL_B3|_RX|4 _PTL_B3|_RX|7 B3_RX  2.058e-12
L_PTL_B3|_RX|P1 _PTL_B3|_RX|2 0  4.795e-13
L_PTL_B3|_RX|P2 _PTL_B3|_RX|5 0  5.431e-13
L_PTL_B3|_RX|P3 _PTL_B3|_RX|8 0  5.339e-13
R_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|101  4.225701121488
R_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|104  3.429952209
R_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|107  2.7439617672
L_PTL_B3|_RX|RB1 _PTL_B3|_RX|101 0  2.38752113364072e-12
L_PTL_B3|_RX|RB2 _PTL_B3|_RX|104 0  1.937922998085e-12
L_PTL_B3|_RX|RB3 _PTL_B3|_RX|107 0  1.550338398468e-12
LI0|_SPL_A|1 A0_RX I0|_SPL_A|D1  2e-12
LI0|_SPL_A|2 I0|_SPL_A|D1 I0|_SPL_A|D2  4.135667696e-12
LI0|_SPL_A|3 I0|_SPL_A|D2 I0|_SPL_A|JCT  9.84682784761905e-13
LI0|_SPL_A|4 I0|_SPL_A|JCT I0|_SPL_A|QA1  9.84682784761905e-13
LI0|_SPL_A|5 I0|_SPL_A|QA1 I0|A1  2e-12
LI0|_SPL_A|6 I0|_SPL_A|JCT I0|_SPL_A|QB1  9.84682784761905e-13
LI0|_SPL_A|7 I0|_SPL_A|QB1 I0|A2  2e-12
LI0|_SPL_B|1 B0_RX I0|_SPL_B|D1  2e-12
LI0|_SPL_B|2 I0|_SPL_B|D1 I0|_SPL_B|D2  4.135667696e-12
LI0|_SPL_B|3 I0|_SPL_B|D2 I0|_SPL_B|JCT  9.84682784761905e-13
LI0|_SPL_B|4 I0|_SPL_B|JCT I0|_SPL_B|QA1  9.84682784761905e-13
LI0|_SPL_B|5 I0|_SPL_B|QA1 I0|B1  2e-12
LI0|_SPL_B|6 I0|_SPL_B|JCT I0|_SPL_B|QB1  9.84682784761905e-13
LI0|_SPL_B|7 I0|_SPL_B|QB1 I0|B2  2e-12
LI0|_DFF_A|1 I0|A1 I0|_DFF_A|A1  2.067833848e-12
LI0|_DFF_A|2 I0|_DFF_A|A1 I0|_DFF_A|A2  4.135667696e-12
LI0|_DFF_A|3 I0|_DFF_A|A3 I0|_DFF_A|A4  8.271335392e-12
LI0|_DFF_A|T T00 I0|_DFF_A|T1  2.067833848e-12
LI0|_DFF_A|4 I0|_DFF_A|T1 I0|_DFF_A|T2  4.135667696e-12
LI0|_DFF_A|5 I0|_DFF_A|A4 I0|_DFF_A|Q1  4.135667696e-12
LI0|_DFF_A|6 I0|_DFF_A|Q1 I0|A1_SYNC  2.067833848e-12
LI0|_DFF_B|1 I0|B1 I0|_DFF_B|A1  2.067833848e-12
LI0|_DFF_B|2 I0|_DFF_B|A1 I0|_DFF_B|A2  4.135667696e-12
LI0|_DFF_B|3 I0|_DFF_B|A3 I0|_DFF_B|A4  8.271335392e-12
LI0|_DFF_B|T T00 I0|_DFF_B|T1  2.067833848e-12
LI0|_DFF_B|4 I0|_DFF_B|T1 I0|_DFF_B|T2  4.135667696e-12
LI0|_DFF_B|5 I0|_DFF_B|A4 I0|_DFF_B|Q1  4.135667696e-12
LI0|_DFF_B|6 I0|_DFF_B|Q1 I0|B1_SYNC  2.067833848e-12
LI0|_XOR|A1 I0|A2 I0|_XOR|A1  2.067833848e-12
LI0|_XOR|A2 I0|_XOR|A1 I0|_XOR|A2  4.135667696e-12
LI0|_XOR|A3 I0|_XOR|A3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|B1 I0|B2 I0|_XOR|B1  2.067833848e-12
LI0|_XOR|B2 I0|_XOR|B1 I0|_XOR|B2  4.135667696e-12
LI0|_XOR|B3 I0|_XOR|B3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|T1 T00 I0|_XOR|T1  2.067833848e-12
LI0|_XOR|T2 I0|_XOR|T1 I0|_XOR|T2  4.135667696e-12
LI0|_XOR|Q2 I0|_XOR|ABTQ I0|_XOR|Q1  4.135667696e-12
LI0|_XOR|Q1 I0|_XOR|Q1 IP0_0  2.067833848e-12
LI0|_AND|A1 I0|A1_SYNC I0|_AND|A1  2.067833848e-12
LI0|_AND|A2 I0|_AND|A1 I0|_AND|A2  4.135667696e-12
LI0|_AND|A3 I0|_AND|A3 I0|_AND|Q3  1.2e-12
LI0|_AND|B1 I0|B1_SYNC I0|_AND|B1  2.067833848e-12
LI0|_AND|B2 I0|_AND|B1 I0|_AND|B2  4.135667696e-12
LI0|_AND|B3 I0|_AND|B3 I0|_AND|Q3  1.2e-12
LI0|_AND|Q3 I0|_AND|Q3 I0|_AND|Q2  4.135667696e-12
LI0|_AND|Q2 I0|_AND|Q2 I0|_AND|Q1  4.135667696e-12
LI0|_AND|Q1 I0|_AND|Q1 IG0_0  2.067833848e-12
LI1|_SPL_A|1 A1_RX I1|_SPL_A|D1  2e-12
LI1|_SPL_A|2 I1|_SPL_A|D1 I1|_SPL_A|D2  4.135667696e-12
LI1|_SPL_A|3 I1|_SPL_A|D2 I1|_SPL_A|JCT  9.84682784761905e-13
LI1|_SPL_A|4 I1|_SPL_A|JCT I1|_SPL_A|QA1  9.84682784761905e-13
LI1|_SPL_A|5 I1|_SPL_A|QA1 I1|A1  2e-12
LI1|_SPL_A|6 I1|_SPL_A|JCT I1|_SPL_A|QB1  9.84682784761905e-13
LI1|_SPL_A|7 I1|_SPL_A|QB1 I1|A2  2e-12
LI1|_SPL_B|1 B1_RX I1|_SPL_B|D1  2e-12
LI1|_SPL_B|2 I1|_SPL_B|D1 I1|_SPL_B|D2  4.135667696e-12
LI1|_SPL_B|3 I1|_SPL_B|D2 I1|_SPL_B|JCT  9.84682784761905e-13
LI1|_SPL_B|4 I1|_SPL_B|JCT I1|_SPL_B|QA1  9.84682784761905e-13
LI1|_SPL_B|5 I1|_SPL_B|QA1 I1|B1  2e-12
LI1|_SPL_B|6 I1|_SPL_B|JCT I1|_SPL_B|QB1  9.84682784761905e-13
LI1|_SPL_B|7 I1|_SPL_B|QB1 I1|B2  2e-12
LI1|_DFF_A|1 I1|A1 I1|_DFF_A|A1  2.067833848e-12
LI1|_DFF_A|2 I1|_DFF_A|A1 I1|_DFF_A|A2  4.135667696e-12
LI1|_DFF_A|3 I1|_DFF_A|A3 I1|_DFF_A|A4  8.271335392e-12
LI1|_DFF_A|T T01 I1|_DFF_A|T1  2.067833848e-12
LI1|_DFF_A|4 I1|_DFF_A|T1 I1|_DFF_A|T2  4.135667696e-12
LI1|_DFF_A|5 I1|_DFF_A|A4 I1|_DFF_A|Q1  4.135667696e-12
LI1|_DFF_A|6 I1|_DFF_A|Q1 I1|A1_SYNC  2.067833848e-12
LI1|_DFF_B|1 I1|B1 I1|_DFF_B|A1  2.067833848e-12
LI1|_DFF_B|2 I1|_DFF_B|A1 I1|_DFF_B|A2  4.135667696e-12
LI1|_DFF_B|3 I1|_DFF_B|A3 I1|_DFF_B|A4  8.271335392e-12
LI1|_DFF_B|T T01 I1|_DFF_B|T1  2.067833848e-12
LI1|_DFF_B|4 I1|_DFF_B|T1 I1|_DFF_B|T2  4.135667696e-12
LI1|_DFF_B|5 I1|_DFF_B|A4 I1|_DFF_B|Q1  4.135667696e-12
LI1|_DFF_B|6 I1|_DFF_B|Q1 I1|B1_SYNC  2.067833848e-12
LI1|_XOR|A1 I1|A2 I1|_XOR|A1  2.067833848e-12
LI1|_XOR|A2 I1|_XOR|A1 I1|_XOR|A2  4.135667696e-12
LI1|_XOR|A3 I1|_XOR|A3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|B1 I1|B2 I1|_XOR|B1  2.067833848e-12
LI1|_XOR|B2 I1|_XOR|B1 I1|_XOR|B2  4.135667696e-12
LI1|_XOR|B3 I1|_XOR|B3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|T1 T01 I1|_XOR|T1  2.067833848e-12
LI1|_XOR|T2 I1|_XOR|T1 I1|_XOR|T2  4.135667696e-12
LI1|_XOR|Q2 I1|_XOR|ABTQ I1|_XOR|Q1  4.135667696e-12
LI1|_XOR|Q1 I1|_XOR|Q1 IP1_0  2.067833848e-12
LI1|_AND|A1 I1|A1_SYNC I1|_AND|A1  2.067833848e-12
LI1|_AND|A2 I1|_AND|A1 I1|_AND|A2  4.135667696e-12
LI1|_AND|A3 I1|_AND|A3 I1|_AND|Q3  1.2e-12
LI1|_AND|B1 I1|B1_SYNC I1|_AND|B1  2.067833848e-12
LI1|_AND|B2 I1|_AND|B1 I1|_AND|B2  4.135667696e-12
LI1|_AND|B3 I1|_AND|B3 I1|_AND|Q3  1.2e-12
LI1|_AND|Q3 I1|_AND|Q3 I1|_AND|Q2  4.135667696e-12
LI1|_AND|Q2 I1|_AND|Q2 I1|_AND|Q1  4.135667696e-12
LI1|_AND|Q1 I1|_AND|Q1 IG1_0  2.067833848e-12
LI2|_SPL_A|1 A2_RX I2|_SPL_A|D1  2e-12
LI2|_SPL_A|2 I2|_SPL_A|D1 I2|_SPL_A|D2  4.135667696e-12
LI2|_SPL_A|3 I2|_SPL_A|D2 I2|_SPL_A|JCT  9.84682784761905e-13
LI2|_SPL_A|4 I2|_SPL_A|JCT I2|_SPL_A|QA1  9.84682784761905e-13
LI2|_SPL_A|5 I2|_SPL_A|QA1 I2|A1  2e-12
LI2|_SPL_A|6 I2|_SPL_A|JCT I2|_SPL_A|QB1  9.84682784761905e-13
LI2|_SPL_A|7 I2|_SPL_A|QB1 I2|A2  2e-12
LI2|_SPL_B|1 B2_RX I2|_SPL_B|D1  2e-12
LI2|_SPL_B|2 I2|_SPL_B|D1 I2|_SPL_B|D2  4.135667696e-12
LI2|_SPL_B|3 I2|_SPL_B|D2 I2|_SPL_B|JCT  9.84682784761905e-13
LI2|_SPL_B|4 I2|_SPL_B|JCT I2|_SPL_B|QA1  9.84682784761905e-13
LI2|_SPL_B|5 I2|_SPL_B|QA1 I2|B1  2e-12
LI2|_SPL_B|6 I2|_SPL_B|JCT I2|_SPL_B|QB1  9.84682784761905e-13
LI2|_SPL_B|7 I2|_SPL_B|QB1 I2|B2  2e-12
LI2|_DFF_A|1 I2|A1 I2|_DFF_A|A1  2.067833848e-12
LI2|_DFF_A|2 I2|_DFF_A|A1 I2|_DFF_A|A2  4.135667696e-12
LI2|_DFF_A|3 I2|_DFF_A|A3 I2|_DFF_A|A4  8.271335392e-12
LI2|_DFF_A|T T02 I2|_DFF_A|T1  2.067833848e-12
LI2|_DFF_A|4 I2|_DFF_A|T1 I2|_DFF_A|T2  4.135667696e-12
LI2|_DFF_A|5 I2|_DFF_A|A4 I2|_DFF_A|Q1  4.135667696e-12
LI2|_DFF_A|6 I2|_DFF_A|Q1 I2|A1_SYNC  2.067833848e-12
LI2|_DFF_B|1 I2|B1 I2|_DFF_B|A1  2.067833848e-12
LI2|_DFF_B|2 I2|_DFF_B|A1 I2|_DFF_B|A2  4.135667696e-12
LI2|_DFF_B|3 I2|_DFF_B|A3 I2|_DFF_B|A4  8.271335392e-12
LI2|_DFF_B|T T02 I2|_DFF_B|T1  2.067833848e-12
LI2|_DFF_B|4 I2|_DFF_B|T1 I2|_DFF_B|T2  4.135667696e-12
LI2|_DFF_B|5 I2|_DFF_B|A4 I2|_DFF_B|Q1  4.135667696e-12
LI2|_DFF_B|6 I2|_DFF_B|Q1 I2|B1_SYNC  2.067833848e-12
LI2|_XOR|A1 I2|A2 I2|_XOR|A1  2.067833848e-12
LI2|_XOR|A2 I2|_XOR|A1 I2|_XOR|A2  4.135667696e-12
LI2|_XOR|A3 I2|_XOR|A3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|B1 I2|B2 I2|_XOR|B1  2.067833848e-12
LI2|_XOR|B2 I2|_XOR|B1 I2|_XOR|B2  4.135667696e-12
LI2|_XOR|B3 I2|_XOR|B3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|T1 T02 I2|_XOR|T1  2.067833848e-12
LI2|_XOR|T2 I2|_XOR|T1 I2|_XOR|T2  4.135667696e-12
LI2|_XOR|Q2 I2|_XOR|ABTQ I2|_XOR|Q1  4.135667696e-12
LI2|_XOR|Q1 I2|_XOR|Q1 IP2_0  2.067833848e-12
LI2|_AND|A1 I2|A1_SYNC I2|_AND|A1  2.067833848e-12
LI2|_AND|A2 I2|_AND|A1 I2|_AND|A2  4.135667696e-12
LI2|_AND|A3 I2|_AND|A3 I2|_AND|Q3  1.2e-12
LI2|_AND|B1 I2|B1_SYNC I2|_AND|B1  2.067833848e-12
LI2|_AND|B2 I2|_AND|B1 I2|_AND|B2  4.135667696e-12
LI2|_AND|B3 I2|_AND|B3 I2|_AND|Q3  1.2e-12
LI2|_AND|Q3 I2|_AND|Q3 I2|_AND|Q2  4.135667696e-12
LI2|_AND|Q2 I2|_AND|Q2 I2|_AND|Q1  4.135667696e-12
LI2|_AND|Q1 I2|_AND|Q1 IG2_0  2.067833848e-12
LI3|_SPL_A|1 A3_RX I3|_SPL_A|D1  2e-12
LI3|_SPL_A|2 I3|_SPL_A|D1 I3|_SPL_A|D2  4.135667696e-12
LI3|_SPL_A|3 I3|_SPL_A|D2 I3|_SPL_A|JCT  9.84682784761905e-13
LI3|_SPL_A|4 I3|_SPL_A|JCT I3|_SPL_A|QA1  9.84682784761905e-13
LI3|_SPL_A|5 I3|_SPL_A|QA1 I3|A1  2e-12
LI3|_SPL_A|6 I3|_SPL_A|JCT I3|_SPL_A|QB1  9.84682784761905e-13
LI3|_SPL_A|7 I3|_SPL_A|QB1 I3|A2  2e-12
LI3|_SPL_B|1 B3_RX I3|_SPL_B|D1  2e-12
LI3|_SPL_B|2 I3|_SPL_B|D1 I3|_SPL_B|D2  4.135667696e-12
LI3|_SPL_B|3 I3|_SPL_B|D2 I3|_SPL_B|JCT  9.84682784761905e-13
LI3|_SPL_B|4 I3|_SPL_B|JCT I3|_SPL_B|QA1  9.84682784761905e-13
LI3|_SPL_B|5 I3|_SPL_B|QA1 I3|B1  2e-12
LI3|_SPL_B|6 I3|_SPL_B|JCT I3|_SPL_B|QB1  9.84682784761905e-13
LI3|_SPL_B|7 I3|_SPL_B|QB1 I3|B2  2e-12
LI3|_DFF_A|1 I3|A1 I3|_DFF_A|A1  2.067833848e-12
LI3|_DFF_A|2 I3|_DFF_A|A1 I3|_DFF_A|A2  4.135667696e-12
LI3|_DFF_A|3 I3|_DFF_A|A3 I3|_DFF_A|A4  8.271335392e-12
LI3|_DFF_A|T T03 I3|_DFF_A|T1  2.067833848e-12
LI3|_DFF_A|4 I3|_DFF_A|T1 I3|_DFF_A|T2  4.135667696e-12
LI3|_DFF_A|5 I3|_DFF_A|A4 I3|_DFF_A|Q1  4.135667696e-12
LI3|_DFF_A|6 I3|_DFF_A|Q1 I3|A1_SYNC  2.067833848e-12
LI3|_DFF_B|1 I3|B1 I3|_DFF_B|A1  2.067833848e-12
LI3|_DFF_B|2 I3|_DFF_B|A1 I3|_DFF_B|A2  4.135667696e-12
LI3|_DFF_B|3 I3|_DFF_B|A3 I3|_DFF_B|A4  8.271335392e-12
LI3|_DFF_B|T T03 I3|_DFF_B|T1  2.067833848e-12
LI3|_DFF_B|4 I3|_DFF_B|T1 I3|_DFF_B|T2  4.135667696e-12
LI3|_DFF_B|5 I3|_DFF_B|A4 I3|_DFF_B|Q1  4.135667696e-12
LI3|_DFF_B|6 I3|_DFF_B|Q1 I3|B1_SYNC  2.067833848e-12
LI3|_XOR|A1 I3|A2 I3|_XOR|A1  2.067833848e-12
LI3|_XOR|A2 I3|_XOR|A1 I3|_XOR|A2  4.135667696e-12
LI3|_XOR|A3 I3|_XOR|A3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|B1 I3|B2 I3|_XOR|B1  2.067833848e-12
LI3|_XOR|B2 I3|_XOR|B1 I3|_XOR|B2  4.135667696e-12
LI3|_XOR|B3 I3|_XOR|B3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|T1 T03 I3|_XOR|T1  2.067833848e-12
LI3|_XOR|T2 I3|_XOR|T1 I3|_XOR|T2  4.135667696e-12
LI3|_XOR|Q2 I3|_XOR|ABTQ I3|_XOR|Q1  4.135667696e-12
LI3|_XOR|Q1 I3|_XOR|Q1 IP3_0  2.067833848e-12
LI3|_AND|A1 I3|A1_SYNC I3|_AND|A1  2.067833848e-12
LI3|_AND|A2 I3|_AND|A1 I3|_AND|A2  4.135667696e-12
LI3|_AND|A3 I3|_AND|A3 I3|_AND|Q3  1.2e-12
LI3|_AND|B1 I3|B1_SYNC I3|_AND|B1  2.067833848e-12
LI3|_AND|B2 I3|_AND|B1 I3|_AND|B2  4.135667696e-12
LI3|_AND|B3 I3|_AND|B3 I3|_AND|Q3  1.2e-12
LI3|_AND|Q3 I3|_AND|Q3 I3|_AND|Q2  4.135667696e-12
LI3|_AND|Q2 I3|_AND|Q2 I3|_AND|Q1  4.135667696e-12
LI3|_AND|Q1 I3|_AND|Q1 IG3_0  2.067833848e-12
B_PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP0_0|_TX|B1 0 _PTL_IP0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP0_0|_TX|B2 0 _PTL_IP0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|3  1.684e-12
L_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|6  3.596e-12
L_PTL_IP0_0|_TX|1 IP0_0 _PTL_IP0_0|_TX|1  2.063e-12
L_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|4  4.123e-12
L_PTL_IP0_0|_TX|3 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|7  2.193e-12
R_PTL_IP0_0|_TX|D _PTL_IP0_0|_TX|7 _PTL_IP0_0|A_PTL  1.36
L_PTL_IP0_0|_TX|P1 _PTL_IP0_0|_TX|2 0  5.254e-13
L_PTL_IP0_0|_TX|P2 _PTL_IP0_0|_TX|5 0  5.141e-13
R_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|101  2.7439617672
R_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|104  2.7439617672
L_PTL_IP0_0|_TX|RB1 _PTL_IP0_0|_TX|101 0  1.550338398468e-12
L_PTL_IP0_0|_TX|RB2 _PTL_IP0_0|_TX|104 0  1.550338398468e-12
B_PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP0_0|_RX|B1 0 _PTL_IP0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|3  2.777e-12
I_PTL_IP0_0|_RX|B2 0 _PTL_IP0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|6  2.685e-12
I_PTL_IP0_0|_RX|B3 0 _PTL_IP0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|9  2.764e-12
L_PTL_IP0_0|_RX|1 _PTL_IP0_0|A_PTL _PTL_IP0_0|_RX|1  1.346e-12
L_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|4  6.348e-12
L_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7  5.197e-12
L_PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7 IP0_0_RX  2.058e-12
L_PTL_IP0_0|_RX|P1 _PTL_IP0_0|_RX|2 0  4.795e-13
L_PTL_IP0_0|_RX|P2 _PTL_IP0_0|_RX|5 0  5.431e-13
L_PTL_IP0_0|_RX|P3 _PTL_IP0_0|_RX|8 0  5.339e-13
R_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|101  4.225701121488
R_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|104  3.429952209
R_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|107  2.7439617672
L_PTL_IP0_0|_RX|RB1 _PTL_IP0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP0_0|_RX|RB2 _PTL_IP0_0|_RX|104 0  1.937922998085e-12
L_PTL_IP0_0|_RX|RB3 _PTL_IP0_0|_RX|107 0  1.550338398468e-12
B_PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG0_0|_TX|B1 0 _PTL_IG0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG0_0|_TX|B2 0 _PTL_IG0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|3  1.684e-12
L_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|6  3.596e-12
L_PTL_IG0_0|_TX|1 IG0_0 _PTL_IG0_0|_TX|1  2.063e-12
L_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|4  4.123e-12
L_PTL_IG0_0|_TX|3 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|7  2.193e-12
R_PTL_IG0_0|_TX|D _PTL_IG0_0|_TX|7 _PTL_IG0_0|A_PTL  1.36
L_PTL_IG0_0|_TX|P1 _PTL_IG0_0|_TX|2 0  5.254e-13
L_PTL_IG0_0|_TX|P2 _PTL_IG0_0|_TX|5 0  5.141e-13
R_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|101  2.7439617672
R_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|104  2.7439617672
L_PTL_IG0_0|_TX|RB1 _PTL_IG0_0|_TX|101 0  1.550338398468e-12
L_PTL_IG0_0|_TX|RB2 _PTL_IG0_0|_TX|104 0  1.550338398468e-12
B_PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG0_0|_RX|B1 0 _PTL_IG0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|3  2.777e-12
I_PTL_IG0_0|_RX|B2 0 _PTL_IG0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|6  2.685e-12
I_PTL_IG0_0|_RX|B3 0 _PTL_IG0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|9  2.764e-12
L_PTL_IG0_0|_RX|1 _PTL_IG0_0|A_PTL _PTL_IG0_0|_RX|1  1.346e-12
L_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|4  6.348e-12
L_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7  5.197e-12
L_PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7 IG0_0_RX  2.058e-12
L_PTL_IG0_0|_RX|P1 _PTL_IG0_0|_RX|2 0  4.795e-13
L_PTL_IG0_0|_RX|P2 _PTL_IG0_0|_RX|5 0  5.431e-13
L_PTL_IG0_0|_RX|P3 _PTL_IG0_0|_RX|8 0  5.339e-13
R_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|101  4.225701121488
R_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|104  3.429952209
R_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|107  2.7439617672
L_PTL_IG0_0|_RX|RB1 _PTL_IG0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG0_0|_RX|RB2 _PTL_IG0_0|_RX|104 0  1.937922998085e-12
L_PTL_IG0_0|_RX|RB3 _PTL_IG0_0|_RX|107 0  1.550338398468e-12
B_PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_0|_TX|B1 0 _PTL_IP1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_0|_TX|B2 0 _PTL_IP1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|3  1.684e-12
L_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|6  3.596e-12
L_PTL_IP1_0|_TX|1 IP1_0 _PTL_IP1_0|_TX|1  2.063e-12
L_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|4  4.123e-12
L_PTL_IP1_0|_TX|3 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|7  2.193e-12
R_PTL_IP1_0|_TX|D _PTL_IP1_0|_TX|7 _PTL_IP1_0|A_PTL  1.36
L_PTL_IP1_0|_TX|P1 _PTL_IP1_0|_TX|2 0  5.254e-13
L_PTL_IP1_0|_TX|P2 _PTL_IP1_0|_TX|5 0  5.141e-13
R_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|101  2.7439617672
R_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|104  2.7439617672
L_PTL_IP1_0|_TX|RB1 _PTL_IP1_0|_TX|101 0  1.550338398468e-12
L_PTL_IP1_0|_TX|RB2 _PTL_IP1_0|_TX|104 0  1.550338398468e-12
B_PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_0|_RX|B1 0 _PTL_IP1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|3  2.777e-12
I_PTL_IP1_0|_RX|B2 0 _PTL_IP1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|6  2.685e-12
I_PTL_IP1_0|_RX|B3 0 _PTL_IP1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|9  2.764e-12
L_PTL_IP1_0|_RX|1 _PTL_IP1_0|A_PTL _PTL_IP1_0|_RX|1  1.346e-12
L_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|4  6.348e-12
L_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7  5.197e-12
L_PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7 IP1_0_RX  2.058e-12
L_PTL_IP1_0|_RX|P1 _PTL_IP1_0|_RX|2 0  4.795e-13
L_PTL_IP1_0|_RX|P2 _PTL_IP1_0|_RX|5 0  5.431e-13
L_PTL_IP1_0|_RX|P3 _PTL_IP1_0|_RX|8 0  5.339e-13
R_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|101  4.225701121488
R_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|104  3.429952209
R_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|107  2.7439617672
L_PTL_IP1_0|_RX|RB1 _PTL_IP1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_0|_RX|RB2 _PTL_IP1_0|_RX|104 0  1.937922998085e-12
L_PTL_IP1_0|_RX|RB3 _PTL_IP1_0|_RX|107 0  1.550338398468e-12
B_PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG1_0|_TX|B1 0 _PTL_IG1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG1_0|_TX|B2 0 _PTL_IG1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|3  1.684e-12
L_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|6  3.596e-12
L_PTL_IG1_0|_TX|1 IG1_0 _PTL_IG1_0|_TX|1  2.063e-12
L_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|4  4.123e-12
L_PTL_IG1_0|_TX|3 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|7  2.193e-12
R_PTL_IG1_0|_TX|D _PTL_IG1_0|_TX|7 _PTL_IG1_0|A_PTL  1.36
L_PTL_IG1_0|_TX|P1 _PTL_IG1_0|_TX|2 0  5.254e-13
L_PTL_IG1_0|_TX|P2 _PTL_IG1_0|_TX|5 0  5.141e-13
R_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|101  2.7439617672
R_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|104  2.7439617672
L_PTL_IG1_0|_TX|RB1 _PTL_IG1_0|_TX|101 0  1.550338398468e-12
L_PTL_IG1_0|_TX|RB2 _PTL_IG1_0|_TX|104 0  1.550338398468e-12
B_PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG1_0|_RX|B1 0 _PTL_IG1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|3  2.777e-12
I_PTL_IG1_0|_RX|B2 0 _PTL_IG1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|6  2.685e-12
I_PTL_IG1_0|_RX|B3 0 _PTL_IG1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|9  2.764e-12
L_PTL_IG1_0|_RX|1 _PTL_IG1_0|A_PTL _PTL_IG1_0|_RX|1  1.346e-12
L_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|4  6.348e-12
L_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7  5.197e-12
L_PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7 IG1_0_RX  2.058e-12
L_PTL_IG1_0|_RX|P1 _PTL_IG1_0|_RX|2 0  4.795e-13
L_PTL_IG1_0|_RX|P2 _PTL_IG1_0|_RX|5 0  5.431e-13
L_PTL_IG1_0|_RX|P3 _PTL_IG1_0|_RX|8 0  5.339e-13
R_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|101  4.225701121488
R_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|104  3.429952209
R_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|107  2.7439617672
L_PTL_IG1_0|_RX|RB1 _PTL_IG1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG1_0|_RX|RB2 _PTL_IG1_0|_RX|104 0  1.937922998085e-12
L_PTL_IG1_0|_RX|RB3 _PTL_IG1_0|_RX|107 0  1.550338398468e-12
B_PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_0|_TX|B1 0 _PTL_IP2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_0|_TX|B2 0 _PTL_IP2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|3  1.684e-12
L_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|6  3.596e-12
L_PTL_IP2_0|_TX|1 IP2_0 _PTL_IP2_0|_TX|1  2.063e-12
L_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|4  4.123e-12
L_PTL_IP2_0|_TX|3 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|7  2.193e-12
R_PTL_IP2_0|_TX|D _PTL_IP2_0|_TX|7 _PTL_IP2_0|A_PTL  1.36
L_PTL_IP2_0|_TX|P1 _PTL_IP2_0|_TX|2 0  5.254e-13
L_PTL_IP2_0|_TX|P2 _PTL_IP2_0|_TX|5 0  5.141e-13
R_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|101  2.7439617672
R_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|104  2.7439617672
L_PTL_IP2_0|_TX|RB1 _PTL_IP2_0|_TX|101 0  1.550338398468e-12
L_PTL_IP2_0|_TX|RB2 _PTL_IP2_0|_TX|104 0  1.550338398468e-12
B_PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_0|_RX|B1 0 _PTL_IP2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|3  2.777e-12
I_PTL_IP2_0|_RX|B2 0 _PTL_IP2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|6  2.685e-12
I_PTL_IP2_0|_RX|B3 0 _PTL_IP2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|9  2.764e-12
L_PTL_IP2_0|_RX|1 _PTL_IP2_0|A_PTL _PTL_IP2_0|_RX|1  1.346e-12
L_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|4  6.348e-12
L_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7  5.197e-12
L_PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7 IP2_0_RX  2.058e-12
L_PTL_IP2_0|_RX|P1 _PTL_IP2_0|_RX|2 0  4.795e-13
L_PTL_IP2_0|_RX|P2 _PTL_IP2_0|_RX|5 0  5.431e-13
L_PTL_IP2_0|_RX|P3 _PTL_IP2_0|_RX|8 0  5.339e-13
R_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|101  4.225701121488
R_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|104  3.429952209
R_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|107  2.7439617672
L_PTL_IP2_0|_RX|RB1 _PTL_IP2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_0|_RX|RB2 _PTL_IP2_0|_RX|104 0  1.937922998085e-12
L_PTL_IP2_0|_RX|RB3 _PTL_IP2_0|_RX|107 0  1.550338398468e-12
B_PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG2_0|_TX|B1 0 _PTL_IG2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG2_0|_TX|B2 0 _PTL_IG2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|3  1.684e-12
L_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|6  3.596e-12
L_PTL_IG2_0|_TX|1 IG2_0 _PTL_IG2_0|_TX|1  2.063e-12
L_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|4  4.123e-12
L_PTL_IG2_0|_TX|3 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|7  2.193e-12
R_PTL_IG2_0|_TX|D _PTL_IG2_0|_TX|7 _PTL_IG2_0|A_PTL  1.36
L_PTL_IG2_0|_TX|P1 _PTL_IG2_0|_TX|2 0  5.254e-13
L_PTL_IG2_0|_TX|P2 _PTL_IG2_0|_TX|5 0  5.141e-13
R_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|101  2.7439617672
R_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|104  2.7439617672
L_PTL_IG2_0|_TX|RB1 _PTL_IG2_0|_TX|101 0  1.550338398468e-12
L_PTL_IG2_0|_TX|RB2 _PTL_IG2_0|_TX|104 0  1.550338398468e-12
B_PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG2_0|_RX|B1 0 _PTL_IG2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|3  2.777e-12
I_PTL_IG2_0|_RX|B2 0 _PTL_IG2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|6  2.685e-12
I_PTL_IG2_0|_RX|B3 0 _PTL_IG2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|9  2.764e-12
L_PTL_IG2_0|_RX|1 _PTL_IG2_0|A_PTL _PTL_IG2_0|_RX|1  1.346e-12
L_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|4  6.348e-12
L_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7  5.197e-12
L_PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7 IG2_0_RX  2.058e-12
L_PTL_IG2_0|_RX|P1 _PTL_IG2_0|_RX|2 0  4.795e-13
L_PTL_IG2_0|_RX|P2 _PTL_IG2_0|_RX|5 0  5.431e-13
L_PTL_IG2_0|_RX|P3 _PTL_IG2_0|_RX|8 0  5.339e-13
R_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|101  4.225701121488
R_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|104  3.429952209
R_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|107  2.7439617672
L_PTL_IG2_0|_RX|RB1 _PTL_IG2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG2_0|_RX|RB2 _PTL_IG2_0|_RX|104 0  1.937922998085e-12
L_PTL_IG2_0|_RX|RB3 _PTL_IG2_0|_RX|107 0  1.550338398468e-12
B_PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_0|_TX|B1 0 _PTL_IP3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_0|_TX|B2 0 _PTL_IP3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|3  1.684e-12
L_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|6  3.596e-12
L_PTL_IP3_0|_TX|1 IP3_0 _PTL_IP3_0|_TX|1  2.063e-12
L_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|4  4.123e-12
L_PTL_IP3_0|_TX|3 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|7  2.193e-12
R_PTL_IP3_0|_TX|D _PTL_IP3_0|_TX|7 _PTL_IP3_0|A_PTL  1.36
L_PTL_IP3_0|_TX|P1 _PTL_IP3_0|_TX|2 0  5.254e-13
L_PTL_IP3_0|_TX|P2 _PTL_IP3_0|_TX|5 0  5.141e-13
R_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|101  2.7439617672
R_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|104  2.7439617672
L_PTL_IP3_0|_TX|RB1 _PTL_IP3_0|_TX|101 0  1.550338398468e-12
L_PTL_IP3_0|_TX|RB2 _PTL_IP3_0|_TX|104 0  1.550338398468e-12
B_PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_0|_RX|B1 0 _PTL_IP3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|3  2.777e-12
I_PTL_IP3_0|_RX|B2 0 _PTL_IP3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|6  2.685e-12
I_PTL_IP3_0|_RX|B3 0 _PTL_IP3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|9  2.764e-12
L_PTL_IP3_0|_RX|1 _PTL_IP3_0|A_PTL _PTL_IP3_0|_RX|1  1.346e-12
L_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|4  6.348e-12
L_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7  5.197e-12
L_PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7 IP3_0_RX  2.058e-12
L_PTL_IP3_0|_RX|P1 _PTL_IP3_0|_RX|2 0  4.795e-13
L_PTL_IP3_0|_RX|P2 _PTL_IP3_0|_RX|5 0  5.431e-13
L_PTL_IP3_0|_RX|P3 _PTL_IP3_0|_RX|8 0  5.339e-13
R_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|101  4.225701121488
R_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|104  3.429952209
R_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|107  2.7439617672
L_PTL_IP3_0|_RX|RB1 _PTL_IP3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_0|_RX|RB2 _PTL_IP3_0|_RX|104 0  1.937922998085e-12
L_PTL_IP3_0|_RX|RB3 _PTL_IP3_0|_RX|107 0  1.550338398468e-12
B_PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG3_0|_TX|B1 0 _PTL_IG3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG3_0|_TX|B2 0 _PTL_IG3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|3  1.684e-12
L_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|6  3.596e-12
L_PTL_IG3_0|_TX|1 IG3_0 _PTL_IG3_0|_TX|1  2.063e-12
L_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|4  4.123e-12
L_PTL_IG3_0|_TX|3 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|7  2.193e-12
R_PTL_IG3_0|_TX|D _PTL_IG3_0|_TX|7 _PTL_IG3_0|A_PTL  1.36
L_PTL_IG3_0|_TX|P1 _PTL_IG3_0|_TX|2 0  5.254e-13
L_PTL_IG3_0|_TX|P2 _PTL_IG3_0|_TX|5 0  5.141e-13
R_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|101  2.7439617672
R_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|104  2.7439617672
L_PTL_IG3_0|_TX|RB1 _PTL_IG3_0|_TX|101 0  1.550338398468e-12
L_PTL_IG3_0|_TX|RB2 _PTL_IG3_0|_TX|104 0  1.550338398468e-12
B_PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG3_0|_RX|B1 0 _PTL_IG3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|3  2.777e-12
I_PTL_IG3_0|_RX|B2 0 _PTL_IG3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|6  2.685e-12
I_PTL_IG3_0|_RX|B3 0 _PTL_IG3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|9  2.764e-12
L_PTL_IG3_0|_RX|1 _PTL_IG3_0|A_PTL _PTL_IG3_0|_RX|1  1.346e-12
L_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|4  6.348e-12
L_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7  5.197e-12
L_PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7 IG3_0_RX  2.058e-12
L_PTL_IG3_0|_RX|P1 _PTL_IG3_0|_RX|2 0  4.795e-13
L_PTL_IG3_0|_RX|P2 _PTL_IG3_0|_RX|5 0  5.431e-13
L_PTL_IG3_0|_RX|P3 _PTL_IG3_0|_RX|8 0  5.339e-13
R_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|101  4.225701121488
R_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|104  3.429952209
R_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|107  2.7439617672
L_PTL_IG3_0|_RX|RB1 _PTL_IG3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG3_0|_RX|RB2 _PTL_IG3_0|_RX|104 0  1.937922998085e-12
L_PTL_IG3_0|_RX|RB3 _PTL_IG3_0|_RX|107 0  1.550338398468e-12
LSPL_IG0_0|I_D1|B SPL_IG0_0|D1 SPL_IG0_0|I_D1|MID  2e-12
ISPL_IG0_0|I_D1|B 0 SPL_IG0_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_D2|B SPL_IG0_0|D2 SPL_IG0_0|I_D2|MID  2e-12
ISPL_IG0_0|I_D2|B 0 SPL_IG0_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG0_0|I_Q1|B SPL_IG0_0|QA1 SPL_IG0_0|I_Q1|MID  2e-12
ISPL_IG0_0|I_Q1|B 0 SPL_IG0_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_Q2|B SPL_IG0_0|QB1 SPL_IG0_0|I_Q2|MID  2e-12
ISPL_IG0_0|I_Q2|B 0 SPL_IG0_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG0_0|1|1 SPL_IG0_0|D1 SPL_IG0_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|1|P SPL_IG0_0|1|MID_SERIES 0  2e-13
RSPL_IG0_0|1|B SPL_IG0_0|D1 SPL_IG0_0|1|MID_SHUNT  2.7439617672
LSPL_IG0_0|1|RB SPL_IG0_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|2|1 SPL_IG0_0|D2 SPL_IG0_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|2|P SPL_IG0_0|2|MID_SERIES 0  2e-13
RSPL_IG0_0|2|B SPL_IG0_0|D2 SPL_IG0_0|2|MID_SHUNT  2.7439617672
LSPL_IG0_0|2|RB SPL_IG0_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|A|1 SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|A|P SPL_IG0_0|A|MID_SERIES 0  2e-13
RSPL_IG0_0|A|B SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SHUNT  2.7439617672
LSPL_IG0_0|A|RB SPL_IG0_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|B|1 SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|B|P SPL_IG0_0|B|MID_SERIES 0  2e-13
RSPL_IG0_0|B|B SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SHUNT  2.7439617672
LSPL_IG0_0|B|RB SPL_IG0_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP1_0|I_D1|B SPL_IP1_0|D1 SPL_IP1_0|I_D1|MID  2e-12
ISPL_IP1_0|I_D1|B 0 SPL_IP1_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_D2|B SPL_IP1_0|D2 SPL_IP1_0|I_D2|MID  2e-12
ISPL_IP1_0|I_D2|B 0 SPL_IP1_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP1_0|I_Q1|B SPL_IP1_0|QA1 SPL_IP1_0|I_Q1|MID  2e-12
ISPL_IP1_0|I_Q1|B 0 SPL_IP1_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_Q2|B SPL_IP1_0|QB1 SPL_IP1_0|I_Q2|MID  2e-12
ISPL_IP1_0|I_Q2|B 0 SPL_IP1_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP1_0|1|1 SPL_IP1_0|D1 SPL_IP1_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|1|P SPL_IP1_0|1|MID_SERIES 0  2e-13
RSPL_IP1_0|1|B SPL_IP1_0|D1 SPL_IP1_0|1|MID_SHUNT  2.7439617672
LSPL_IP1_0|1|RB SPL_IP1_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|2|1 SPL_IP1_0|D2 SPL_IP1_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|2|P SPL_IP1_0|2|MID_SERIES 0  2e-13
RSPL_IP1_0|2|B SPL_IP1_0|D2 SPL_IP1_0|2|MID_SHUNT  2.7439617672
LSPL_IP1_0|2|RB SPL_IP1_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|A|1 SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|A|P SPL_IP1_0|A|MID_SERIES 0  2e-13
RSPL_IP1_0|A|B SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SHUNT  2.7439617672
LSPL_IP1_0|A|RB SPL_IP1_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|B|1 SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|B|P SPL_IP1_0|B|MID_SERIES 0  2e-13
RSPL_IP1_0|B|B SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SHUNT  2.7439617672
LSPL_IP1_0|B|RB SPL_IP1_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|1 IP2_0_RX SPL_IP2_0|SPL1|D1  2e-12
LSPL_IP2_0|SPL1|2 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|D2  4.135667696e-12
LSPL_IP2_0|SPL1|3 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL1|4 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL1|5 SPL_IP2_0|SPL1|QA1 IP2_0_TO2  2e-12
LSPL_IP2_0|SPL1|6 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL1|7 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|QTMP  2e-12
LSPL_IP2_0|SPL2|1 SPL_IP2_0|QTMP SPL_IP2_0|SPL2|D1  2e-12
LSPL_IP2_0|SPL2|2 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|D2  4.135667696e-12
LSPL_IP2_0|SPL2|3 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL2|4 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL2|5 SPL_IP2_0|SPL2|QA1 IP2_0_TO3  2e-12
LSPL_IP2_0|SPL2|6 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL2|7 SPL_IP2_0|SPL2|QB1 IP2_0_OUT  2e-12
LSPL_IG2_0|I_D1|B SPL_IG2_0|D1 SPL_IG2_0|I_D1|MID  2e-12
ISPL_IG2_0|I_D1|B 0 SPL_IG2_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_D2|B SPL_IG2_0|D2 SPL_IG2_0|I_D2|MID  2e-12
ISPL_IG2_0|I_D2|B 0 SPL_IG2_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG2_0|I_Q1|B SPL_IG2_0|QA1 SPL_IG2_0|I_Q1|MID  2e-12
ISPL_IG2_0|I_Q1|B 0 SPL_IG2_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_Q2|B SPL_IG2_0|QB1 SPL_IG2_0|I_Q2|MID  2e-12
ISPL_IG2_0|I_Q2|B 0 SPL_IG2_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG2_0|1|1 SPL_IG2_0|D1 SPL_IG2_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|1|P SPL_IG2_0|1|MID_SERIES 0  2e-13
RSPL_IG2_0|1|B SPL_IG2_0|D1 SPL_IG2_0|1|MID_SHUNT  2.7439617672
LSPL_IG2_0|1|RB SPL_IG2_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|2|1 SPL_IG2_0|D2 SPL_IG2_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|2|P SPL_IG2_0|2|MID_SERIES 0  2e-13
RSPL_IG2_0|2|B SPL_IG2_0|D2 SPL_IG2_0|2|MID_SHUNT  2.7439617672
LSPL_IG2_0|2|RB SPL_IG2_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|A|1 SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|A|P SPL_IG2_0|A|MID_SERIES 0  2e-13
RSPL_IG2_0|A|B SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SHUNT  2.7439617672
LSPL_IG2_0|A|RB SPL_IG2_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|B|1 SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|B|P SPL_IG2_0|B|MID_SERIES 0  2e-13
RSPL_IG2_0|B|B SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SHUNT  2.7439617672
LSPL_IG2_0|B|RB SPL_IG2_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP3_0|I_D1|B SPL_IP3_0|D1 SPL_IP3_0|I_D1|MID  2e-12
ISPL_IP3_0|I_D1|B 0 SPL_IP3_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_D2|B SPL_IP3_0|D2 SPL_IP3_0|I_D2|MID  2e-12
ISPL_IP3_0|I_D2|B 0 SPL_IP3_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP3_0|I_Q1|B SPL_IP3_0|QA1 SPL_IP3_0|I_Q1|MID  2e-12
ISPL_IP3_0|I_Q1|B 0 SPL_IP3_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_Q2|B SPL_IP3_0|QB1 SPL_IP3_0|I_Q2|MID  2e-12
ISPL_IP3_0|I_Q2|B 0 SPL_IP3_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP3_0|1|1 SPL_IP3_0|D1 SPL_IP3_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|1|P SPL_IP3_0|1|MID_SERIES 0  2e-13
RSPL_IP3_0|1|B SPL_IP3_0|D1 SPL_IP3_0|1|MID_SHUNT  2.7439617672
LSPL_IP3_0|1|RB SPL_IP3_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|2|1 SPL_IP3_0|D2 SPL_IP3_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|2|P SPL_IP3_0|2|MID_SERIES 0  2e-13
RSPL_IP3_0|2|B SPL_IP3_0|D2 SPL_IP3_0|2|MID_SHUNT  2.7439617672
LSPL_IP3_0|2|RB SPL_IP3_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|A|1 SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|A|P SPL_IP3_0|A|MID_SERIES 0  2e-13
RSPL_IP3_0|A|B SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SHUNT  2.7439617672
LSPL_IP3_0|A|RB SPL_IP3_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|B|1 SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|B|P SPL_IP3_0|B|MID_SERIES 0  2e-13
RSPL_IP3_0|B|B SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SHUNT  2.7439617672
LSPL_IP3_0|B|RB SPL_IP3_0|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|1 IP0_0_RX _PG0_01|P|A1  2.067833848e-12
L_PG0_01|P|2 _PG0_01|P|A1 _PG0_01|P|A2  4.135667696e-12
L_PG0_01|P|3 _PG0_01|P|A3 _PG0_01|P|A4  8.271335392e-12
L_PG0_01|P|T T04 _PG0_01|P|T1  2.067833848e-12
L_PG0_01|P|4 _PG0_01|P|T1 _PG0_01|P|T2  4.135667696e-12
L_PG0_01|P|5 _PG0_01|P|A4 _PG0_01|P|Q1  4.135667696e-12
L_PG0_01|P|6 _PG0_01|P|Q1 P0_1  2.067833848e-12
L_PG0_01|G|1 IG0_0_TO0 _PG0_01|G|A1  2.067833848e-12
L_PG0_01|G|2 _PG0_01|G|A1 _PG0_01|G|A2  4.135667696e-12
L_PG0_01|G|3 _PG0_01|G|A3 _PG0_01|G|A4  8.271335392e-12
L_PG0_01|G|T T04 _PG0_01|G|T1  2.067833848e-12
L_PG0_01|G|4 _PG0_01|G|T1 _PG0_01|G|T2  4.135667696e-12
L_PG0_01|G|5 _PG0_01|G|A4 _PG0_01|G|Q1  4.135667696e-12
L_PG0_01|G|6 _PG0_01|G|Q1 G0_1  2.067833848e-12
L_PG1_01|_SPL_G1|1 IG1_0_RX _PG1_01|_SPL_G1|D1  2e-12
L_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|D2  4.135667696e-12
L_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG1_01|_SPL_G1|5 _PG1_01|_SPL_G1|QA1 _PG1_01|G1_COPY_1  2e-12
L_PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|QB1 _PG1_01|G1_COPY_2  2e-12
L_PG1_01|_PG|A1 IP1_0_TO1 _PG1_01|_PG|A1  2.067833848e-12
L_PG1_01|_PG|A2 _PG1_01|_PG|A1 _PG1_01|_PG|A2  4.135667696e-12
L_PG1_01|_PG|A3 _PG1_01|_PG|A3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|B1 _PG1_01|G1_COPY_1 _PG1_01|_PG|B1  2.067833848e-12
L_PG1_01|_PG|B2 _PG1_01|_PG|B1 _PG1_01|_PG|B2  4.135667696e-12
L_PG1_01|_PG|B3 _PG1_01|_PG|B3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|Q3 _PG1_01|_PG|Q3 _PG1_01|_PG|Q2  4.135667696e-12
L_PG1_01|_PG|Q2 _PG1_01|_PG|Q2 _PG1_01|_PG|Q1  4.135667696e-12
L_PG1_01|_PG|Q1 _PG1_01|_PG|Q1 _PG1_01|PG  2.067833848e-12
L_PG1_01|_GG|A1 IG0_0_TO1 _PG1_01|_GG|A1  2.067833848e-12
L_PG1_01|_GG|A2 _PG1_01|_GG|A1 _PG1_01|_GG|A2  4.135667696e-12
L_PG1_01|_GG|A3 _PG1_01|_GG|A3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|B1 _PG1_01|G1_COPY_2 _PG1_01|_GG|B1  2.067833848e-12
L_PG1_01|_GG|B2 _PG1_01|_GG|B1 _PG1_01|_GG|B2  4.135667696e-12
L_PG1_01|_GG|B3 _PG1_01|_GG|B3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|Q3 _PG1_01|_GG|Q3 _PG1_01|_GG|Q2  4.135667696e-12
L_PG1_01|_GG|Q2 _PG1_01|_GG|Q2 _PG1_01|_GG|Q1  4.135667696e-12
L_PG1_01|_GG|Q1 _PG1_01|_GG|Q1 _PG1_01|GG  2.067833848e-12
L_PG1_01|_DFF_PG|1 _PG1_01|PG _PG1_01|_DFF_PG|A1  2.067833848e-12
L_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|A2  4.135667696e-12
L_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|A4  8.271335392e-12
L_PG1_01|_DFF_PG|T T05 _PG1_01|_DFF_PG|T1  2.067833848e-12
L_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T2  4.135667696e-12
L_PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|Q1  4.135667696e-12
L_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|Q1 _PG1_01|PG_SYNC  2.067833848e-12
L_PG1_01|_DFF_GG|1 _PG1_01|GG _PG1_01|_DFF_GG|A1  2.067833848e-12
L_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|A2  4.135667696e-12
L_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|A4  8.271335392e-12
L_PG1_01|_DFF_GG|T T05 _PG1_01|_DFF_GG|T1  2.067833848e-12
L_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T2  4.135667696e-12
L_PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|Q1  4.135667696e-12
L_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|Q1 _PG1_01|GG_SYNC  2.067833848e-12
L_PG1_01|_AND_G|A1 _PG1_01|PG_SYNC _PG1_01|_AND_G|A1  2.067833848e-12
L_PG1_01|_AND_G|A2 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A2  4.135667696e-12
L_PG1_01|_AND_G|A3 _PG1_01|_AND_G|A3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|B1 _PG1_01|GG_SYNC _PG1_01|_AND_G|B1  2.067833848e-12
L_PG1_01|_AND_G|B2 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B2  4.135667696e-12
L_PG1_01|_AND_G|B3 _PG1_01|_AND_G|B3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q2  4.135667696e-12
L_PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q1  4.135667696e-12
L_PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1 G1_1  2.067833848e-12
L_PG2_01|P|1 IP2_0_TO2 _PG2_01|P|A1  2.067833848e-12
L_PG2_01|P|2 _PG2_01|P|A1 _PG2_01|P|A2  4.135667696e-12
L_PG2_01|P|3 _PG2_01|P|A3 _PG2_01|P|A4  8.271335392e-12
L_PG2_01|P|T T06 _PG2_01|P|T1  2.067833848e-12
L_PG2_01|P|4 _PG2_01|P|T1 _PG2_01|P|T2  4.135667696e-12
L_PG2_01|P|5 _PG2_01|P|A4 _PG2_01|P|Q1  4.135667696e-12
L_PG2_01|P|6 _PG2_01|P|Q1 P2_1  2.067833848e-12
L_PG2_01|G|1 IG2_0_TO2 _PG2_01|G|A1  2.067833848e-12
L_PG2_01|G|2 _PG2_01|G|A1 _PG2_01|G|A2  4.135667696e-12
L_PG2_01|G|3 _PG2_01|G|A3 _PG2_01|G|A4  8.271335392e-12
L_PG2_01|G|T T06 _PG2_01|G|T1  2.067833848e-12
L_PG2_01|G|4 _PG2_01|G|T1 _PG2_01|G|T2  4.135667696e-12
L_PG2_01|G|5 _PG2_01|G|A4 _PG2_01|G|Q1  4.135667696e-12
L_PG2_01|G|6 _PG2_01|G|Q1 G2_1  2.067833848e-12
L_PG3_01|_SPL_G1|1 IG3_0_RX _PG3_01|_SPL_G1|D1  2e-12
L_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|D2  4.135667696e-12
L_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_G1|5 _PG3_01|_SPL_G1|QA1 _PG3_01|G1_COPY_1  2e-12
L_PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|QB1 _PG3_01|G1_COPY_2  2e-12
L_PG3_01|_SPL_P1|1 IP3_0_TO1 _PG3_01|_SPL_P1|D1  2e-12
L_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|D2  4.135667696e-12
L_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_P1|5 _PG3_01|_SPL_P1|QA1 _PG3_01|P1_COPY_1  2e-12
L_PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|QB1 _PG3_01|P1_COPY_2  2e-12
L_PG3_01|_PG|A1 _PG3_01|P1_COPY_1 _PG3_01|_PG|A1  2.067833848e-12
L_PG3_01|_PG|A2 _PG3_01|_PG|A1 _PG3_01|_PG|A2  4.135667696e-12
L_PG3_01|_PG|A3 _PG3_01|_PG|A3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|B1 _PG3_01|G1_COPY_1 _PG3_01|_PG|B1  2.067833848e-12
L_PG3_01|_PG|B2 _PG3_01|_PG|B1 _PG3_01|_PG|B2  4.135667696e-12
L_PG3_01|_PG|B3 _PG3_01|_PG|B3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|Q3 _PG3_01|_PG|Q3 _PG3_01|_PG|Q2  4.135667696e-12
L_PG3_01|_PG|Q2 _PG3_01|_PG|Q2 _PG3_01|_PG|Q1  4.135667696e-12
L_PG3_01|_PG|Q1 _PG3_01|_PG|Q1 _PG3_01|PG  2.067833848e-12
L_PG3_01|_GG|A1 IG2_0_TO3 _PG3_01|_GG|A1  2.067833848e-12
L_PG3_01|_GG|A2 _PG3_01|_GG|A1 _PG3_01|_GG|A2  4.135667696e-12
L_PG3_01|_GG|A3 _PG3_01|_GG|A3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|B1 _PG3_01|G1_COPY_2 _PG3_01|_GG|B1  2.067833848e-12
L_PG3_01|_GG|B2 _PG3_01|_GG|B1 _PG3_01|_GG|B2  4.135667696e-12
L_PG3_01|_GG|B3 _PG3_01|_GG|B3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|Q3 _PG3_01|_GG|Q3 _PG3_01|_GG|Q2  4.135667696e-12
L_PG3_01|_GG|Q2 _PG3_01|_GG|Q2 _PG3_01|_GG|Q1  4.135667696e-12
L_PG3_01|_GG|Q1 _PG3_01|_GG|Q1 _PG3_01|GG  2.067833848e-12
L_PG3_01|_DFF_P0|1 IP2_0_TO3 _PG3_01|_DFF_P0|A1  2.067833848e-12
L_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|A2  4.135667696e-12
L_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|A4  8.271335392e-12
L_PG3_01|_DFF_P0|T T07 _PG3_01|_DFF_P0|T1  2.067833848e-12
L_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T2  4.135667696e-12
L_PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|Q1  4.135667696e-12
L_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|Q1 _PG3_01|P0_SYNC  2.067833848e-12
L_PG3_01|_DFF_P1|1 _PG3_01|P1_COPY_2 _PG3_01|_DFF_P1|A1  2.067833848e-12
L_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|A2  4.135667696e-12
L_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|A4  8.271335392e-12
L_PG3_01|_DFF_P1|T T07 _PG3_01|_DFF_P1|T1  2.067833848e-12
L_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T2  4.135667696e-12
L_PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|Q1  4.135667696e-12
L_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|Q1 _PG3_01|P1_SYNC  2.067833848e-12
L_PG3_01|_DFF_PG|1 _PG3_01|PG _PG3_01|_DFF_PG|A1  2.067833848e-12
L_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|A2  4.135667696e-12
L_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|A4  8.271335392e-12
L_PG3_01|_DFF_PG|T T07 _PG3_01|_DFF_PG|T1  2.067833848e-12
L_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T2  4.135667696e-12
L_PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|Q1  4.135667696e-12
L_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|Q1 _PG3_01|PG_SYNC  2.067833848e-12
L_PG3_01|_DFF_GG|1 _PG3_01|GG _PG3_01|_DFF_GG|A1  2.067833848e-12
L_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|A2  4.135667696e-12
L_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|A4  8.271335392e-12
L_PG3_01|_DFF_GG|T T07 _PG3_01|_DFF_GG|T1  2.067833848e-12
L_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T2  4.135667696e-12
L_PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|Q1  4.135667696e-12
L_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|Q1 _PG3_01|GG_SYNC  2.067833848e-12
L_PG3_01|_AND_G|A1 _PG3_01|PG_SYNC _PG3_01|_AND_G|A1  2.067833848e-12
L_PG3_01|_AND_G|A2 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A2  4.135667696e-12
L_PG3_01|_AND_G|A3 _PG3_01|_AND_G|A3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|B1 _PG3_01|GG_SYNC _PG3_01|_AND_G|B1  2.067833848e-12
L_PG3_01|_AND_G|B2 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B2  4.135667696e-12
L_PG3_01|_AND_G|B3 _PG3_01|_AND_G|B3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q2  4.135667696e-12
L_PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q1  4.135667696e-12
L_PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1 G3_1  2.067833848e-12
L_PG3_01|_AND_P|A1 _PG3_01|P0_SYNC _PG3_01|_AND_P|A1  2.067833848e-12
L_PG3_01|_AND_P|A2 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A2  4.135667696e-12
L_PG3_01|_AND_P|A3 _PG3_01|_AND_P|A3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|B1 _PG3_01|P1_SYNC _PG3_01|_AND_P|B1  2.067833848e-12
L_PG3_01|_AND_P|B2 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B2  4.135667696e-12
L_PG3_01|_AND_P|B3 _PG3_01|_AND_P|B3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q2  4.135667696e-12
L_PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q1  4.135667696e-12
L_PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1 P3_1  2.067833848e-12
L_DFF_IP1_01|I_1|B _DFF_IP1_01|A1 _DFF_IP1_01|I_1|MID  2e-12
I_DFF_IP1_01|I_1|B 0 _DFF_IP1_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_3|B _DFF_IP1_01|A3 _DFF_IP1_01|I_3|MID  2e-12
I_DFF_IP1_01|I_3|B 0 _DFF_IP1_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_01|I_T|B _DFF_IP1_01|T1 _DFF_IP1_01|I_T|MID  2e-12
I_DFF_IP1_01|I_T|B 0 _DFF_IP1_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_6|B _DFF_IP1_01|Q1 _DFF_IP1_01|I_6|MID  2e-12
I_DFF_IP1_01|I_6|B 0 _DFF_IP1_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_01|1|1 _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|1|P _DFF_IP1_01|1|MID_SERIES 0  2e-13
R_DFF_IP1_01|1|B _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SHUNT  2.7439617672
L_DFF_IP1_01|1|RB _DFF_IP1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|23|1 _DFF_IP1_01|A2 _DFF_IP1_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|23|B _DFF_IP1_01|A2 _DFF_IP1_01|23|MID_SHUNT  3.84154647408
L_DFF_IP1_01|23|RB _DFF_IP1_01|23|MID_SHUNT _DFF_IP1_01|A3  2.1704737578552e-12
B_DFF_IP1_01|3|1 _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|3|P _DFF_IP1_01|3|MID_SERIES 0  2e-13
R_DFF_IP1_01|3|B _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SHUNT  2.7439617672
L_DFF_IP1_01|3|RB _DFF_IP1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|4|1 _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|4|P _DFF_IP1_01|4|MID_SERIES 0  2e-13
R_DFF_IP1_01|4|B _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SHUNT  2.7439617672
L_DFF_IP1_01|4|RB _DFF_IP1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|T|1 _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|T|P _DFF_IP1_01|T|MID_SERIES 0  2e-13
R_DFF_IP1_01|T|B _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SHUNT  2.7439617672
L_DFF_IP1_01|T|RB _DFF_IP1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|45|1 _DFF_IP1_01|T2 _DFF_IP1_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|45|B _DFF_IP1_01|T2 _DFF_IP1_01|45|MID_SHUNT  3.84154647408
L_DFF_IP1_01|45|RB _DFF_IP1_01|45|MID_SHUNT _DFF_IP1_01|A4  2.1704737578552e-12
B_DFF_IP1_01|6|1 _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|6|P _DFF_IP1_01|6|MID_SERIES 0  2e-13
R_DFF_IP1_01|6|B _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SHUNT  2.7439617672
L_DFF_IP1_01|6|RB _DFF_IP1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_01|I_1|B _DFF_IP2_01|A1 _DFF_IP2_01|I_1|MID  2e-12
I_DFF_IP2_01|I_1|B 0 _DFF_IP2_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_3|B _DFF_IP2_01|A3 _DFF_IP2_01|I_3|MID  2e-12
I_DFF_IP2_01|I_3|B 0 _DFF_IP2_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_01|I_T|B _DFF_IP2_01|T1 _DFF_IP2_01|I_T|MID  2e-12
I_DFF_IP2_01|I_T|B 0 _DFF_IP2_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_6|B _DFF_IP2_01|Q1 _DFF_IP2_01|I_6|MID  2e-12
I_DFF_IP2_01|I_6|B 0 _DFF_IP2_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_01|1|1 _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|1|P _DFF_IP2_01|1|MID_SERIES 0  2e-13
R_DFF_IP2_01|1|B _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SHUNT  2.7439617672
L_DFF_IP2_01|1|RB _DFF_IP2_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|23|1 _DFF_IP2_01|A2 _DFF_IP2_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|23|B _DFF_IP2_01|A2 _DFF_IP2_01|23|MID_SHUNT  3.84154647408
L_DFF_IP2_01|23|RB _DFF_IP2_01|23|MID_SHUNT _DFF_IP2_01|A3  2.1704737578552e-12
B_DFF_IP2_01|3|1 _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|3|P _DFF_IP2_01|3|MID_SERIES 0  2e-13
R_DFF_IP2_01|3|B _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SHUNT  2.7439617672
L_DFF_IP2_01|3|RB _DFF_IP2_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|4|1 _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|4|P _DFF_IP2_01|4|MID_SERIES 0  2e-13
R_DFF_IP2_01|4|B _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SHUNT  2.7439617672
L_DFF_IP2_01|4|RB _DFF_IP2_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|T|1 _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|T|P _DFF_IP2_01|T|MID_SERIES 0  2e-13
R_DFF_IP2_01|T|B _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SHUNT  2.7439617672
L_DFF_IP2_01|T|RB _DFF_IP2_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|45|1 _DFF_IP2_01|T2 _DFF_IP2_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|45|B _DFF_IP2_01|T2 _DFF_IP2_01|45|MID_SHUNT  3.84154647408
L_DFF_IP2_01|45|RB _DFF_IP2_01|45|MID_SHUNT _DFF_IP2_01|A4  2.1704737578552e-12
B_DFF_IP2_01|6|1 _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|6|P _DFF_IP2_01|6|MID_SERIES 0  2e-13
R_DFF_IP2_01|6|B _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SHUNT  2.7439617672
L_DFF_IP2_01|6|RB _DFF_IP2_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_01|I_1|B _DFF_IP3_01|A1 _DFF_IP3_01|I_1|MID  2e-12
I_DFF_IP3_01|I_1|B 0 _DFF_IP3_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_3|B _DFF_IP3_01|A3 _DFF_IP3_01|I_3|MID  2e-12
I_DFF_IP3_01|I_3|B 0 _DFF_IP3_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_01|I_T|B _DFF_IP3_01|T1 _DFF_IP3_01|I_T|MID  2e-12
I_DFF_IP3_01|I_T|B 0 _DFF_IP3_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_6|B _DFF_IP3_01|Q1 _DFF_IP3_01|I_6|MID  2e-12
I_DFF_IP3_01|I_6|B 0 _DFF_IP3_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_01|1|1 _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|1|P _DFF_IP3_01|1|MID_SERIES 0  2e-13
R_DFF_IP3_01|1|B _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SHUNT  2.7439617672
L_DFF_IP3_01|1|RB _DFF_IP3_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|23|1 _DFF_IP3_01|A2 _DFF_IP3_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|23|B _DFF_IP3_01|A2 _DFF_IP3_01|23|MID_SHUNT  3.84154647408
L_DFF_IP3_01|23|RB _DFF_IP3_01|23|MID_SHUNT _DFF_IP3_01|A3  2.1704737578552e-12
B_DFF_IP3_01|3|1 _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|3|P _DFF_IP3_01|3|MID_SERIES 0  2e-13
R_DFF_IP3_01|3|B _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SHUNT  2.7439617672
L_DFF_IP3_01|3|RB _DFF_IP3_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|4|1 _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|4|P _DFF_IP3_01|4|MID_SERIES 0  2e-13
R_DFF_IP3_01|4|B _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SHUNT  2.7439617672
L_DFF_IP3_01|4|RB _DFF_IP3_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|T|1 _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|T|P _DFF_IP3_01|T|MID_SERIES 0  2e-13
R_DFF_IP3_01|T|B _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SHUNT  2.7439617672
L_DFF_IP3_01|T|RB _DFF_IP3_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|45|1 _DFF_IP3_01|T2 _DFF_IP3_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|45|B _DFF_IP3_01|T2 _DFF_IP3_01|45|MID_SHUNT  3.84154647408
L_DFF_IP3_01|45|RB _DFF_IP3_01|45|MID_SHUNT _DFF_IP3_01|A4  2.1704737578552e-12
B_DFF_IP3_01|6|1 _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|6|P _DFF_IP3_01|6|MID_SERIES 0  2e-13
R_DFF_IP3_01|6|B _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SHUNT  2.7439617672
L_DFF_IP3_01|6|RB _DFF_IP3_01|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_P0_1|_TX|1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|2 JJMIT AREA=2.5
B_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|5 JJMIT AREA=2.5
I_PTL_P0_1|_TX|B1 0 _PTL_P0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_1|_TX|B2 0 _PTL_P0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|3  1.684e-12
L_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|6  3.596e-12
L_PTL_P0_1|_TX|1 P0_1 _PTL_P0_1|_TX|1  2.063e-12
L_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|4  4.123e-12
L_PTL_P0_1|_TX|3 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|7  2.193e-12
R_PTL_P0_1|_TX|D _PTL_P0_1|_TX|7 _PTL_P0_1|A_PTL  1.36
L_PTL_P0_1|_TX|P1 _PTL_P0_1|_TX|2 0  5.254e-13
L_PTL_P0_1|_TX|P2 _PTL_P0_1|_TX|5 0  5.141e-13
R_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|101  2.7439617672
R_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|104  2.7439617672
L_PTL_P0_1|_TX|RB1 _PTL_P0_1|_TX|101 0  1.550338398468e-12
L_PTL_P0_1|_TX|RB2 _PTL_P0_1|_TX|104 0  1.550338398468e-12
B_PTL_P0_1|_RX|1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|5 JJMIT AREA=2.0
B_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|8 JJMIT AREA=2.5
I_PTL_P0_1|_RX|B1 0 _PTL_P0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|3  2.777e-12
I_PTL_P0_1|_RX|B2 0 _PTL_P0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|6  2.685e-12
I_PTL_P0_1|_RX|B3 0 _PTL_P0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|9  2.764e-12
L_PTL_P0_1|_RX|1 _PTL_P0_1|A_PTL _PTL_P0_1|_RX|1  1.346e-12
L_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|4  6.348e-12
L_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7  5.197e-12
L_PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7 P0_1_RX  2.058e-12
L_PTL_P0_1|_RX|P1 _PTL_P0_1|_RX|2 0  4.795e-13
L_PTL_P0_1|_RX|P2 _PTL_P0_1|_RX|5 0  5.431e-13
L_PTL_P0_1|_RX|P3 _PTL_P0_1|_RX|8 0  5.339e-13
R_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|101  4.225701121488
R_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|104  3.429952209
R_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|107  2.7439617672
L_PTL_P0_1|_RX|RB1 _PTL_P0_1|_RX|101 0  2.38752113364072e-12
L_PTL_P0_1|_RX|RB2 _PTL_P0_1|_RX|104 0  1.937922998085e-12
L_PTL_P0_1|_RX|RB3 _PTL_P0_1|_RX|107 0  1.550338398468e-12
B_PTL_G0_1|_TX|1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|2 JJMIT AREA=2.5
B_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|5 JJMIT AREA=2.5
I_PTL_G0_1|_TX|B1 0 _PTL_G0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_1|_TX|B2 0 _PTL_G0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|3  1.684e-12
L_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|6  3.596e-12
L_PTL_G0_1|_TX|1 G0_1 _PTL_G0_1|_TX|1  2.063e-12
L_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|4  4.123e-12
L_PTL_G0_1|_TX|3 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|7  2.193e-12
R_PTL_G0_1|_TX|D _PTL_G0_1|_TX|7 _PTL_G0_1|A_PTL  1.36
L_PTL_G0_1|_TX|P1 _PTL_G0_1|_TX|2 0  5.254e-13
L_PTL_G0_1|_TX|P2 _PTL_G0_1|_TX|5 0  5.141e-13
R_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|101  2.7439617672
R_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|104  2.7439617672
L_PTL_G0_1|_TX|RB1 _PTL_G0_1|_TX|101 0  1.550338398468e-12
L_PTL_G0_1|_TX|RB2 _PTL_G0_1|_TX|104 0  1.550338398468e-12
B_PTL_G0_1|_RX|1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|5 JJMIT AREA=2.0
B_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|8 JJMIT AREA=2.5
I_PTL_G0_1|_RX|B1 0 _PTL_G0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|3  2.777e-12
I_PTL_G0_1|_RX|B2 0 _PTL_G0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|6  2.685e-12
I_PTL_G0_1|_RX|B3 0 _PTL_G0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|9  2.764e-12
L_PTL_G0_1|_RX|1 _PTL_G0_1|A_PTL _PTL_G0_1|_RX|1  1.346e-12
L_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|4  6.348e-12
L_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7  5.197e-12
L_PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7 G0_1_RX  2.058e-12
L_PTL_G0_1|_RX|P1 _PTL_G0_1|_RX|2 0  4.795e-13
L_PTL_G0_1|_RX|P2 _PTL_G0_1|_RX|5 0  5.431e-13
L_PTL_G0_1|_RX|P3 _PTL_G0_1|_RX|8 0  5.339e-13
R_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|101  4.225701121488
R_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|104  3.429952209
R_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|107  2.7439617672
L_PTL_G0_1|_RX|RB1 _PTL_G0_1|_RX|101 0  2.38752113364072e-12
L_PTL_G0_1|_RX|RB2 _PTL_G0_1|_RX|104 0  1.937922998085e-12
L_PTL_G0_1|_RX|RB3 _PTL_G0_1|_RX|107 0  1.550338398468e-12
B_PTL_G1_1|_TX|1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|2 JJMIT AREA=2.5
B_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|5 JJMIT AREA=2.5
I_PTL_G1_1|_TX|B1 0 _PTL_G1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_1|_TX|B2 0 _PTL_G1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|3  1.684e-12
L_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|6  3.596e-12
L_PTL_G1_1|_TX|1 G1_1 _PTL_G1_1|_TX|1  2.063e-12
L_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|4  4.123e-12
L_PTL_G1_1|_TX|3 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|7  2.193e-12
R_PTL_G1_1|_TX|D _PTL_G1_1|_TX|7 _PTL_G1_1|A_PTL  1.36
L_PTL_G1_1|_TX|P1 _PTL_G1_1|_TX|2 0  5.254e-13
L_PTL_G1_1|_TX|P2 _PTL_G1_1|_TX|5 0  5.141e-13
R_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|101  2.7439617672
R_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|104  2.7439617672
L_PTL_G1_1|_TX|RB1 _PTL_G1_1|_TX|101 0  1.550338398468e-12
L_PTL_G1_1|_TX|RB2 _PTL_G1_1|_TX|104 0  1.550338398468e-12
B_PTL_G1_1|_RX|1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|5 JJMIT AREA=2.0
B_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|8 JJMIT AREA=2.5
I_PTL_G1_1|_RX|B1 0 _PTL_G1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|3  2.777e-12
I_PTL_G1_1|_RX|B2 0 _PTL_G1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|6  2.685e-12
I_PTL_G1_1|_RX|B3 0 _PTL_G1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|9  2.764e-12
L_PTL_G1_1|_RX|1 _PTL_G1_1|A_PTL _PTL_G1_1|_RX|1  1.346e-12
L_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|4  6.348e-12
L_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7  5.197e-12
L_PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7 G1_1_RX  2.058e-12
L_PTL_G1_1|_RX|P1 _PTL_G1_1|_RX|2 0  4.795e-13
L_PTL_G1_1|_RX|P2 _PTL_G1_1|_RX|5 0  5.431e-13
L_PTL_G1_1|_RX|P3 _PTL_G1_1|_RX|8 0  5.339e-13
R_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|101  4.225701121488
R_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|104  3.429952209
R_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|107  2.7439617672
L_PTL_G1_1|_RX|RB1 _PTL_G1_1|_RX|101 0  2.38752113364072e-12
L_PTL_G1_1|_RX|RB2 _PTL_G1_1|_RX|104 0  1.937922998085e-12
L_PTL_G1_1|_RX|RB3 _PTL_G1_1|_RX|107 0  1.550338398468e-12
B_PTL_P2_1|_TX|1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|2 JJMIT AREA=2.5
B_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|5 JJMIT AREA=2.5
I_PTL_P2_1|_TX|B1 0 _PTL_P2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P2_1|_TX|B2 0 _PTL_P2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|3  1.684e-12
L_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|6  3.596e-12
L_PTL_P2_1|_TX|1 P2_1 _PTL_P2_1|_TX|1  2.063e-12
L_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|4  4.123e-12
L_PTL_P2_1|_TX|3 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|7  2.193e-12
R_PTL_P2_1|_TX|D _PTL_P2_1|_TX|7 _PTL_P2_1|A_PTL  1.36
L_PTL_P2_1|_TX|P1 _PTL_P2_1|_TX|2 0  5.254e-13
L_PTL_P2_1|_TX|P2 _PTL_P2_1|_TX|5 0  5.141e-13
R_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|101  2.7439617672
R_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|104  2.7439617672
L_PTL_P2_1|_TX|RB1 _PTL_P2_1|_TX|101 0  1.550338398468e-12
L_PTL_P2_1|_TX|RB2 _PTL_P2_1|_TX|104 0  1.550338398468e-12
B_PTL_P2_1|_RX|1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|5 JJMIT AREA=2.0
B_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|8 JJMIT AREA=2.5
I_PTL_P2_1|_RX|B1 0 _PTL_P2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|3  2.777e-12
I_PTL_P2_1|_RX|B2 0 _PTL_P2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|6  2.685e-12
I_PTL_P2_1|_RX|B3 0 _PTL_P2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|9  2.764e-12
L_PTL_P2_1|_RX|1 _PTL_P2_1|A_PTL _PTL_P2_1|_RX|1  1.346e-12
L_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|4  6.348e-12
L_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7  5.197e-12
L_PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7 P2_1_RX  2.058e-12
L_PTL_P2_1|_RX|P1 _PTL_P2_1|_RX|2 0  4.795e-13
L_PTL_P2_1|_RX|P2 _PTL_P2_1|_RX|5 0  5.431e-13
L_PTL_P2_1|_RX|P3 _PTL_P2_1|_RX|8 0  5.339e-13
R_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|101  4.225701121488
R_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|104  3.429952209
R_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|107  2.7439617672
L_PTL_P2_1|_RX|RB1 _PTL_P2_1|_RX|101 0  2.38752113364072e-12
L_PTL_P2_1|_RX|RB2 _PTL_P2_1|_RX|104 0  1.937922998085e-12
L_PTL_P2_1|_RX|RB3 _PTL_P2_1|_RX|107 0  1.550338398468e-12
B_PTL_G2_1|_TX|1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|2 JJMIT AREA=2.5
B_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|5 JJMIT AREA=2.5
I_PTL_G2_1|_TX|B1 0 _PTL_G2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_1|_TX|B2 0 _PTL_G2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|3  1.684e-12
L_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|6  3.596e-12
L_PTL_G2_1|_TX|1 G2_1 _PTL_G2_1|_TX|1  2.063e-12
L_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|4  4.123e-12
L_PTL_G2_1|_TX|3 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|7  2.193e-12
R_PTL_G2_1|_TX|D _PTL_G2_1|_TX|7 _PTL_G2_1|A_PTL  1.36
L_PTL_G2_1|_TX|P1 _PTL_G2_1|_TX|2 0  5.254e-13
L_PTL_G2_1|_TX|P2 _PTL_G2_1|_TX|5 0  5.141e-13
R_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|101  2.7439617672
R_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|104  2.7439617672
L_PTL_G2_1|_TX|RB1 _PTL_G2_1|_TX|101 0  1.550338398468e-12
L_PTL_G2_1|_TX|RB2 _PTL_G2_1|_TX|104 0  1.550338398468e-12
B_PTL_G2_1|_RX|1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|5 JJMIT AREA=2.0
B_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|8 JJMIT AREA=2.5
I_PTL_G2_1|_RX|B1 0 _PTL_G2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|3  2.777e-12
I_PTL_G2_1|_RX|B2 0 _PTL_G2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|6  2.685e-12
I_PTL_G2_1|_RX|B3 0 _PTL_G2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|9  2.764e-12
L_PTL_G2_1|_RX|1 _PTL_G2_1|A_PTL _PTL_G2_1|_RX|1  1.346e-12
L_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|4  6.348e-12
L_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7  5.197e-12
L_PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7 G2_1_RX  2.058e-12
L_PTL_G2_1|_RX|P1 _PTL_G2_1|_RX|2 0  4.795e-13
L_PTL_G2_1|_RX|P2 _PTL_G2_1|_RX|5 0  5.431e-13
L_PTL_G2_1|_RX|P3 _PTL_G2_1|_RX|8 0  5.339e-13
R_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|101  4.225701121488
R_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|104  3.429952209
R_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|107  2.7439617672
L_PTL_G2_1|_RX|RB1 _PTL_G2_1|_RX|101 0  2.38752113364072e-12
L_PTL_G2_1|_RX|RB2 _PTL_G2_1|_RX|104 0  1.937922998085e-12
L_PTL_G2_1|_RX|RB3 _PTL_G2_1|_RX|107 0  1.550338398468e-12
B_PTL_P3_1|_TX|1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|2 JJMIT AREA=2.5
B_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|5 JJMIT AREA=2.5
I_PTL_P3_1|_TX|B1 0 _PTL_P3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P3_1|_TX|B2 0 _PTL_P3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|3  1.684e-12
L_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|6  3.596e-12
L_PTL_P3_1|_TX|1 P3_1 _PTL_P3_1|_TX|1  2.063e-12
L_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|4  4.123e-12
L_PTL_P3_1|_TX|3 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|7  2.193e-12
R_PTL_P3_1|_TX|D _PTL_P3_1|_TX|7 _PTL_P3_1|A_PTL  1.36
L_PTL_P3_1|_TX|P1 _PTL_P3_1|_TX|2 0  5.254e-13
L_PTL_P3_1|_TX|P2 _PTL_P3_1|_TX|5 0  5.141e-13
R_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|101  2.7439617672
R_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|104  2.7439617672
L_PTL_P3_1|_TX|RB1 _PTL_P3_1|_TX|101 0  1.550338398468e-12
L_PTL_P3_1|_TX|RB2 _PTL_P3_1|_TX|104 0  1.550338398468e-12
B_PTL_P3_1|_RX|1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|5 JJMIT AREA=2.0
B_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|8 JJMIT AREA=2.5
I_PTL_P3_1|_RX|B1 0 _PTL_P3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|3  2.777e-12
I_PTL_P3_1|_RX|B2 0 _PTL_P3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|6  2.685e-12
I_PTL_P3_1|_RX|B3 0 _PTL_P3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|9  2.764e-12
L_PTL_P3_1|_RX|1 _PTL_P3_1|A_PTL _PTL_P3_1|_RX|1  1.346e-12
L_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|4  6.348e-12
L_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7  5.197e-12
L_PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7 P3_1_RX  2.058e-12
L_PTL_P3_1|_RX|P1 _PTL_P3_1|_RX|2 0  4.795e-13
L_PTL_P3_1|_RX|P2 _PTL_P3_1|_RX|5 0  5.431e-13
L_PTL_P3_1|_RX|P3 _PTL_P3_1|_RX|8 0  5.339e-13
R_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|101  4.225701121488
R_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|104  3.429952209
R_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|107  2.7439617672
L_PTL_P3_1|_RX|RB1 _PTL_P3_1|_RX|101 0  2.38752113364072e-12
L_PTL_P3_1|_RX|RB2 _PTL_P3_1|_RX|104 0  1.937922998085e-12
L_PTL_P3_1|_RX|RB3 _PTL_P3_1|_RX|107 0  1.550338398468e-12
B_PTL_G3_1|_TX|1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|2 JJMIT AREA=2.5
B_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|5 JJMIT AREA=2.5
I_PTL_G3_1|_TX|B1 0 _PTL_G3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_1|_TX|B2 0 _PTL_G3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|3  1.684e-12
L_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|6  3.596e-12
L_PTL_G3_1|_TX|1 G3_1 _PTL_G3_1|_TX|1  2.063e-12
L_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|4  4.123e-12
L_PTL_G3_1|_TX|3 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|7  2.193e-12
R_PTL_G3_1|_TX|D _PTL_G3_1|_TX|7 _PTL_G3_1|A_PTL  1.36
L_PTL_G3_1|_TX|P1 _PTL_G3_1|_TX|2 0  5.254e-13
L_PTL_G3_1|_TX|P2 _PTL_G3_1|_TX|5 0  5.141e-13
R_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|101  2.7439617672
R_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|104  2.7439617672
L_PTL_G3_1|_TX|RB1 _PTL_G3_1|_TX|101 0  1.550338398468e-12
L_PTL_G3_1|_TX|RB2 _PTL_G3_1|_TX|104 0  1.550338398468e-12
B_PTL_G3_1|_RX|1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|5 JJMIT AREA=2.0
B_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|8 JJMIT AREA=2.5
I_PTL_G3_1|_RX|B1 0 _PTL_G3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|3  2.777e-12
I_PTL_G3_1|_RX|B2 0 _PTL_G3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|6  2.685e-12
I_PTL_G3_1|_RX|B3 0 _PTL_G3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|9  2.764e-12
L_PTL_G3_1|_RX|1 _PTL_G3_1|A_PTL _PTL_G3_1|_RX|1  1.346e-12
L_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|4  6.348e-12
L_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7  5.197e-12
L_PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7 G3_1_RX  2.058e-12
L_PTL_G3_1|_RX|P1 _PTL_G3_1|_RX|2 0  4.795e-13
L_PTL_G3_1|_RX|P2 _PTL_G3_1|_RX|5 0  5.431e-13
L_PTL_G3_1|_RX|P3 _PTL_G3_1|_RX|8 0  5.339e-13
R_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|101  4.225701121488
R_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|104  3.429952209
R_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|107  2.7439617672
L_PTL_G3_1|_RX|RB1 _PTL_G3_1|_RX|101 0  2.38752113364072e-12
L_PTL_G3_1|_RX|RB2 _PTL_G3_1|_RX|104 0  1.937922998085e-12
L_PTL_G3_1|_RX|RB3 _PTL_G3_1|_RX|107 0  1.550338398468e-12
B_PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_1|_TX|B1 0 _PTL_IP1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_1|_TX|B2 0 _PTL_IP1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|3  1.684e-12
L_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|6  3.596e-12
L_PTL_IP1_1|_TX|1 IP1_1_OUT _PTL_IP1_1|_TX|1  2.063e-12
L_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|4  4.123e-12
L_PTL_IP1_1|_TX|3 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|7  2.193e-12
R_PTL_IP1_1|_TX|D _PTL_IP1_1|_TX|7 _PTL_IP1_1|A_PTL  1.36
L_PTL_IP1_1|_TX|P1 _PTL_IP1_1|_TX|2 0  5.254e-13
L_PTL_IP1_1|_TX|P2 _PTL_IP1_1|_TX|5 0  5.141e-13
R_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|101  2.7439617672
R_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|104  2.7439617672
L_PTL_IP1_1|_TX|RB1 _PTL_IP1_1|_TX|101 0  1.550338398468e-12
L_PTL_IP1_1|_TX|RB2 _PTL_IP1_1|_TX|104 0  1.550338398468e-12
B_PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_1|_RX|B1 0 _PTL_IP1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|3  2.777e-12
I_PTL_IP1_1|_RX|B2 0 _PTL_IP1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|6  2.685e-12
I_PTL_IP1_1|_RX|B3 0 _PTL_IP1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|9  2.764e-12
L_PTL_IP1_1|_RX|1 _PTL_IP1_1|A_PTL _PTL_IP1_1|_RX|1  1.346e-12
L_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|4  6.348e-12
L_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7  5.197e-12
L_PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7 IP1_1_OUT_RX  2.058e-12
L_PTL_IP1_1|_RX|P1 _PTL_IP1_1|_RX|2 0  4.795e-13
L_PTL_IP1_1|_RX|P2 _PTL_IP1_1|_RX|5 0  5.431e-13
L_PTL_IP1_1|_RX|P3 _PTL_IP1_1|_RX|8 0  5.339e-13
R_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|101  4.225701121488
R_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|104  3.429952209
R_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|107  2.7439617672
L_PTL_IP1_1|_RX|RB1 _PTL_IP1_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_1|_RX|RB2 _PTL_IP1_1|_RX|104 0  1.937922998085e-12
L_PTL_IP1_1|_RX|RB3 _PTL_IP1_1|_RX|107 0  1.550338398468e-12
B_PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_1|_TX|B1 0 _PTL_IP2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_1|_TX|B2 0 _PTL_IP2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|3  1.684e-12
L_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|6  3.596e-12
L_PTL_IP2_1|_TX|1 IP2_1_OUT _PTL_IP2_1|_TX|1  2.063e-12
L_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|4  4.123e-12
L_PTL_IP2_1|_TX|3 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|7  2.193e-12
R_PTL_IP2_1|_TX|D _PTL_IP2_1|_TX|7 _PTL_IP2_1|A_PTL  1.36
L_PTL_IP2_1|_TX|P1 _PTL_IP2_1|_TX|2 0  5.254e-13
L_PTL_IP2_1|_TX|P2 _PTL_IP2_1|_TX|5 0  5.141e-13
R_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|101  2.7439617672
R_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|104  2.7439617672
L_PTL_IP2_1|_TX|RB1 _PTL_IP2_1|_TX|101 0  1.550338398468e-12
L_PTL_IP2_1|_TX|RB2 _PTL_IP2_1|_TX|104 0  1.550338398468e-12
B_PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_1|_RX|B1 0 _PTL_IP2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|3  2.777e-12
I_PTL_IP2_1|_RX|B2 0 _PTL_IP2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|6  2.685e-12
I_PTL_IP2_1|_RX|B3 0 _PTL_IP2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|9  2.764e-12
L_PTL_IP2_1|_RX|1 _PTL_IP2_1|A_PTL _PTL_IP2_1|_RX|1  1.346e-12
L_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|4  6.348e-12
L_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7  5.197e-12
L_PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7 IP2_1_OUT_RX  2.058e-12
L_PTL_IP2_1|_RX|P1 _PTL_IP2_1|_RX|2 0  4.795e-13
L_PTL_IP2_1|_RX|P2 _PTL_IP2_1|_RX|5 0  5.431e-13
L_PTL_IP2_1|_RX|P3 _PTL_IP2_1|_RX|8 0  5.339e-13
R_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|101  4.225701121488
R_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|104  3.429952209
R_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|107  2.7439617672
L_PTL_IP2_1|_RX|RB1 _PTL_IP2_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_1|_RX|RB2 _PTL_IP2_1|_RX|104 0  1.937922998085e-12
L_PTL_IP2_1|_RX|RB3 _PTL_IP2_1|_RX|107 0  1.550338398468e-12
B_PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_1|_TX|B1 0 _PTL_IP3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_1|_TX|B2 0 _PTL_IP3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|3  1.684e-12
L_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|6  3.596e-12
L_PTL_IP3_1|_TX|1 IP3_1_OUT _PTL_IP3_1|_TX|1  2.063e-12
L_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|4  4.123e-12
L_PTL_IP3_1|_TX|3 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|7  2.193e-12
R_PTL_IP3_1|_TX|D _PTL_IP3_1|_TX|7 _PTL_IP3_1|A_PTL  1.36
L_PTL_IP3_1|_TX|P1 _PTL_IP3_1|_TX|2 0  5.254e-13
L_PTL_IP3_1|_TX|P2 _PTL_IP3_1|_TX|5 0  5.141e-13
R_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|101  2.7439617672
R_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|104  2.7439617672
L_PTL_IP3_1|_TX|RB1 _PTL_IP3_1|_TX|101 0  1.550338398468e-12
L_PTL_IP3_1|_TX|RB2 _PTL_IP3_1|_TX|104 0  1.550338398468e-12
B_PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_1|_RX|B1 0 _PTL_IP3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|3  2.777e-12
I_PTL_IP3_1|_RX|B2 0 _PTL_IP3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|6  2.685e-12
I_PTL_IP3_1|_RX|B3 0 _PTL_IP3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|9  2.764e-12
L_PTL_IP3_1|_RX|1 _PTL_IP3_1|A_PTL _PTL_IP3_1|_RX|1  1.346e-12
L_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|4  6.348e-12
L_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7  5.197e-12
L_PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7 IP3_1_OUT_RX  2.058e-12
L_PTL_IP3_1|_RX|P1 _PTL_IP3_1|_RX|2 0  4.795e-13
L_PTL_IP3_1|_RX|P2 _PTL_IP3_1|_RX|5 0  5.431e-13
L_PTL_IP3_1|_RX|P3 _PTL_IP3_1|_RX|8 0  5.339e-13
R_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|101  4.225701121488
R_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|104  3.429952209
R_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|107  2.7439617672
L_PTL_IP3_1|_RX|RB1 _PTL_IP3_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_1|_RX|RB2 _PTL_IP3_1|_RX|104 0  1.937922998085e-12
L_PTL_IP3_1|_RX|RB3 _PTL_IP3_1|_RX|107 0  1.550338398468e-12
LSPL_G1_1|SPL1|1 G1_1_RX SPL_G1_1|SPL1|D1  2e-12
LSPL_G1_1|SPL1|2 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|D2  4.135667696e-12
LSPL_G1_1|SPL1|3 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|JCT  9.84682784761905e-13
LSPL_G1_1|SPL1|4 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QA1  9.84682784761905e-13
LSPL_G1_1|SPL1|5 SPL_G1_1|SPL1|QA1 G1_1_TO1  2e-12
LSPL_G1_1|SPL1|6 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QB1  9.84682784761905e-13
LSPL_G1_1|SPL1|7 SPL_G1_1|SPL1|QB1 SPL_G1_1|QTMP  2e-12
LSPL_G1_1|SPL2|1 SPL_G1_1|QTMP SPL_G1_1|SPL2|D1  2e-12
LSPL_G1_1|SPL2|2 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|D2  4.135667696e-12
LSPL_G1_1|SPL2|3 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|JCT  9.84682784761905e-13
LSPL_G1_1|SPL2|4 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QA1  9.84682784761905e-13
LSPL_G1_1|SPL2|5 SPL_G1_1|SPL2|QA1 G1_1_TO2  2e-12
LSPL_G1_1|SPL2|6 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QB1  9.84682784761905e-13
LSPL_G1_1|SPL2|7 SPL_G1_1|SPL2|QB1 G1_1_TO3  2e-12
L_PG0_12|P|1 P0_1_RX _PG0_12|P|A1  2.067833848e-12
L_PG0_12|P|2 _PG0_12|P|A1 _PG0_12|P|A2  4.135667696e-12
L_PG0_12|P|3 _PG0_12|P|A3 _PG0_12|P|A4  8.271335392e-12
L_PG0_12|P|T T08 _PG0_12|P|T1  2.067833848e-12
L_PG0_12|P|4 _PG0_12|P|T1 _PG0_12|P|T2  4.135667696e-12
L_PG0_12|P|5 _PG0_12|P|A4 _PG0_12|P|Q1  4.135667696e-12
L_PG0_12|P|6 _PG0_12|P|Q1 P0_2  2.067833848e-12
L_PG0_12|G|1 G0_1_RX _PG0_12|G|A1  2.067833848e-12
L_PG0_12|G|2 _PG0_12|G|A1 _PG0_12|G|A2  4.135667696e-12
L_PG0_12|G|3 _PG0_12|G|A3 _PG0_12|G|A4  8.271335392e-12
L_PG0_12|G|T T08 _PG0_12|G|T1  2.067833848e-12
L_PG0_12|G|4 _PG0_12|G|T1 _PG0_12|G|T2  4.135667696e-12
L_PG0_12|G|5 _PG0_12|G|A4 _PG0_12|G|Q1  4.135667696e-12
L_PG0_12|G|6 _PG0_12|G|Q1 G0_2  2.067833848e-12
L_PG1_12|I_1|B _PG1_12|A1 _PG1_12|I_1|MID  2e-12
I_PG1_12|I_1|B 0 _PG1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_3|B _PG1_12|A3 _PG1_12|I_3|MID  2e-12
I_PG1_12|I_3|B 0 _PG1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_12|I_T|B _PG1_12|T1 _PG1_12|I_T|MID  2e-12
I_PG1_12|I_T|B 0 _PG1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_6|B _PG1_12|Q1 _PG1_12|I_6|MID  2e-12
I_PG1_12|I_6|B 0 _PG1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_12|1|1 _PG1_12|A1 _PG1_12|1|MID_SERIES JJMIT AREA=2.5
L_PG1_12|1|P _PG1_12|1|MID_SERIES 0  2e-13
R_PG1_12|1|B _PG1_12|A1 _PG1_12|1|MID_SHUNT  2.7439617672
L_PG1_12|1|RB _PG1_12|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|23|1 _PG1_12|A2 _PG1_12|A3 JJMIT AREA=1.7857142857142858
R_PG1_12|23|B _PG1_12|A2 _PG1_12|23|MID_SHUNT  3.84154647408
L_PG1_12|23|RB _PG1_12|23|MID_SHUNT _PG1_12|A3  2.1704737578552e-12
B_PG1_12|3|1 _PG1_12|A3 _PG1_12|3|MID_SERIES JJMIT AREA=2.5
L_PG1_12|3|P _PG1_12|3|MID_SERIES 0  2e-13
R_PG1_12|3|B _PG1_12|A3 _PG1_12|3|MID_SHUNT  2.7439617672
L_PG1_12|3|RB _PG1_12|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|4|1 _PG1_12|A4 _PG1_12|4|MID_SERIES JJMIT AREA=2.5
L_PG1_12|4|P _PG1_12|4|MID_SERIES 0  2e-13
R_PG1_12|4|B _PG1_12|A4 _PG1_12|4|MID_SHUNT  2.7439617672
L_PG1_12|4|RB _PG1_12|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|T|1 _PG1_12|T1 _PG1_12|T|MID_SERIES JJMIT AREA=2.5
L_PG1_12|T|P _PG1_12|T|MID_SERIES 0  2e-13
R_PG1_12|T|B _PG1_12|T1 _PG1_12|T|MID_SHUNT  2.7439617672
L_PG1_12|T|RB _PG1_12|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|45|1 _PG1_12|T2 _PG1_12|A4 JJMIT AREA=1.7857142857142858
R_PG1_12|45|B _PG1_12|T2 _PG1_12|45|MID_SHUNT  3.84154647408
L_PG1_12|45|RB _PG1_12|45|MID_SHUNT _PG1_12|A4  2.1704737578552e-12
B_PG1_12|6|1 _PG1_12|Q1 _PG1_12|6|MID_SERIES JJMIT AREA=2.5
L_PG1_12|6|P _PG1_12|6|MID_SERIES 0  2e-13
R_PG1_12|6|B _PG1_12|Q1 _PG1_12|6|MID_SHUNT  2.7439617672
L_PG1_12|6|RB _PG1_12|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|1 G2_1_RX _PG2_12|_SPL_G1|D1  2e-12
L_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|D2  4.135667696e-12
L_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG2_12|_SPL_G1|5 _PG2_12|_SPL_G1|QA1 _PG2_12|G1_COPY_1  2e-12
L_PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|QB1 _PG2_12|G1_COPY_2  2e-12
L_PG2_12|_PG|A1 P2_1_RX _PG2_12|_PG|A1  2.067833848e-12
L_PG2_12|_PG|A2 _PG2_12|_PG|A1 _PG2_12|_PG|A2  4.135667696e-12
L_PG2_12|_PG|A3 _PG2_12|_PG|A3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|B1 _PG2_12|G1_COPY_1 _PG2_12|_PG|B1  2.067833848e-12
L_PG2_12|_PG|B2 _PG2_12|_PG|B1 _PG2_12|_PG|B2  4.135667696e-12
L_PG2_12|_PG|B3 _PG2_12|_PG|B3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|Q3 _PG2_12|_PG|Q3 _PG2_12|_PG|Q2  4.135667696e-12
L_PG2_12|_PG|Q2 _PG2_12|_PG|Q2 _PG2_12|_PG|Q1  4.135667696e-12
L_PG2_12|_PG|Q1 _PG2_12|_PG|Q1 _PG2_12|PG  2.067833848e-12
L_PG2_12|_GG|A1 G1_1_TO2 _PG2_12|_GG|A1  2.067833848e-12
L_PG2_12|_GG|A2 _PG2_12|_GG|A1 _PG2_12|_GG|A2  4.135667696e-12
L_PG2_12|_GG|A3 _PG2_12|_GG|A3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|B1 _PG2_12|G1_COPY_2 _PG2_12|_GG|B1  2.067833848e-12
L_PG2_12|_GG|B2 _PG2_12|_GG|B1 _PG2_12|_GG|B2  4.135667696e-12
L_PG2_12|_GG|B3 _PG2_12|_GG|B3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|Q3 _PG2_12|_GG|Q3 _PG2_12|_GG|Q2  4.135667696e-12
L_PG2_12|_GG|Q2 _PG2_12|_GG|Q2 _PG2_12|_GG|Q1  4.135667696e-12
L_PG2_12|_GG|Q1 _PG2_12|_GG|Q1 _PG2_12|GG  2.067833848e-12
L_PG2_12|_DFF_PG|1 _PG2_12|PG _PG2_12|_DFF_PG|A1  2.067833848e-12
L_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|A2  4.135667696e-12
L_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|A4  8.271335392e-12
L_PG2_12|_DFF_PG|T T10 _PG2_12|_DFF_PG|T1  2.067833848e-12
L_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T2  4.135667696e-12
L_PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|Q1  4.135667696e-12
L_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|Q1 _PG2_12|PG_SYNC  2.067833848e-12
L_PG2_12|_DFF_GG|1 _PG2_12|GG _PG2_12|_DFF_GG|A1  2.067833848e-12
L_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|A2  4.135667696e-12
L_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|A4  8.271335392e-12
L_PG2_12|_DFF_GG|T T10 _PG2_12|_DFF_GG|T1  2.067833848e-12
L_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T2  4.135667696e-12
L_PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|Q1  4.135667696e-12
L_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|Q1 _PG2_12|GG_SYNC  2.067833848e-12
L_PG2_12|_AND_G|A1 _PG2_12|PG_SYNC _PG2_12|_AND_G|A1  2.067833848e-12
L_PG2_12|_AND_G|A2 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A2  4.135667696e-12
L_PG2_12|_AND_G|A3 _PG2_12|_AND_G|A3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|B1 _PG2_12|GG_SYNC _PG2_12|_AND_G|B1  2.067833848e-12
L_PG2_12|_AND_G|B2 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B2  4.135667696e-12
L_PG2_12|_AND_G|B3 _PG2_12|_AND_G|B3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q2  4.135667696e-12
L_PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q1  4.135667696e-12
L_PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1 G2_2  2.067833848e-12
L_PG3_12|_SPL_G1|1 G3_1_RX _PG3_12|_SPL_G1|D1  2e-12
L_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|D2  4.135667696e-12
L_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_12|_SPL_G1|5 _PG3_12|_SPL_G1|QA1 _PG3_12|G1_COPY_1  2e-12
L_PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|QB1 _PG3_12|G1_COPY_2  2e-12
L_PG3_12|_PG|A1 P3_1_RX _PG3_12|_PG|A1  2.067833848e-12
L_PG3_12|_PG|A2 _PG3_12|_PG|A1 _PG3_12|_PG|A2  4.135667696e-12
L_PG3_12|_PG|A3 _PG3_12|_PG|A3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|B1 _PG3_12|G1_COPY_1 _PG3_12|_PG|B1  2.067833848e-12
L_PG3_12|_PG|B2 _PG3_12|_PG|B1 _PG3_12|_PG|B2  4.135667696e-12
L_PG3_12|_PG|B3 _PG3_12|_PG|B3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|Q3 _PG3_12|_PG|Q3 _PG3_12|_PG|Q2  4.135667696e-12
L_PG3_12|_PG|Q2 _PG3_12|_PG|Q2 _PG3_12|_PG|Q1  4.135667696e-12
L_PG3_12|_PG|Q1 _PG3_12|_PG|Q1 _PG3_12|PG  2.067833848e-12
L_PG3_12|_GG|A1 G1_1_TO3 _PG3_12|_GG|A1  2.067833848e-12
L_PG3_12|_GG|A2 _PG3_12|_GG|A1 _PG3_12|_GG|A2  4.135667696e-12
L_PG3_12|_GG|A3 _PG3_12|_GG|A3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|B1 _PG3_12|G1_COPY_2 _PG3_12|_GG|B1  2.067833848e-12
L_PG3_12|_GG|B2 _PG3_12|_GG|B1 _PG3_12|_GG|B2  4.135667696e-12
L_PG3_12|_GG|B3 _PG3_12|_GG|B3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|Q3 _PG3_12|_GG|Q3 _PG3_12|_GG|Q2  4.135667696e-12
L_PG3_12|_GG|Q2 _PG3_12|_GG|Q2 _PG3_12|_GG|Q1  4.135667696e-12
L_PG3_12|_GG|Q1 _PG3_12|_GG|Q1 _PG3_12|GG  2.067833848e-12
L_PG3_12|_DFF_PG|1 _PG3_12|PG _PG3_12|_DFF_PG|A1  2.067833848e-12
L_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|A2  4.135667696e-12
L_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|A4  8.271335392e-12
L_PG3_12|_DFF_PG|T T11 _PG3_12|_DFF_PG|T1  2.067833848e-12
L_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T2  4.135667696e-12
L_PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|Q1  4.135667696e-12
L_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|Q1 _PG3_12|PG_SYNC  2.067833848e-12
L_PG3_12|_DFF_GG|1 _PG3_12|GG _PG3_12|_DFF_GG|A1  2.067833848e-12
L_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|A2  4.135667696e-12
L_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|A4  8.271335392e-12
L_PG3_12|_DFF_GG|T T11 _PG3_12|_DFF_GG|T1  2.067833848e-12
L_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T2  4.135667696e-12
L_PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|Q1  4.135667696e-12
L_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|Q1 _PG3_12|GG_SYNC  2.067833848e-12
L_PG3_12|_AND_G|A1 _PG3_12|PG_SYNC _PG3_12|_AND_G|A1  2.067833848e-12
L_PG3_12|_AND_G|A2 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A2  4.135667696e-12
L_PG3_12|_AND_G|A3 _PG3_12|_AND_G|A3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|B1 _PG3_12|GG_SYNC _PG3_12|_AND_G|B1  2.067833848e-12
L_PG3_12|_AND_G|B2 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B2  4.135667696e-12
L_PG3_12|_AND_G|B3 _PG3_12|_AND_G|B3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q2  4.135667696e-12
L_PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q1  4.135667696e-12
L_PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1 G3_2  2.067833848e-12
L_DFF_IP1_12|I_1|B _DFF_IP1_12|A1 _DFF_IP1_12|I_1|MID  2e-12
I_DFF_IP1_12|I_1|B 0 _DFF_IP1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_3|B _DFF_IP1_12|A3 _DFF_IP1_12|I_3|MID  2e-12
I_DFF_IP1_12|I_3|B 0 _DFF_IP1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_12|I_T|B _DFF_IP1_12|T1 _DFF_IP1_12|I_T|MID  2e-12
I_DFF_IP1_12|I_T|B 0 _DFF_IP1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_6|B _DFF_IP1_12|Q1 _DFF_IP1_12|I_6|MID  2e-12
I_DFF_IP1_12|I_6|B 0 _DFF_IP1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_12|1|1 _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|1|P _DFF_IP1_12|1|MID_SERIES 0  2e-13
R_DFF_IP1_12|1|B _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SHUNT  2.7439617672
L_DFF_IP1_12|1|RB _DFF_IP1_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|23|1 _DFF_IP1_12|A2 _DFF_IP1_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|23|B _DFF_IP1_12|A2 _DFF_IP1_12|23|MID_SHUNT  3.84154647408
L_DFF_IP1_12|23|RB _DFF_IP1_12|23|MID_SHUNT _DFF_IP1_12|A3  2.1704737578552e-12
B_DFF_IP1_12|3|1 _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|3|P _DFF_IP1_12|3|MID_SERIES 0  2e-13
R_DFF_IP1_12|3|B _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SHUNT  2.7439617672
L_DFF_IP1_12|3|RB _DFF_IP1_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|4|1 _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|4|P _DFF_IP1_12|4|MID_SERIES 0  2e-13
R_DFF_IP1_12|4|B _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SHUNT  2.7439617672
L_DFF_IP1_12|4|RB _DFF_IP1_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|T|1 _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|T|P _DFF_IP1_12|T|MID_SERIES 0  2e-13
R_DFF_IP1_12|T|B _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SHUNT  2.7439617672
L_DFF_IP1_12|T|RB _DFF_IP1_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|45|1 _DFF_IP1_12|T2 _DFF_IP1_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|45|B _DFF_IP1_12|T2 _DFF_IP1_12|45|MID_SHUNT  3.84154647408
L_DFF_IP1_12|45|RB _DFF_IP1_12|45|MID_SHUNT _DFF_IP1_12|A4  2.1704737578552e-12
B_DFF_IP1_12|6|1 _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|6|P _DFF_IP1_12|6|MID_SERIES 0  2e-13
R_DFF_IP1_12|6|B _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SHUNT  2.7439617672
L_DFF_IP1_12|6|RB _DFF_IP1_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_12|I_1|B _DFF_IP2_12|A1 _DFF_IP2_12|I_1|MID  2e-12
I_DFF_IP2_12|I_1|B 0 _DFF_IP2_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_3|B _DFF_IP2_12|A3 _DFF_IP2_12|I_3|MID  2e-12
I_DFF_IP2_12|I_3|B 0 _DFF_IP2_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_12|I_T|B _DFF_IP2_12|T1 _DFF_IP2_12|I_T|MID  2e-12
I_DFF_IP2_12|I_T|B 0 _DFF_IP2_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_6|B _DFF_IP2_12|Q1 _DFF_IP2_12|I_6|MID  2e-12
I_DFF_IP2_12|I_6|B 0 _DFF_IP2_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_12|1|1 _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|1|P _DFF_IP2_12|1|MID_SERIES 0  2e-13
R_DFF_IP2_12|1|B _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SHUNT  2.7439617672
L_DFF_IP2_12|1|RB _DFF_IP2_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|23|1 _DFF_IP2_12|A2 _DFF_IP2_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|23|B _DFF_IP2_12|A2 _DFF_IP2_12|23|MID_SHUNT  3.84154647408
L_DFF_IP2_12|23|RB _DFF_IP2_12|23|MID_SHUNT _DFF_IP2_12|A3  2.1704737578552e-12
B_DFF_IP2_12|3|1 _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|3|P _DFF_IP2_12|3|MID_SERIES 0  2e-13
R_DFF_IP2_12|3|B _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SHUNT  2.7439617672
L_DFF_IP2_12|3|RB _DFF_IP2_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|4|1 _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|4|P _DFF_IP2_12|4|MID_SERIES 0  2e-13
R_DFF_IP2_12|4|B _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SHUNT  2.7439617672
L_DFF_IP2_12|4|RB _DFF_IP2_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|T|1 _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|T|P _DFF_IP2_12|T|MID_SERIES 0  2e-13
R_DFF_IP2_12|T|B _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SHUNT  2.7439617672
L_DFF_IP2_12|T|RB _DFF_IP2_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|45|1 _DFF_IP2_12|T2 _DFF_IP2_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|45|B _DFF_IP2_12|T2 _DFF_IP2_12|45|MID_SHUNT  3.84154647408
L_DFF_IP2_12|45|RB _DFF_IP2_12|45|MID_SHUNT _DFF_IP2_12|A4  2.1704737578552e-12
B_DFF_IP2_12|6|1 _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|6|P _DFF_IP2_12|6|MID_SERIES 0  2e-13
R_DFF_IP2_12|6|B _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SHUNT  2.7439617672
L_DFF_IP2_12|6|RB _DFF_IP2_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_12|I_1|B _DFF_IP3_12|A1 _DFF_IP3_12|I_1|MID  2e-12
I_DFF_IP3_12|I_1|B 0 _DFF_IP3_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_3|B _DFF_IP3_12|A3 _DFF_IP3_12|I_3|MID  2e-12
I_DFF_IP3_12|I_3|B 0 _DFF_IP3_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_12|I_T|B _DFF_IP3_12|T1 _DFF_IP3_12|I_T|MID  2e-12
I_DFF_IP3_12|I_T|B 0 _DFF_IP3_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_6|B _DFF_IP3_12|Q1 _DFF_IP3_12|I_6|MID  2e-12
I_DFF_IP3_12|I_6|B 0 _DFF_IP3_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_12|1|1 _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|1|P _DFF_IP3_12|1|MID_SERIES 0  2e-13
R_DFF_IP3_12|1|B _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SHUNT  2.7439617672
L_DFF_IP3_12|1|RB _DFF_IP3_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|23|1 _DFF_IP3_12|A2 _DFF_IP3_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|23|B _DFF_IP3_12|A2 _DFF_IP3_12|23|MID_SHUNT  3.84154647408
L_DFF_IP3_12|23|RB _DFF_IP3_12|23|MID_SHUNT _DFF_IP3_12|A3  2.1704737578552e-12
B_DFF_IP3_12|3|1 _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|3|P _DFF_IP3_12|3|MID_SERIES 0  2e-13
R_DFF_IP3_12|3|B _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SHUNT  2.7439617672
L_DFF_IP3_12|3|RB _DFF_IP3_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|4|1 _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|4|P _DFF_IP3_12|4|MID_SERIES 0  2e-13
R_DFF_IP3_12|4|B _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SHUNT  2.7439617672
L_DFF_IP3_12|4|RB _DFF_IP3_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|T|1 _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|T|P _DFF_IP3_12|T|MID_SERIES 0  2e-13
R_DFF_IP3_12|T|B _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SHUNT  2.7439617672
L_DFF_IP3_12|T|RB _DFF_IP3_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|45|1 _DFF_IP3_12|T2 _DFF_IP3_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|45|B _DFF_IP3_12|T2 _DFF_IP3_12|45|MID_SHUNT  3.84154647408
L_DFF_IP3_12|45|RB _DFF_IP3_12|45|MID_SHUNT _DFF_IP3_12|A4  2.1704737578552e-12
B_DFF_IP3_12|6|1 _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|6|P _DFF_IP3_12|6|MID_SERIES 0  2e-13
R_DFF_IP3_12|6|B _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SHUNT  2.7439617672
L_DFF_IP3_12|6|RB _DFF_IP3_12|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_P0_2|_TX|1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|2 JJMIT AREA=2.5
B_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|5 JJMIT AREA=2.5
I_PTL_P0_2|_TX|B1 0 _PTL_P0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_2|_TX|B2 0 _PTL_P0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|3  1.684e-12
L_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|6  3.596e-12
L_PTL_P0_2|_TX|1 P0_2 _PTL_P0_2|_TX|1  2.063e-12
L_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|4  4.123e-12
L_PTL_P0_2|_TX|3 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|7  2.193e-12
R_PTL_P0_2|_TX|D _PTL_P0_2|_TX|7 _PTL_P0_2|A_PTL  1.36
L_PTL_P0_2|_TX|P1 _PTL_P0_2|_TX|2 0  5.254e-13
L_PTL_P0_2|_TX|P2 _PTL_P0_2|_TX|5 0  5.141e-13
R_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|101  2.7439617672
R_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|104  2.7439617672
L_PTL_P0_2|_TX|RB1 _PTL_P0_2|_TX|101 0  1.550338398468e-12
L_PTL_P0_2|_TX|RB2 _PTL_P0_2|_TX|104 0  1.550338398468e-12
B_PTL_P0_2|_RX|1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|5 JJMIT AREA=2.0
B_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|8 JJMIT AREA=2.5
I_PTL_P0_2|_RX|B1 0 _PTL_P0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|3  2.777e-12
I_PTL_P0_2|_RX|B2 0 _PTL_P0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|6  2.685e-12
I_PTL_P0_2|_RX|B3 0 _PTL_P0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|9  2.764e-12
L_PTL_P0_2|_RX|1 _PTL_P0_2|A_PTL _PTL_P0_2|_RX|1  1.346e-12
L_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|4  6.348e-12
L_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7  5.197e-12
L_PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7 _PTL_P0_2|A_PTL_RX  2.058e-12
L_PTL_P0_2|_RX|P1 _PTL_P0_2|_RX|2 0  4.795e-13
L_PTL_P0_2|_RX|P2 _PTL_P0_2|_RX|5 0  5.431e-13
L_PTL_P0_2|_RX|P3 _PTL_P0_2|_RX|8 0  5.339e-13
R_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|101  4.225701121488
R_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|104  3.429952209
R_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|107  2.7439617672
L_PTL_P0_2|_RX|RB1 _PTL_P0_2|_RX|101 0  2.38752113364072e-12
L_PTL_P0_2|_RX|RB2 _PTL_P0_2|_RX|104 0  1.937922998085e-12
L_PTL_P0_2|_RX|RB3 _PTL_P0_2|_RX|107 0  1.550338398468e-12
B_PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|2 JJMIT AREA=2.5
B_PTL_P0_2|_JTL|2 _PTL_P0_2|_JTL|6 _PTL_P0_2|_JTL|7 JJMIT AREA=2.5
I_PTL_P0_2|_JTL|B1 0 _PTL_P0_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_P0_2|_JTL|1 _PTL_P0_2|A_PTL_RX _PTL_P0_2|_JTL|1  2.067833848e-12
L_PTL_P0_2|_JTL|2 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|4  2.067833848e-12
L_PTL_P0_2|_JTL|3 _PTL_P0_2|_JTL|4 _PTL_P0_2|_JTL|6  2.067833848e-12
L_PTL_P0_2|_JTL|4 _PTL_P0_2|_JTL|6 P0_2_RX  2.067833848e-12
L_PTL_P0_2|_JTL|P1 _PTL_P0_2|_JTL|2 0  2e-13
L_PTL_P0_2|_JTL|P2 _PTL_P0_2|_JTL|7 0  2e-13
L_PTL_P0_2|_JTL|B1 _PTL_P0_2|_JTL|5 _PTL_P0_2|_JTL|4  2e-12
R_PTL_P0_2|_JTL|B1 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|3  2.7439617672
R_PTL_P0_2|_JTL|B2 _PTL_P0_2|_JTL|6 _PTL_P0_2|_JTL|8  2.7439617672
L_PTL_P0_2|_JTL|RB1 _PTL_P0_2|_JTL|3 0  1.750338398468e-12
L_PTL_P0_2|_JTL|RB2 _PTL_P0_2|_JTL|8 0  1.750338398468e-12
B_PTL_G0_2|_TX|1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|2 JJMIT AREA=2.5
B_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|5 JJMIT AREA=2.5
I_PTL_G0_2|_TX|B1 0 _PTL_G0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_2|_TX|B2 0 _PTL_G0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|3  1.684e-12
L_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|6  3.596e-12
L_PTL_G0_2|_TX|1 G0_2 _PTL_G0_2|_TX|1  2.063e-12
L_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|4  4.123e-12
L_PTL_G0_2|_TX|3 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|7  2.193e-12
R_PTL_G0_2|_TX|D _PTL_G0_2|_TX|7 _PTL_G0_2|A_PTL  1.36
L_PTL_G0_2|_TX|P1 _PTL_G0_2|_TX|2 0  5.254e-13
L_PTL_G0_2|_TX|P2 _PTL_G0_2|_TX|5 0  5.141e-13
R_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|101  2.7439617672
R_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|104  2.7439617672
L_PTL_G0_2|_TX|RB1 _PTL_G0_2|_TX|101 0  1.550338398468e-12
L_PTL_G0_2|_TX|RB2 _PTL_G0_2|_TX|104 0  1.550338398468e-12
B_PTL_G0_2|_RX|1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|5 JJMIT AREA=2.0
B_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|8 JJMIT AREA=2.5
I_PTL_G0_2|_RX|B1 0 _PTL_G0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|3  2.777e-12
I_PTL_G0_2|_RX|B2 0 _PTL_G0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|6  2.685e-12
I_PTL_G0_2|_RX|B3 0 _PTL_G0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|9  2.764e-12
L_PTL_G0_2|_RX|1 _PTL_G0_2|A_PTL _PTL_G0_2|_RX|1  1.346e-12
L_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|4  6.348e-12
L_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7  5.197e-12
L_PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7 _PTL_G0_2|A_PTL_RX  2.058e-12
L_PTL_G0_2|_RX|P1 _PTL_G0_2|_RX|2 0  4.795e-13
L_PTL_G0_2|_RX|P2 _PTL_G0_2|_RX|5 0  5.431e-13
L_PTL_G0_2|_RX|P3 _PTL_G0_2|_RX|8 0  5.339e-13
R_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|101  4.225701121488
R_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|104  3.429952209
R_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|107  2.7439617672
L_PTL_G0_2|_RX|RB1 _PTL_G0_2|_RX|101 0  2.38752113364072e-12
L_PTL_G0_2|_RX|RB2 _PTL_G0_2|_RX|104 0  1.937922998085e-12
L_PTL_G0_2|_RX|RB3 _PTL_G0_2|_RX|107 0  1.550338398468e-12
B_PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G0_2|_JTL|2 _PTL_G0_2|_JTL|6 _PTL_G0_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G0_2|_JTL|B1 0 _PTL_G0_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G0_2|_JTL|1 _PTL_G0_2|A_PTL_RX _PTL_G0_2|_JTL|1  2.067833848e-12
L_PTL_G0_2|_JTL|2 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|4  2.067833848e-12
L_PTL_G0_2|_JTL|3 _PTL_G0_2|_JTL|4 _PTL_G0_2|_JTL|6  2.067833848e-12
L_PTL_G0_2|_JTL|4 _PTL_G0_2|_JTL|6 G0_2_RX  2.067833848e-12
L_PTL_G0_2|_JTL|P1 _PTL_G0_2|_JTL|2 0  2e-13
L_PTL_G0_2|_JTL|P2 _PTL_G0_2|_JTL|7 0  2e-13
L_PTL_G0_2|_JTL|B1 _PTL_G0_2|_JTL|5 _PTL_G0_2|_JTL|4  2e-12
R_PTL_G0_2|_JTL|B1 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|3  2.7439617672
R_PTL_G0_2|_JTL|B2 _PTL_G0_2|_JTL|6 _PTL_G0_2|_JTL|8  2.7439617672
L_PTL_G0_2|_JTL|RB1 _PTL_G0_2|_JTL|3 0  1.750338398468e-12
L_PTL_G0_2|_JTL|RB2 _PTL_G0_2|_JTL|8 0  1.750338398468e-12
B_PTL_G1_2|_TX|1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|2 JJMIT AREA=2.5
B_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|5 JJMIT AREA=2.5
I_PTL_G1_2|_TX|B1 0 _PTL_G1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_2|_TX|B2 0 _PTL_G1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|3  1.684e-12
L_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|6  3.596e-12
L_PTL_G1_2|_TX|1 G1_2 _PTL_G1_2|_TX|1  2.063e-12
L_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|4  4.123e-12
L_PTL_G1_2|_TX|3 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|7  2.193e-12
R_PTL_G1_2|_TX|D _PTL_G1_2|_TX|7 _PTL_G1_2|A_PTL  1.36
L_PTL_G1_2|_TX|P1 _PTL_G1_2|_TX|2 0  5.254e-13
L_PTL_G1_2|_TX|P2 _PTL_G1_2|_TX|5 0  5.141e-13
R_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|101  2.7439617672
R_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|104  2.7439617672
L_PTL_G1_2|_TX|RB1 _PTL_G1_2|_TX|101 0  1.550338398468e-12
L_PTL_G1_2|_TX|RB2 _PTL_G1_2|_TX|104 0  1.550338398468e-12
B_PTL_G1_2|_RX|1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|5 JJMIT AREA=2.0
B_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|8 JJMIT AREA=2.5
I_PTL_G1_2|_RX|B1 0 _PTL_G1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|3  2.777e-12
I_PTL_G1_2|_RX|B2 0 _PTL_G1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|6  2.685e-12
I_PTL_G1_2|_RX|B3 0 _PTL_G1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|9  2.764e-12
L_PTL_G1_2|_RX|1 _PTL_G1_2|A_PTL _PTL_G1_2|_RX|1  1.346e-12
L_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|4  6.348e-12
L_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7  5.197e-12
L_PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7 _PTL_G1_2|A_PTL_RX  2.058e-12
L_PTL_G1_2|_RX|P1 _PTL_G1_2|_RX|2 0  4.795e-13
L_PTL_G1_2|_RX|P2 _PTL_G1_2|_RX|5 0  5.431e-13
L_PTL_G1_2|_RX|P3 _PTL_G1_2|_RX|8 0  5.339e-13
R_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|101  4.225701121488
R_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|104  3.429952209
R_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|107  2.7439617672
L_PTL_G1_2|_RX|RB1 _PTL_G1_2|_RX|101 0  2.38752113364072e-12
L_PTL_G1_2|_RX|RB2 _PTL_G1_2|_RX|104 0  1.937922998085e-12
L_PTL_G1_2|_RX|RB3 _PTL_G1_2|_RX|107 0  1.550338398468e-12
B_PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G1_2|_JTL|2 _PTL_G1_2|_JTL|6 _PTL_G1_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G1_2|_JTL|B1 0 _PTL_G1_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G1_2|_JTL|1 _PTL_G1_2|A_PTL_RX _PTL_G1_2|_JTL|1  2.067833848e-12
L_PTL_G1_2|_JTL|2 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|4  2.067833848e-12
L_PTL_G1_2|_JTL|3 _PTL_G1_2|_JTL|4 _PTL_G1_2|_JTL|6  2.067833848e-12
L_PTL_G1_2|_JTL|4 _PTL_G1_2|_JTL|6 G1_2_RX  2.067833848e-12
L_PTL_G1_2|_JTL|P1 _PTL_G1_2|_JTL|2 0  2e-13
L_PTL_G1_2|_JTL|P2 _PTL_G1_2|_JTL|7 0  2e-13
L_PTL_G1_2|_JTL|B1 _PTL_G1_2|_JTL|5 _PTL_G1_2|_JTL|4  2e-12
R_PTL_G1_2|_JTL|B1 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|3  2.7439617672
R_PTL_G1_2|_JTL|B2 _PTL_G1_2|_JTL|6 _PTL_G1_2|_JTL|8  2.7439617672
L_PTL_G1_2|_JTL|RB1 _PTL_G1_2|_JTL|3 0  1.750338398468e-12
L_PTL_G1_2|_JTL|RB2 _PTL_G1_2|_JTL|8 0  1.750338398468e-12
B_PTL_G2_2|_TX|1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|2 JJMIT AREA=2.5
B_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|5 JJMIT AREA=2.5
I_PTL_G2_2|_TX|B1 0 _PTL_G2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_2|_TX|B2 0 _PTL_G2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|3  1.684e-12
L_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|6  3.596e-12
L_PTL_G2_2|_TX|1 G2_2 _PTL_G2_2|_TX|1  2.063e-12
L_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|4  4.123e-12
L_PTL_G2_2|_TX|3 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|7  2.193e-12
R_PTL_G2_2|_TX|D _PTL_G2_2|_TX|7 _PTL_G2_2|A_PTL  1.36
L_PTL_G2_2|_TX|P1 _PTL_G2_2|_TX|2 0  5.254e-13
L_PTL_G2_2|_TX|P2 _PTL_G2_2|_TX|5 0  5.141e-13
R_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|101  2.7439617672
R_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|104  2.7439617672
L_PTL_G2_2|_TX|RB1 _PTL_G2_2|_TX|101 0  1.550338398468e-12
L_PTL_G2_2|_TX|RB2 _PTL_G2_2|_TX|104 0  1.550338398468e-12
B_PTL_G2_2|_RX|1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|5 JJMIT AREA=2.0
B_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|8 JJMIT AREA=2.5
I_PTL_G2_2|_RX|B1 0 _PTL_G2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|3  2.777e-12
I_PTL_G2_2|_RX|B2 0 _PTL_G2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|6  2.685e-12
I_PTL_G2_2|_RX|B3 0 _PTL_G2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|9  2.764e-12
L_PTL_G2_2|_RX|1 _PTL_G2_2|A_PTL _PTL_G2_2|_RX|1  1.346e-12
L_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|4  6.348e-12
L_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7  5.197e-12
L_PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7 _PTL_G2_2|A_PTL_RX  2.058e-12
L_PTL_G2_2|_RX|P1 _PTL_G2_2|_RX|2 0  4.795e-13
L_PTL_G2_2|_RX|P2 _PTL_G2_2|_RX|5 0  5.431e-13
L_PTL_G2_2|_RX|P3 _PTL_G2_2|_RX|8 0  5.339e-13
R_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|101  4.225701121488
R_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|104  3.429952209
R_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|107  2.7439617672
L_PTL_G2_2|_RX|RB1 _PTL_G2_2|_RX|101 0  2.38752113364072e-12
L_PTL_G2_2|_RX|RB2 _PTL_G2_2|_RX|104 0  1.937922998085e-12
L_PTL_G2_2|_RX|RB3 _PTL_G2_2|_RX|107 0  1.550338398468e-12
B_PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G2_2|_JTL|2 _PTL_G2_2|_JTL|6 _PTL_G2_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G2_2|_JTL|B1 0 _PTL_G2_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G2_2|_JTL|1 _PTL_G2_2|A_PTL_RX _PTL_G2_2|_JTL|1  2.067833848e-12
L_PTL_G2_2|_JTL|2 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|4  2.067833848e-12
L_PTL_G2_2|_JTL|3 _PTL_G2_2|_JTL|4 _PTL_G2_2|_JTL|6  2.067833848e-12
L_PTL_G2_2|_JTL|4 _PTL_G2_2|_JTL|6 G2_2_RX  2.067833848e-12
L_PTL_G2_2|_JTL|P1 _PTL_G2_2|_JTL|2 0  2e-13
L_PTL_G2_2|_JTL|P2 _PTL_G2_2|_JTL|7 0  2e-13
L_PTL_G2_2|_JTL|B1 _PTL_G2_2|_JTL|5 _PTL_G2_2|_JTL|4  2e-12
R_PTL_G2_2|_JTL|B1 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|3  2.7439617672
R_PTL_G2_2|_JTL|B2 _PTL_G2_2|_JTL|6 _PTL_G2_2|_JTL|8  2.7439617672
L_PTL_G2_2|_JTL|RB1 _PTL_G2_2|_JTL|3 0  1.750338398468e-12
L_PTL_G2_2|_JTL|RB2 _PTL_G2_2|_JTL|8 0  1.750338398468e-12
B_PTL_G3_2|_TX|1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|2 JJMIT AREA=2.5
B_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|5 JJMIT AREA=2.5
I_PTL_G3_2|_TX|B1 0 _PTL_G3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_2|_TX|B2 0 _PTL_G3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|3  1.684e-12
L_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|6  3.596e-12
L_PTL_G3_2|_TX|1 G3_2 _PTL_G3_2|_TX|1  2.063e-12
L_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|4  4.123e-12
L_PTL_G3_2|_TX|3 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|7  2.193e-12
R_PTL_G3_2|_TX|D _PTL_G3_2|_TX|7 _PTL_G3_2|A_PTL  1.36
L_PTL_G3_2|_TX|P1 _PTL_G3_2|_TX|2 0  5.254e-13
L_PTL_G3_2|_TX|P2 _PTL_G3_2|_TX|5 0  5.141e-13
R_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|101  2.7439617672
R_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|104  2.7439617672
L_PTL_G3_2|_TX|RB1 _PTL_G3_2|_TX|101 0  1.550338398468e-12
L_PTL_G3_2|_TX|RB2 _PTL_G3_2|_TX|104 0  1.550338398468e-12
B_PTL_G3_2|_RX|1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|5 JJMIT AREA=2.0
B_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|8 JJMIT AREA=2.5
I_PTL_G3_2|_RX|B1 0 _PTL_G3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|3  2.777e-12
I_PTL_G3_2|_RX|B2 0 _PTL_G3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|6  2.685e-12
I_PTL_G3_2|_RX|B3 0 _PTL_G3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|9  2.764e-12
L_PTL_G3_2|_RX|1 _PTL_G3_2|A_PTL _PTL_G3_2|_RX|1  1.346e-12
L_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|4  6.348e-12
L_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7  5.197e-12
L_PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7 _PTL_G3_2|A_PTL_RX  2.058e-12
L_PTL_G3_2|_RX|P1 _PTL_G3_2|_RX|2 0  4.795e-13
L_PTL_G3_2|_RX|P2 _PTL_G3_2|_RX|5 0  5.431e-13
L_PTL_G3_2|_RX|P3 _PTL_G3_2|_RX|8 0  5.339e-13
R_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|101  4.225701121488
R_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|104  3.429952209
R_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|107  2.7439617672
L_PTL_G3_2|_RX|RB1 _PTL_G3_2|_RX|101 0  2.38752113364072e-12
L_PTL_G3_2|_RX|RB2 _PTL_G3_2|_RX|104 0  1.937922998085e-12
L_PTL_G3_2|_RX|RB3 _PTL_G3_2|_RX|107 0  1.550338398468e-12
B_PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G3_2|_JTL|2 _PTL_G3_2|_JTL|6 _PTL_G3_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G3_2|_JTL|B1 0 _PTL_G3_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G3_2|_JTL|1 _PTL_G3_2|A_PTL_RX _PTL_G3_2|_JTL|1  2.067833848e-12
L_PTL_G3_2|_JTL|2 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|4  2.067833848e-12
L_PTL_G3_2|_JTL|3 _PTL_G3_2|_JTL|4 _PTL_G3_2|_JTL|6  2.067833848e-12
L_PTL_G3_2|_JTL|4 _PTL_G3_2|_JTL|6 G3_2_RX  2.067833848e-12
L_PTL_G3_2|_JTL|P1 _PTL_G3_2|_JTL|2 0  2e-13
L_PTL_G3_2|_JTL|P2 _PTL_G3_2|_JTL|7 0  2e-13
L_PTL_G3_2|_JTL|B1 _PTL_G3_2|_JTL|5 _PTL_G3_2|_JTL|4  2e-12
R_PTL_G3_2|_JTL|B1 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|3  2.7439617672
R_PTL_G3_2|_JTL|B2 _PTL_G3_2|_JTL|6 _PTL_G3_2|_JTL|8  2.7439617672
L_PTL_G3_2|_JTL|RB1 _PTL_G3_2|_JTL|3 0  1.750338398468e-12
L_PTL_G3_2|_JTL|RB2 _PTL_G3_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_2|_TX|B1 0 _PTL_IP1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_2|_TX|B2 0 _PTL_IP1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|3  1.684e-12
L_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|6  3.596e-12
L_PTL_IP1_2|_TX|1 IP1_2_OUT _PTL_IP1_2|_TX|1  2.063e-12
L_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|4  4.123e-12
L_PTL_IP1_2|_TX|3 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|7  2.193e-12
R_PTL_IP1_2|_TX|D _PTL_IP1_2|_TX|7 _PTL_IP1_2|A_PTL  1.36
L_PTL_IP1_2|_TX|P1 _PTL_IP1_2|_TX|2 0  5.254e-13
L_PTL_IP1_2|_TX|P2 _PTL_IP1_2|_TX|5 0  5.141e-13
R_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|101  2.7439617672
R_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|104  2.7439617672
L_PTL_IP1_2|_TX|RB1 _PTL_IP1_2|_TX|101 0  1.550338398468e-12
L_PTL_IP1_2|_TX|RB2 _PTL_IP1_2|_TX|104 0  1.550338398468e-12
B_PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_2|_RX|B1 0 _PTL_IP1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|3  2.777e-12
I_PTL_IP1_2|_RX|B2 0 _PTL_IP1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|6  2.685e-12
I_PTL_IP1_2|_RX|B3 0 _PTL_IP1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|9  2.764e-12
L_PTL_IP1_2|_RX|1 _PTL_IP1_2|A_PTL _PTL_IP1_2|_RX|1  1.346e-12
L_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|4  6.348e-12
L_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7  5.197e-12
L_PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7 _PTL_IP1_2|A_PTL_RX  2.058e-12
L_PTL_IP1_2|_RX|P1 _PTL_IP1_2|_RX|2 0  4.795e-13
L_PTL_IP1_2|_RX|P2 _PTL_IP1_2|_RX|5 0  5.431e-13
L_PTL_IP1_2|_RX|P3 _PTL_IP1_2|_RX|8 0  5.339e-13
R_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|101  4.225701121488
R_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|104  3.429952209
R_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|107  2.7439617672
L_PTL_IP1_2|_RX|RB1 _PTL_IP1_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_2|_RX|RB2 _PTL_IP1_2|_RX|104 0  1.937922998085e-12
L_PTL_IP1_2|_RX|RB3 _PTL_IP1_2|_RX|107 0  1.550338398468e-12
B_PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP1_2|_JTL|2 _PTL_IP1_2|_JTL|6 _PTL_IP1_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP1_2|_JTL|B1 0 _PTL_IP1_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP1_2|_JTL|1 _PTL_IP1_2|A_PTL_RX _PTL_IP1_2|_JTL|1  2.067833848e-12
L_PTL_IP1_2|_JTL|2 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|4  2.067833848e-12
L_PTL_IP1_2|_JTL|3 _PTL_IP1_2|_JTL|4 _PTL_IP1_2|_JTL|6  2.067833848e-12
L_PTL_IP1_2|_JTL|4 _PTL_IP1_2|_JTL|6 IP1_2_OUT_RX  2.067833848e-12
L_PTL_IP1_2|_JTL|P1 _PTL_IP1_2|_JTL|2 0  2e-13
L_PTL_IP1_2|_JTL|P2 _PTL_IP1_2|_JTL|7 0  2e-13
L_PTL_IP1_2|_JTL|B1 _PTL_IP1_2|_JTL|5 _PTL_IP1_2|_JTL|4  2e-12
R_PTL_IP1_2|_JTL|B1 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|3  2.7439617672
R_PTL_IP1_2|_JTL|B2 _PTL_IP1_2|_JTL|6 _PTL_IP1_2|_JTL|8  2.7439617672
L_PTL_IP1_2|_JTL|RB1 _PTL_IP1_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP1_2|_JTL|RB2 _PTL_IP1_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_2|_TX|B1 0 _PTL_IP2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_2|_TX|B2 0 _PTL_IP2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|3  1.684e-12
L_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|6  3.596e-12
L_PTL_IP2_2|_TX|1 IP2_2_OUT _PTL_IP2_2|_TX|1  2.063e-12
L_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|4  4.123e-12
L_PTL_IP2_2|_TX|3 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|7  2.193e-12
R_PTL_IP2_2|_TX|D _PTL_IP2_2|_TX|7 _PTL_IP2_2|A_PTL  1.36
L_PTL_IP2_2|_TX|P1 _PTL_IP2_2|_TX|2 0  5.254e-13
L_PTL_IP2_2|_TX|P2 _PTL_IP2_2|_TX|5 0  5.141e-13
R_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|101  2.7439617672
R_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|104  2.7439617672
L_PTL_IP2_2|_TX|RB1 _PTL_IP2_2|_TX|101 0  1.550338398468e-12
L_PTL_IP2_2|_TX|RB2 _PTL_IP2_2|_TX|104 0  1.550338398468e-12
B_PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_2|_RX|B1 0 _PTL_IP2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|3  2.777e-12
I_PTL_IP2_2|_RX|B2 0 _PTL_IP2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|6  2.685e-12
I_PTL_IP2_2|_RX|B3 0 _PTL_IP2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|9  2.764e-12
L_PTL_IP2_2|_RX|1 _PTL_IP2_2|A_PTL _PTL_IP2_2|_RX|1  1.346e-12
L_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|4  6.348e-12
L_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7  5.197e-12
L_PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7 _PTL_IP2_2|A_PTL_RX  2.058e-12
L_PTL_IP2_2|_RX|P1 _PTL_IP2_2|_RX|2 0  4.795e-13
L_PTL_IP2_2|_RX|P2 _PTL_IP2_2|_RX|5 0  5.431e-13
L_PTL_IP2_2|_RX|P3 _PTL_IP2_2|_RX|8 0  5.339e-13
R_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|101  4.225701121488
R_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|104  3.429952209
R_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|107  2.7439617672
L_PTL_IP2_2|_RX|RB1 _PTL_IP2_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_2|_RX|RB2 _PTL_IP2_2|_RX|104 0  1.937922998085e-12
L_PTL_IP2_2|_RX|RB3 _PTL_IP2_2|_RX|107 0  1.550338398468e-12
B_PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP2_2|_JTL|2 _PTL_IP2_2|_JTL|6 _PTL_IP2_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP2_2|_JTL|B1 0 _PTL_IP2_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP2_2|_JTL|1 _PTL_IP2_2|A_PTL_RX _PTL_IP2_2|_JTL|1  2.067833848e-12
L_PTL_IP2_2|_JTL|2 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|4  2.067833848e-12
L_PTL_IP2_2|_JTL|3 _PTL_IP2_2|_JTL|4 _PTL_IP2_2|_JTL|6  2.067833848e-12
L_PTL_IP2_2|_JTL|4 _PTL_IP2_2|_JTL|6 IP2_2_OUT_RX  2.067833848e-12
L_PTL_IP2_2|_JTL|P1 _PTL_IP2_2|_JTL|2 0  2e-13
L_PTL_IP2_2|_JTL|P2 _PTL_IP2_2|_JTL|7 0  2e-13
L_PTL_IP2_2|_JTL|B1 _PTL_IP2_2|_JTL|5 _PTL_IP2_2|_JTL|4  2e-12
R_PTL_IP2_2|_JTL|B1 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|3  2.7439617672
R_PTL_IP2_2|_JTL|B2 _PTL_IP2_2|_JTL|6 _PTL_IP2_2|_JTL|8  2.7439617672
L_PTL_IP2_2|_JTL|RB1 _PTL_IP2_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP2_2|_JTL|RB2 _PTL_IP2_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_2|_TX|B1 0 _PTL_IP3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_2|_TX|B2 0 _PTL_IP3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|3  1.684e-12
L_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|6  3.596e-12
L_PTL_IP3_2|_TX|1 IP3_2_OUT _PTL_IP3_2|_TX|1  2.063e-12
L_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|4  4.123e-12
L_PTL_IP3_2|_TX|3 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|7  2.193e-12
R_PTL_IP3_2|_TX|D _PTL_IP3_2|_TX|7 _PTL_IP3_2|A_PTL  1.36
L_PTL_IP3_2|_TX|P1 _PTL_IP3_2|_TX|2 0  5.254e-13
L_PTL_IP3_2|_TX|P2 _PTL_IP3_2|_TX|5 0  5.141e-13
R_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|101  2.7439617672
R_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|104  2.7439617672
L_PTL_IP3_2|_TX|RB1 _PTL_IP3_2|_TX|101 0  1.550338398468e-12
L_PTL_IP3_2|_TX|RB2 _PTL_IP3_2|_TX|104 0  1.550338398468e-12
B_PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_2|_RX|B1 0 _PTL_IP3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|3  2.777e-12
I_PTL_IP3_2|_RX|B2 0 _PTL_IP3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|6  2.685e-12
I_PTL_IP3_2|_RX|B3 0 _PTL_IP3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|9  2.764e-12
L_PTL_IP3_2|_RX|1 _PTL_IP3_2|A_PTL _PTL_IP3_2|_RX|1  1.346e-12
L_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|4  6.348e-12
L_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7  5.197e-12
L_PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7 _PTL_IP3_2|A_PTL_RX  2.058e-12
L_PTL_IP3_2|_RX|P1 _PTL_IP3_2|_RX|2 0  4.795e-13
L_PTL_IP3_2|_RX|P2 _PTL_IP3_2|_RX|5 0  5.431e-13
L_PTL_IP3_2|_RX|P3 _PTL_IP3_2|_RX|8 0  5.339e-13
R_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|101  4.225701121488
R_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|104  3.429952209
R_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|107  2.7439617672
L_PTL_IP3_2|_RX|RB1 _PTL_IP3_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_2|_RX|RB2 _PTL_IP3_2|_RX|104 0  1.937922998085e-12
L_PTL_IP3_2|_RX|RB3 _PTL_IP3_2|_RX|107 0  1.550338398468e-12
B_PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP3_2|_JTL|2 _PTL_IP3_2|_JTL|6 _PTL_IP3_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP3_2|_JTL|B1 0 _PTL_IP3_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP3_2|_JTL|1 _PTL_IP3_2|A_PTL_RX _PTL_IP3_2|_JTL|1  2.067833848e-12
L_PTL_IP3_2|_JTL|2 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|4  2.067833848e-12
L_PTL_IP3_2|_JTL|3 _PTL_IP3_2|_JTL|4 _PTL_IP3_2|_JTL|6  2.067833848e-12
L_PTL_IP3_2|_JTL|4 _PTL_IP3_2|_JTL|6 IP3_2_OUT_RX  2.067833848e-12
L_PTL_IP3_2|_JTL|P1 _PTL_IP3_2|_JTL|2 0  2e-13
L_PTL_IP3_2|_JTL|P2 _PTL_IP3_2|_JTL|7 0  2e-13
L_PTL_IP3_2|_JTL|B1 _PTL_IP3_2|_JTL|5 _PTL_IP3_2|_JTL|4  2e-12
R_PTL_IP3_2|_JTL|B1 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|3  2.7439617672
R_PTL_IP3_2|_JTL|B2 _PTL_IP3_2|_JTL|6 _PTL_IP3_2|_JTL|8  2.7439617672
L_PTL_IP3_2|_JTL|RB1 _PTL_IP3_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP3_2|_JTL|RB2 _PTL_IP3_2|_JTL|8 0  1.750338398468e-12
L_S0|I_1|B _S0|A1 _S0|I_1|MID  2e-12
I_S0|I_1|B 0 _S0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_3|B _S0|A3 _S0|I_3|MID  2e-12
I_S0|I_3|B 0 _S0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0|I_T|B _S0|T1 _S0|I_T|MID  2e-12
I_S0|I_T|B 0 _S0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_6|B _S0|Q1 _S0|I_6|MID  2e-12
I_S0|I_6|B 0 _S0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0|1|1 _S0|A1 _S0|1|MID_SERIES JJMIT AREA=2.5
L_S0|1|P _S0|1|MID_SERIES 0  2e-13
R_S0|1|B _S0|A1 _S0|1|MID_SHUNT  2.7439617672
L_S0|1|RB _S0|1|MID_SHUNT 0  1.550338398468e-12
B_S0|23|1 _S0|A2 _S0|A3 JJMIT AREA=1.7857142857142858
R_S0|23|B _S0|A2 _S0|23|MID_SHUNT  3.84154647408
L_S0|23|RB _S0|23|MID_SHUNT _S0|A3  2.1704737578552e-12
B_S0|3|1 _S0|A3 _S0|3|MID_SERIES JJMIT AREA=2.5
L_S0|3|P _S0|3|MID_SERIES 0  2e-13
R_S0|3|B _S0|A3 _S0|3|MID_SHUNT  2.7439617672
L_S0|3|RB _S0|3|MID_SHUNT 0  1.550338398468e-12
B_S0|4|1 _S0|A4 _S0|4|MID_SERIES JJMIT AREA=2.5
L_S0|4|P _S0|4|MID_SERIES 0  2e-13
R_S0|4|B _S0|A4 _S0|4|MID_SHUNT  2.7439617672
L_S0|4|RB _S0|4|MID_SHUNT 0  1.550338398468e-12
B_S0|T|1 _S0|T1 _S0|T|MID_SERIES JJMIT AREA=2.5
L_S0|T|P _S0|T|MID_SERIES 0  2e-13
R_S0|T|B _S0|T1 _S0|T|MID_SHUNT  2.7439617672
L_S0|T|RB _S0|T|MID_SHUNT 0  1.550338398468e-12
B_S0|45|1 _S0|T2 _S0|A4 JJMIT AREA=1.7857142857142858
R_S0|45|B _S0|T2 _S0|45|MID_SHUNT  3.84154647408
L_S0|45|RB _S0|45|MID_SHUNT _S0|A4  2.1704737578552e-12
B_S0|6|1 _S0|Q1 _S0|6|MID_SERIES JJMIT AREA=2.5
L_S0|6|P _S0|6|MID_SERIES 0  2e-13
R_S0|6|B _S0|Q1 _S0|6|MID_SHUNT  2.7439617672
L_S0|6|RB _S0|6|MID_SHUNT 0  1.550338398468e-12
L_S1|I_A1|B _S1|A1 _S1|I_A1|MID  2e-12
I_S1|I_A1|B 0 _S1|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_A3|B _S1|A3 _S1|I_A3|MID  2e-12
I_S1|I_A3|B 0 _S1|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B1|B _S1|B1 _S1|I_B1|MID  2e-12
I_S1|I_B1|B 0 _S1|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B3|B _S1|B3 _S1|I_B3|MID  2e-12
I_S1|I_B3|B 0 _S1|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_Q1|B _S1|Q1 _S1|I_Q1|MID  2e-12
I_S1|I_Q1|B 0 _S1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S1|A1|1 _S1|A1 _S1|A1|MID_SERIES JJMIT AREA=2.5
L_S1|A1|P _S1|A1|MID_SERIES 0  5e-13
R_S1|A1|B _S1|A1 _S1|A1|MID_SHUNT  2.7439617672
L_S1|A1|RB _S1|A1|MID_SHUNT 0  2.050338398468e-12
B_S1|A2|1 _S1|A2 _S1|A2|MID_SERIES JJMIT AREA=2.5
L_S1|A2|P _S1|A2|MID_SERIES 0  5e-13
R_S1|A2|B _S1|A2 _S1|A2|MID_SHUNT  2.7439617672
L_S1|A2|RB _S1|A2|MID_SHUNT 0  2.050338398468e-12
B_S1|A3|1 _S1|A2 _S1|A3|MID_SERIES JJMIT AREA=2.5
L_S1|A3|P _S1|A3|MID_SERIES _S1|A3  1.2e-12
R_S1|A3|B _S1|A2 _S1|A3|MID_SHUNT  2.7439617672
L_S1|A3|RB _S1|A3|MID_SHUNT _S1|A3  2.050338398468e-12
B_S1|B1|1 _S1|B1 _S1|B1|MID_SERIES JJMIT AREA=2.5
L_S1|B1|P _S1|B1|MID_SERIES 0  5e-13
R_S1|B1|B _S1|B1 _S1|B1|MID_SHUNT  2.7439617672
L_S1|B1|RB _S1|B1|MID_SHUNT 0  2.050338398468e-12
B_S1|B2|1 _S1|B2 _S1|B2|MID_SERIES JJMIT AREA=2.5
L_S1|B2|P _S1|B2|MID_SERIES 0  5e-13
R_S1|B2|B _S1|B2 _S1|B2|MID_SHUNT  2.7439617672
L_S1|B2|RB _S1|B2|MID_SHUNT 0  2.050338398468e-12
B_S1|B3|1 _S1|B2 _S1|B3|MID_SERIES JJMIT AREA=2.5
L_S1|B3|P _S1|B3|MID_SERIES _S1|B3  1.2e-12
R_S1|B3|B _S1|B2 _S1|B3|MID_SHUNT  2.7439617672
L_S1|B3|RB _S1|B3|MID_SHUNT _S1|B3  2.050338398468e-12
B_S1|T1|1 _S1|T1 _S1|T1|MID_SERIES JJMIT AREA=2.5
L_S1|T1|P _S1|T1|MID_SERIES 0  5e-13
R_S1|T1|B _S1|T1 _S1|T1|MID_SHUNT  2.7439617672
L_S1|T1|RB _S1|T1|MID_SHUNT 0  2.050338398468e-12
B_S1|T2|1 _S1|T2 _S1|ABTQ JJMIT AREA=2.0
R_S1|T2|B _S1|T2 _S1|T2|MID_SHUNT  3.429952209
L_S1|T2|RB _S1|T2|MID_SHUNT _S1|ABTQ  2.437922998085e-12
B_S1|AB|1 _S1|AB _S1|AB|MID_SERIES JJMIT AREA=1.5
L_S1|AB|P _S1|AB|MID_SERIES _S1|ABTQ  1.2e-12
R_S1|AB|B _S1|AB _S1|AB|MID_SHUNT  4.573269612
L_S1|AB|RB _S1|AB|MID_SHUNT _S1|ABTQ  3.08389733078e-12
B_S1|ABTQ|1 _S1|ABTQ _S1|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S1|ABTQ|P _S1|ABTQ|MID_SERIES 0  5e-13
R_S1|ABTQ|B _S1|ABTQ _S1|ABTQ|MID_SHUNT  3.6586156896
L_S1|ABTQ|RB _S1|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S1|Q1|1 _S1|Q1 _S1|Q1|MID_SERIES JJMIT AREA=2.5
L_S1|Q1|P _S1|Q1|MID_SERIES 0  5e-13
R_S1|Q1|B _S1|Q1 _S1|Q1|MID_SHUNT  2.7439617672
L_S1|Q1|RB _S1|Q1|MID_SHUNT 0  2.050338398468e-12
L_S2|I_A1|B _S2|A1 _S2|I_A1|MID  2e-12
I_S2|I_A1|B 0 _S2|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_A3|B _S2|A3 _S2|I_A3|MID  2e-12
I_S2|I_A3|B 0 _S2|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B1|B _S2|B1 _S2|I_B1|MID  2e-12
I_S2|I_B1|B 0 _S2|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B3|B _S2|B3 _S2|I_B3|MID  2e-12
I_S2|I_B3|B 0 _S2|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_Q1|B _S2|Q1 _S2|I_Q1|MID  2e-12
I_S2|I_Q1|B 0 _S2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S2|A1|1 _S2|A1 _S2|A1|MID_SERIES JJMIT AREA=2.5
L_S2|A1|P _S2|A1|MID_SERIES 0  5e-13
R_S2|A1|B _S2|A1 _S2|A1|MID_SHUNT  2.7439617672
L_S2|A1|RB _S2|A1|MID_SHUNT 0  2.050338398468e-12
B_S2|A2|1 _S2|A2 _S2|A2|MID_SERIES JJMIT AREA=2.5
L_S2|A2|P _S2|A2|MID_SERIES 0  5e-13
R_S2|A2|B _S2|A2 _S2|A2|MID_SHUNT  2.7439617672
L_S2|A2|RB _S2|A2|MID_SHUNT 0  2.050338398468e-12
B_S2|A3|1 _S2|A2 _S2|A3|MID_SERIES JJMIT AREA=2.5
L_S2|A3|P _S2|A3|MID_SERIES _S2|A3  1.2e-12
R_S2|A3|B _S2|A2 _S2|A3|MID_SHUNT  2.7439617672
L_S2|A3|RB _S2|A3|MID_SHUNT _S2|A3  2.050338398468e-12
B_S2|B1|1 _S2|B1 _S2|B1|MID_SERIES JJMIT AREA=2.5
L_S2|B1|P _S2|B1|MID_SERIES 0  5e-13
R_S2|B1|B _S2|B1 _S2|B1|MID_SHUNT  2.7439617672
L_S2|B1|RB _S2|B1|MID_SHUNT 0  2.050338398468e-12
B_S2|B2|1 _S2|B2 _S2|B2|MID_SERIES JJMIT AREA=2.5
L_S2|B2|P _S2|B2|MID_SERIES 0  5e-13
R_S2|B2|B _S2|B2 _S2|B2|MID_SHUNT  2.7439617672
L_S2|B2|RB _S2|B2|MID_SHUNT 0  2.050338398468e-12
B_S2|B3|1 _S2|B2 _S2|B3|MID_SERIES JJMIT AREA=2.5
L_S2|B3|P _S2|B3|MID_SERIES _S2|B3  1.2e-12
R_S2|B3|B _S2|B2 _S2|B3|MID_SHUNT  2.7439617672
L_S2|B3|RB _S2|B3|MID_SHUNT _S2|B3  2.050338398468e-12
B_S2|T1|1 _S2|T1 _S2|T1|MID_SERIES JJMIT AREA=2.5
L_S2|T1|P _S2|T1|MID_SERIES 0  5e-13
R_S2|T1|B _S2|T1 _S2|T1|MID_SHUNT  2.7439617672
L_S2|T1|RB _S2|T1|MID_SHUNT 0  2.050338398468e-12
B_S2|T2|1 _S2|T2 _S2|ABTQ JJMIT AREA=2.0
R_S2|T2|B _S2|T2 _S2|T2|MID_SHUNT  3.429952209
L_S2|T2|RB _S2|T2|MID_SHUNT _S2|ABTQ  2.437922998085e-12
B_S2|AB|1 _S2|AB _S2|AB|MID_SERIES JJMIT AREA=1.5
L_S2|AB|P _S2|AB|MID_SERIES _S2|ABTQ  1.2e-12
R_S2|AB|B _S2|AB _S2|AB|MID_SHUNT  4.573269612
L_S2|AB|RB _S2|AB|MID_SHUNT _S2|ABTQ  3.08389733078e-12
B_S2|ABTQ|1 _S2|ABTQ _S2|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S2|ABTQ|P _S2|ABTQ|MID_SERIES 0  5e-13
R_S2|ABTQ|B _S2|ABTQ _S2|ABTQ|MID_SHUNT  3.6586156896
L_S2|ABTQ|RB _S2|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S2|Q1|1 _S2|Q1 _S2|Q1|MID_SERIES JJMIT AREA=2.5
L_S2|Q1|P _S2|Q1|MID_SERIES 0  5e-13
R_S2|Q1|B _S2|Q1 _S2|Q1|MID_SHUNT  2.7439617672
L_S2|Q1|RB _S2|Q1|MID_SHUNT 0  2.050338398468e-12
L_S3|I_A1|B _S3|A1 _S3|I_A1|MID  2e-12
I_S3|I_A1|B 0 _S3|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_A3|B _S3|A3 _S3|I_A3|MID  2e-12
I_S3|I_A3|B 0 _S3|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B1|B _S3|B1 _S3|I_B1|MID  2e-12
I_S3|I_B1|B 0 _S3|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B3|B _S3|B3 _S3|I_B3|MID  2e-12
I_S3|I_B3|B 0 _S3|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_Q1|B _S3|Q1 _S3|I_Q1|MID  2e-12
I_S3|I_Q1|B 0 _S3|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S3|A1|1 _S3|A1 _S3|A1|MID_SERIES JJMIT AREA=2.5
L_S3|A1|P _S3|A1|MID_SERIES 0  5e-13
R_S3|A1|B _S3|A1 _S3|A1|MID_SHUNT  2.7439617672
L_S3|A1|RB _S3|A1|MID_SHUNT 0  2.050338398468e-12
B_S3|A2|1 _S3|A2 _S3|A2|MID_SERIES JJMIT AREA=2.5
L_S3|A2|P _S3|A2|MID_SERIES 0  5e-13
R_S3|A2|B _S3|A2 _S3|A2|MID_SHUNT  2.7439617672
L_S3|A2|RB _S3|A2|MID_SHUNT 0  2.050338398468e-12
B_S3|A3|1 _S3|A2 _S3|A3|MID_SERIES JJMIT AREA=2.5
L_S3|A3|P _S3|A3|MID_SERIES _S3|A3  1.2e-12
R_S3|A3|B _S3|A2 _S3|A3|MID_SHUNT  2.7439617672
L_S3|A3|RB _S3|A3|MID_SHUNT _S3|A3  2.050338398468e-12
B_S3|B1|1 _S3|B1 _S3|B1|MID_SERIES JJMIT AREA=2.5
L_S3|B1|P _S3|B1|MID_SERIES 0  5e-13
R_S3|B1|B _S3|B1 _S3|B1|MID_SHUNT  2.7439617672
L_S3|B1|RB _S3|B1|MID_SHUNT 0  2.050338398468e-12
B_S3|B2|1 _S3|B2 _S3|B2|MID_SERIES JJMIT AREA=2.5
L_S3|B2|P _S3|B2|MID_SERIES 0  5e-13
R_S3|B2|B _S3|B2 _S3|B2|MID_SHUNT  2.7439617672
L_S3|B2|RB _S3|B2|MID_SHUNT 0  2.050338398468e-12
B_S3|B3|1 _S3|B2 _S3|B3|MID_SERIES JJMIT AREA=2.5
L_S3|B3|P _S3|B3|MID_SERIES _S3|B3  1.2e-12
R_S3|B3|B _S3|B2 _S3|B3|MID_SHUNT  2.7439617672
L_S3|B3|RB _S3|B3|MID_SHUNT _S3|B3  2.050338398468e-12
B_S3|T1|1 _S3|T1 _S3|T1|MID_SERIES JJMIT AREA=2.5
L_S3|T1|P _S3|T1|MID_SERIES 0  5e-13
R_S3|T1|B _S3|T1 _S3|T1|MID_SHUNT  2.7439617672
L_S3|T1|RB _S3|T1|MID_SHUNT 0  2.050338398468e-12
B_S3|T2|1 _S3|T2 _S3|ABTQ JJMIT AREA=2.0
R_S3|T2|B _S3|T2 _S3|T2|MID_SHUNT  3.429952209
L_S3|T2|RB _S3|T2|MID_SHUNT _S3|ABTQ  2.437922998085e-12
B_S3|AB|1 _S3|AB _S3|AB|MID_SERIES JJMIT AREA=1.5
L_S3|AB|P _S3|AB|MID_SERIES _S3|ABTQ  1.2e-12
R_S3|AB|B _S3|AB _S3|AB|MID_SHUNT  4.573269612
L_S3|AB|RB _S3|AB|MID_SHUNT _S3|ABTQ  3.08389733078e-12
B_S3|ABTQ|1 _S3|ABTQ _S3|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S3|ABTQ|P _S3|ABTQ|MID_SERIES 0  5e-13
R_S3|ABTQ|B _S3|ABTQ _S3|ABTQ|MID_SHUNT  3.6586156896
L_S3|ABTQ|RB _S3|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S3|Q1|1 _S3|Q1 _S3|Q1|MID_SERIES JJMIT AREA=2.5
L_S3|Q1|P _S3|Q1|MID_SERIES 0  5e-13
R_S3|Q1|B _S3|Q1 _S3|Q1|MID_SHUNT  2.7439617672
L_S3|Q1|RB _S3|Q1|MID_SHUNT 0  2.050338398468e-12
L_S4|I_1|B _S4|A1 _S4|I_1|MID  2e-12
I_S4|I_1|B 0 _S4|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_3|B _S4|A3 _S4|I_3|MID  2e-12
I_S4|I_3|B 0 _S4|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S4|I_T|B _S4|T1 _S4|I_T|MID  2e-12
I_S4|I_T|B 0 _S4|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_6|B _S4|Q1 _S4|I_6|MID  2e-12
I_S4|I_6|B 0 _S4|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S4|1|1 _S4|A1 _S4|1|MID_SERIES JJMIT AREA=2.5
L_S4|1|P _S4|1|MID_SERIES 0  2e-13
R_S4|1|B _S4|A1 _S4|1|MID_SHUNT  2.7439617672
L_S4|1|RB _S4|1|MID_SHUNT 0  1.550338398468e-12
B_S4|23|1 _S4|A2 _S4|A3 JJMIT AREA=1.7857142857142858
R_S4|23|B _S4|A2 _S4|23|MID_SHUNT  3.84154647408
L_S4|23|RB _S4|23|MID_SHUNT _S4|A3  2.1704737578552e-12
B_S4|3|1 _S4|A3 _S4|3|MID_SERIES JJMIT AREA=2.5
L_S4|3|P _S4|3|MID_SERIES 0  2e-13
R_S4|3|B _S4|A3 _S4|3|MID_SHUNT  2.7439617672
L_S4|3|RB _S4|3|MID_SHUNT 0  1.550338398468e-12
B_S4|4|1 _S4|A4 _S4|4|MID_SERIES JJMIT AREA=2.5
L_S4|4|P _S4|4|MID_SERIES 0  2e-13
R_S4|4|B _S4|A4 _S4|4|MID_SHUNT  2.7439617672
L_S4|4|RB _S4|4|MID_SHUNT 0  1.550338398468e-12
B_S4|T|1 _S4|T1 _S4|T|MID_SERIES JJMIT AREA=2.5
L_S4|T|P _S4|T|MID_SERIES 0  2e-13
R_S4|T|B _S4|T1 _S4|T|MID_SHUNT  2.7439617672
L_S4|T|RB _S4|T|MID_SHUNT 0  1.550338398468e-12
B_S4|45|1 _S4|T2 _S4|A4 JJMIT AREA=1.7857142857142858
R_S4|45|B _S4|T2 _S4|45|MID_SHUNT  3.84154647408
L_S4|45|RB _S4|45|MID_SHUNT _S4|A4  2.1704737578552e-12
B_S4|6|1 _S4|Q1 _S4|6|MID_SERIES JJMIT AREA=2.5
L_S4|6|P _S4|6|MID_SERIES 0  2e-13
R_S4|6|B _S4|Q1 _S4|6|MID_SHUNT  2.7439617672
L_S4|6|RB _S4|6|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_A|I_D1|B I0|_SPL_A|D1 I0|_SPL_A|I_D1|MID  2e-12
II0|_SPL_A|I_D1|B 0 I0|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_D2|B I0|_SPL_A|D2 I0|_SPL_A|I_D2|MID  2e-12
II0|_SPL_A|I_D2|B 0 I0|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_A|I_Q1|B I0|_SPL_A|QA1 I0|_SPL_A|I_Q1|MID  2e-12
II0|_SPL_A|I_Q1|B 0 I0|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_Q2|B I0|_SPL_A|QB1 I0|_SPL_A|I_Q2|MID  2e-12
II0|_SPL_A|I_Q2|B 0 I0|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_A|1|1 I0|_SPL_A|D1 I0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|1|P I0|_SPL_A|1|MID_SERIES 0  2e-13
RI0|_SPL_A|1|B I0|_SPL_A|D1 I0|_SPL_A|1|MID_SHUNT  2.7439617672
LI0|_SPL_A|1|RB I0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|2|1 I0|_SPL_A|D2 I0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|2|P I0|_SPL_A|2|MID_SERIES 0  2e-13
RI0|_SPL_A|2|B I0|_SPL_A|D2 I0|_SPL_A|2|MID_SHUNT  2.7439617672
LI0|_SPL_A|2|RB I0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|A|1 I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|A|P I0|_SPL_A|A|MID_SERIES 0  2e-13
RI0|_SPL_A|A|B I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SHUNT  2.7439617672
LI0|_SPL_A|A|RB I0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|B|1 I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|B|P I0|_SPL_A|B|MID_SERIES 0  2e-13
RI0|_SPL_A|B|B I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SHUNT  2.7439617672
LI0|_SPL_A|B|RB I0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_B|I_D1|B I0|_SPL_B|D1 I0|_SPL_B|I_D1|MID  2e-12
II0|_SPL_B|I_D1|B 0 I0|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_D2|B I0|_SPL_B|D2 I0|_SPL_B|I_D2|MID  2e-12
II0|_SPL_B|I_D2|B 0 I0|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_B|I_Q1|B I0|_SPL_B|QA1 I0|_SPL_B|I_Q1|MID  2e-12
II0|_SPL_B|I_Q1|B 0 I0|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_Q2|B I0|_SPL_B|QB1 I0|_SPL_B|I_Q2|MID  2e-12
II0|_SPL_B|I_Q2|B 0 I0|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_B|1|1 I0|_SPL_B|D1 I0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|1|P I0|_SPL_B|1|MID_SERIES 0  2e-13
RI0|_SPL_B|1|B I0|_SPL_B|D1 I0|_SPL_B|1|MID_SHUNT  2.7439617672
LI0|_SPL_B|1|RB I0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|2|1 I0|_SPL_B|D2 I0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|2|P I0|_SPL_B|2|MID_SERIES 0  2e-13
RI0|_SPL_B|2|B I0|_SPL_B|D2 I0|_SPL_B|2|MID_SHUNT  2.7439617672
LI0|_SPL_B|2|RB I0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|A|1 I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|A|P I0|_SPL_B|A|MID_SERIES 0  2e-13
RI0|_SPL_B|A|B I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SHUNT  2.7439617672
LI0|_SPL_B|A|RB I0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|B|1 I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|B|P I0|_SPL_B|B|MID_SERIES 0  2e-13
RI0|_SPL_B|B|B I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SHUNT  2.7439617672
LI0|_SPL_B|B|RB I0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_A|I_1|B I0|_DFF_A|A1 I0|_DFF_A|I_1|MID  2e-12
II0|_DFF_A|I_1|B 0 I0|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_3|B I0|_DFF_A|A3 I0|_DFF_A|I_3|MID  2e-12
II0|_DFF_A|I_3|B 0 I0|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_A|I_T|B I0|_DFF_A|T1 I0|_DFF_A|I_T|MID  2e-12
II0|_DFF_A|I_T|B 0 I0|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_6|B I0|_DFF_A|Q1 I0|_DFF_A|I_6|MID  2e-12
II0|_DFF_A|I_6|B 0 I0|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_A|1|1 I0|_DFF_A|A1 I0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|1|P I0|_DFF_A|1|MID_SERIES 0  2e-13
RI0|_DFF_A|1|B I0|_DFF_A|A1 I0|_DFF_A|1|MID_SHUNT  2.7439617672
LI0|_DFF_A|1|RB I0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|23|1 I0|_DFF_A|A2 I0|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|23|B I0|_DFF_A|A2 I0|_DFF_A|23|MID_SHUNT  3.84154647408
LI0|_DFF_A|23|RB I0|_DFF_A|23|MID_SHUNT I0|_DFF_A|A3  2.1704737578552e-12
BI0|_DFF_A|3|1 I0|_DFF_A|A3 I0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|3|P I0|_DFF_A|3|MID_SERIES 0  2e-13
RI0|_DFF_A|3|B I0|_DFF_A|A3 I0|_DFF_A|3|MID_SHUNT  2.7439617672
LI0|_DFF_A|3|RB I0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|4|1 I0|_DFF_A|A4 I0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|4|P I0|_DFF_A|4|MID_SERIES 0  2e-13
RI0|_DFF_A|4|B I0|_DFF_A|A4 I0|_DFF_A|4|MID_SHUNT  2.7439617672
LI0|_DFF_A|4|RB I0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|T|1 I0|_DFF_A|T1 I0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|T|P I0|_DFF_A|T|MID_SERIES 0  2e-13
RI0|_DFF_A|T|B I0|_DFF_A|T1 I0|_DFF_A|T|MID_SHUNT  2.7439617672
LI0|_DFF_A|T|RB I0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|45|1 I0|_DFF_A|T2 I0|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|45|B I0|_DFF_A|T2 I0|_DFF_A|45|MID_SHUNT  3.84154647408
LI0|_DFF_A|45|RB I0|_DFF_A|45|MID_SHUNT I0|_DFF_A|A4  2.1704737578552e-12
BI0|_DFF_A|6|1 I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|6|P I0|_DFF_A|6|MID_SERIES 0  2e-13
RI0|_DFF_A|6|B I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SHUNT  2.7439617672
LI0|_DFF_A|6|RB I0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_B|I_1|B I0|_DFF_B|A1 I0|_DFF_B|I_1|MID  2e-12
II0|_DFF_B|I_1|B 0 I0|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_3|B I0|_DFF_B|A3 I0|_DFF_B|I_3|MID  2e-12
II0|_DFF_B|I_3|B 0 I0|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_B|I_T|B I0|_DFF_B|T1 I0|_DFF_B|I_T|MID  2e-12
II0|_DFF_B|I_T|B 0 I0|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_6|B I0|_DFF_B|Q1 I0|_DFF_B|I_6|MID  2e-12
II0|_DFF_B|I_6|B 0 I0|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_B|1|1 I0|_DFF_B|A1 I0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|1|P I0|_DFF_B|1|MID_SERIES 0  2e-13
RI0|_DFF_B|1|B I0|_DFF_B|A1 I0|_DFF_B|1|MID_SHUNT  2.7439617672
LI0|_DFF_B|1|RB I0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|23|1 I0|_DFF_B|A2 I0|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|23|B I0|_DFF_B|A2 I0|_DFF_B|23|MID_SHUNT  3.84154647408
LI0|_DFF_B|23|RB I0|_DFF_B|23|MID_SHUNT I0|_DFF_B|A3  2.1704737578552e-12
BI0|_DFF_B|3|1 I0|_DFF_B|A3 I0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|3|P I0|_DFF_B|3|MID_SERIES 0  2e-13
RI0|_DFF_B|3|B I0|_DFF_B|A3 I0|_DFF_B|3|MID_SHUNT  2.7439617672
LI0|_DFF_B|3|RB I0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|4|1 I0|_DFF_B|A4 I0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|4|P I0|_DFF_B|4|MID_SERIES 0  2e-13
RI0|_DFF_B|4|B I0|_DFF_B|A4 I0|_DFF_B|4|MID_SHUNT  2.7439617672
LI0|_DFF_B|4|RB I0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|T|1 I0|_DFF_B|T1 I0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|T|P I0|_DFF_B|T|MID_SERIES 0  2e-13
RI0|_DFF_B|T|B I0|_DFF_B|T1 I0|_DFF_B|T|MID_SHUNT  2.7439617672
LI0|_DFF_B|T|RB I0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|45|1 I0|_DFF_B|T2 I0|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|45|B I0|_DFF_B|T2 I0|_DFF_B|45|MID_SHUNT  3.84154647408
LI0|_DFF_B|45|RB I0|_DFF_B|45|MID_SHUNT I0|_DFF_B|A4  2.1704737578552e-12
BI0|_DFF_B|6|1 I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|6|P I0|_DFF_B|6|MID_SERIES 0  2e-13
RI0|_DFF_B|6|B I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SHUNT  2.7439617672
LI0|_DFF_B|6|RB I0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI0|_XOR|I_A1|B I0|_XOR|A1 I0|_XOR|I_A1|MID  2e-12
II0|_XOR|I_A1|B 0 I0|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_A3|B I0|_XOR|A3 I0|_XOR|I_A3|MID  2e-12
II0|_XOR|I_A3|B 0 I0|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B1|B I0|_XOR|B1 I0|_XOR|I_B1|MID  2e-12
II0|_XOR|I_B1|B 0 I0|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B3|B I0|_XOR|B3 I0|_XOR|I_B3|MID  2e-12
II0|_XOR|I_B3|B 0 I0|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_Q1|B I0|_XOR|Q1 I0|_XOR|I_Q1|MID  2e-12
II0|_XOR|I_Q1|B 0 I0|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_XOR|A1|1 I0|_XOR|A1 I0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A1|P I0|_XOR|A1|MID_SERIES 0  5e-13
RI0|_XOR|A1|B I0|_XOR|A1 I0|_XOR|A1|MID_SHUNT  2.7439617672
LI0|_XOR|A1|RB I0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A2|1 I0|_XOR|A2 I0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A2|P I0|_XOR|A2|MID_SERIES 0  5e-13
RI0|_XOR|A2|B I0|_XOR|A2 I0|_XOR|A2|MID_SHUNT  2.7439617672
LI0|_XOR|A2|RB I0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A3|1 I0|_XOR|A2 I0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A3|P I0|_XOR|A3|MID_SERIES I0|_XOR|A3  1.2e-12
RI0|_XOR|A3|B I0|_XOR|A2 I0|_XOR|A3|MID_SHUNT  2.7439617672
LI0|_XOR|A3|RB I0|_XOR|A3|MID_SHUNT I0|_XOR|A3  2.050338398468e-12
BI0|_XOR|B1|1 I0|_XOR|B1 I0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B1|P I0|_XOR|B1|MID_SERIES 0  5e-13
RI0|_XOR|B1|B I0|_XOR|B1 I0|_XOR|B1|MID_SHUNT  2.7439617672
LI0|_XOR|B1|RB I0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B2|1 I0|_XOR|B2 I0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B2|P I0|_XOR|B2|MID_SERIES 0  5e-13
RI0|_XOR|B2|B I0|_XOR|B2 I0|_XOR|B2|MID_SHUNT  2.7439617672
LI0|_XOR|B2|RB I0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B3|1 I0|_XOR|B2 I0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B3|P I0|_XOR|B3|MID_SERIES I0|_XOR|B3  1.2e-12
RI0|_XOR|B3|B I0|_XOR|B2 I0|_XOR|B3|MID_SHUNT  2.7439617672
LI0|_XOR|B3|RB I0|_XOR|B3|MID_SHUNT I0|_XOR|B3  2.050338398468e-12
BI0|_XOR|T1|1 I0|_XOR|T1 I0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|T1|P I0|_XOR|T1|MID_SERIES 0  5e-13
RI0|_XOR|T1|B I0|_XOR|T1 I0|_XOR|T1|MID_SHUNT  2.7439617672
LI0|_XOR|T1|RB I0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|T2|1 I0|_XOR|T2 I0|_XOR|ABTQ JJMIT AREA=2.0
RI0|_XOR|T2|B I0|_XOR|T2 I0|_XOR|T2|MID_SHUNT  3.429952209
LI0|_XOR|T2|RB I0|_XOR|T2|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|AB|1 I0|_XOR|AB I0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI0|_XOR|AB|P I0|_XOR|AB|MID_SERIES I0|_XOR|ABTQ  1.2e-12
RI0|_XOR|AB|B I0|_XOR|AB I0|_XOR|AB|MID_SHUNT  3.429952209
LI0|_XOR|AB|RB I0|_XOR|AB|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|ABTQ|1 I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|ABTQ|P I0|_XOR|ABTQ|MID_SERIES 0  5e-13
RI0|_XOR|ABTQ|B I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI0|_XOR|ABTQ|RB I0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|Q1|1 I0|_XOR|Q1 I0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|Q1|P I0|_XOR|Q1|MID_SERIES 0  5e-13
RI0|_XOR|Q1|B I0|_XOR|Q1 I0|_XOR|Q1|MID_SHUNT  2.7439617672
LI0|_XOR|Q1|RB I0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI0|_AND|I_A1|B I0|_AND|A1 I0|_AND|I_A1|MID  2e-12
II0|_AND|I_A1|B 0 I0|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_B1|B I0|_AND|B1 I0|_AND|I_B1|MID  2e-12
II0|_AND|I_B1|B 0 I0|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q3|B I0|_AND|Q3 I0|_AND|I_Q3|MID  2e-12
II0|_AND|I_Q3|B 0 I0|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0|_AND|I_Q2|B I0|_AND|Q2 I0|_AND|I_Q2|MID  2e-12
II0|_AND|I_Q2|B 0 I0|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q1|B I0|_AND|Q1 I0|_AND|I_Q1|MID  2e-12
II0|_AND|I_Q1|B 0 I0|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_AND|A1|1 I0|_AND|A1 I0|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A1|P I0|_AND|A1|MID_SERIES 0  2e-13
RI0|_AND|A1|B I0|_AND|A1 I0|_AND|A1|MID_SHUNT  2.7439617672
LI0|_AND|A1|RB I0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A2|1 I0|_AND|A2 I0|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A2|P I0|_AND|A2|MID_SERIES 0  2e-13
RI0|_AND|A2|B I0|_AND|A2 I0|_AND|A2|MID_SHUNT  2.7439617672
LI0|_AND|A2|RB I0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A12|1 I0|_AND|A2 I0|_AND|A3 JJMIT AREA=1.7857142857142858
RI0|_AND|A12|B I0|_AND|A2 I0|_AND|A12|MID_SHUNT  3.84154647408
LI0|_AND|A12|RB I0|_AND|A12|MID_SHUNT I0|_AND|A3  2.1704737578552e-12
BI0|_AND|B1|1 I0|_AND|B1 I0|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B1|P I0|_AND|B1|MID_SERIES 0  2e-13
RI0|_AND|B1|B I0|_AND|B1 I0|_AND|B1|MID_SHUNT  2.7439617672
LI0|_AND|B1|RB I0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B2|1 I0|_AND|B2 I0|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B2|P I0|_AND|B2|MID_SERIES 0  2e-13
RI0|_AND|B2|B I0|_AND|B2 I0|_AND|B2|MID_SHUNT  2.7439617672
LI0|_AND|B2|RB I0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B12|1 I0|_AND|B2 I0|_AND|B3 JJMIT AREA=1.7857142857142858
RI0|_AND|B12|B I0|_AND|B2 I0|_AND|B12|MID_SHUNT  3.84154647408
LI0|_AND|B12|RB I0|_AND|B12|MID_SHUNT I0|_AND|B3  2.1704737578552e-12
BI0|_AND|Q2|1 I0|_AND|Q2 I0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q2|P I0|_AND|Q2|MID_SERIES 0  2e-13
RI0|_AND|Q2|B I0|_AND|Q2 I0|_AND|Q2|MID_SHUNT  2.7439617672
LI0|_AND|Q2|RB I0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|Q1|1 I0|_AND|Q1 I0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q1|P I0|_AND|Q1|MID_SERIES 0  2e-13
RI0|_AND|Q1|B I0|_AND|Q1 I0|_AND|Q1|MID_SHUNT  2.7439617672
LI0|_AND|Q1|RB I0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_A|I_D1|B I1|_SPL_A|D1 I1|_SPL_A|I_D1|MID  2e-12
II1|_SPL_A|I_D1|B 0 I1|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_D2|B I1|_SPL_A|D2 I1|_SPL_A|I_D2|MID  2e-12
II1|_SPL_A|I_D2|B 0 I1|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_A|I_Q1|B I1|_SPL_A|QA1 I1|_SPL_A|I_Q1|MID  2e-12
II1|_SPL_A|I_Q1|B 0 I1|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_Q2|B I1|_SPL_A|QB1 I1|_SPL_A|I_Q2|MID  2e-12
II1|_SPL_A|I_Q2|B 0 I1|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_A|1|1 I1|_SPL_A|D1 I1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|1|P I1|_SPL_A|1|MID_SERIES 0  2e-13
RI1|_SPL_A|1|B I1|_SPL_A|D1 I1|_SPL_A|1|MID_SHUNT  2.7439617672
LI1|_SPL_A|1|RB I1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|2|1 I1|_SPL_A|D2 I1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|2|P I1|_SPL_A|2|MID_SERIES 0  2e-13
RI1|_SPL_A|2|B I1|_SPL_A|D2 I1|_SPL_A|2|MID_SHUNT  2.7439617672
LI1|_SPL_A|2|RB I1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|A|1 I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|A|P I1|_SPL_A|A|MID_SERIES 0  2e-13
RI1|_SPL_A|A|B I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SHUNT  2.7439617672
LI1|_SPL_A|A|RB I1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|B|1 I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|B|P I1|_SPL_A|B|MID_SERIES 0  2e-13
RI1|_SPL_A|B|B I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SHUNT  2.7439617672
LI1|_SPL_A|B|RB I1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_B|I_D1|B I1|_SPL_B|D1 I1|_SPL_B|I_D1|MID  2e-12
II1|_SPL_B|I_D1|B 0 I1|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_D2|B I1|_SPL_B|D2 I1|_SPL_B|I_D2|MID  2e-12
II1|_SPL_B|I_D2|B 0 I1|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_B|I_Q1|B I1|_SPL_B|QA1 I1|_SPL_B|I_Q1|MID  2e-12
II1|_SPL_B|I_Q1|B 0 I1|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_Q2|B I1|_SPL_B|QB1 I1|_SPL_B|I_Q2|MID  2e-12
II1|_SPL_B|I_Q2|B 0 I1|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_B|1|1 I1|_SPL_B|D1 I1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|1|P I1|_SPL_B|1|MID_SERIES 0  2e-13
RI1|_SPL_B|1|B I1|_SPL_B|D1 I1|_SPL_B|1|MID_SHUNT  2.7439617672
LI1|_SPL_B|1|RB I1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|2|1 I1|_SPL_B|D2 I1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|2|P I1|_SPL_B|2|MID_SERIES 0  2e-13
RI1|_SPL_B|2|B I1|_SPL_B|D2 I1|_SPL_B|2|MID_SHUNT  2.7439617672
LI1|_SPL_B|2|RB I1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|A|1 I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|A|P I1|_SPL_B|A|MID_SERIES 0  2e-13
RI1|_SPL_B|A|B I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SHUNT  2.7439617672
LI1|_SPL_B|A|RB I1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|B|1 I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|B|P I1|_SPL_B|B|MID_SERIES 0  2e-13
RI1|_SPL_B|B|B I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SHUNT  2.7439617672
LI1|_SPL_B|B|RB I1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_A|I_1|B I1|_DFF_A|A1 I1|_DFF_A|I_1|MID  2e-12
II1|_DFF_A|I_1|B 0 I1|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_3|B I1|_DFF_A|A3 I1|_DFF_A|I_3|MID  2e-12
II1|_DFF_A|I_3|B 0 I1|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_A|I_T|B I1|_DFF_A|T1 I1|_DFF_A|I_T|MID  2e-12
II1|_DFF_A|I_T|B 0 I1|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_6|B I1|_DFF_A|Q1 I1|_DFF_A|I_6|MID  2e-12
II1|_DFF_A|I_6|B 0 I1|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_A|1|1 I1|_DFF_A|A1 I1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|1|P I1|_DFF_A|1|MID_SERIES 0  2e-13
RI1|_DFF_A|1|B I1|_DFF_A|A1 I1|_DFF_A|1|MID_SHUNT  2.7439617672
LI1|_DFF_A|1|RB I1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|23|1 I1|_DFF_A|A2 I1|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|23|B I1|_DFF_A|A2 I1|_DFF_A|23|MID_SHUNT  3.84154647408
LI1|_DFF_A|23|RB I1|_DFF_A|23|MID_SHUNT I1|_DFF_A|A3  2.1704737578552e-12
BI1|_DFF_A|3|1 I1|_DFF_A|A3 I1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|3|P I1|_DFF_A|3|MID_SERIES 0  2e-13
RI1|_DFF_A|3|B I1|_DFF_A|A3 I1|_DFF_A|3|MID_SHUNT  2.7439617672
LI1|_DFF_A|3|RB I1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|4|1 I1|_DFF_A|A4 I1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|4|P I1|_DFF_A|4|MID_SERIES 0  2e-13
RI1|_DFF_A|4|B I1|_DFF_A|A4 I1|_DFF_A|4|MID_SHUNT  2.7439617672
LI1|_DFF_A|4|RB I1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|T|1 I1|_DFF_A|T1 I1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|T|P I1|_DFF_A|T|MID_SERIES 0  2e-13
RI1|_DFF_A|T|B I1|_DFF_A|T1 I1|_DFF_A|T|MID_SHUNT  2.7439617672
LI1|_DFF_A|T|RB I1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|45|1 I1|_DFF_A|T2 I1|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|45|B I1|_DFF_A|T2 I1|_DFF_A|45|MID_SHUNT  3.84154647408
LI1|_DFF_A|45|RB I1|_DFF_A|45|MID_SHUNT I1|_DFF_A|A4  2.1704737578552e-12
BI1|_DFF_A|6|1 I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|6|P I1|_DFF_A|6|MID_SERIES 0  2e-13
RI1|_DFF_A|6|B I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SHUNT  2.7439617672
LI1|_DFF_A|6|RB I1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_B|I_1|B I1|_DFF_B|A1 I1|_DFF_B|I_1|MID  2e-12
II1|_DFF_B|I_1|B 0 I1|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_3|B I1|_DFF_B|A3 I1|_DFF_B|I_3|MID  2e-12
II1|_DFF_B|I_3|B 0 I1|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_B|I_T|B I1|_DFF_B|T1 I1|_DFF_B|I_T|MID  2e-12
II1|_DFF_B|I_T|B 0 I1|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_6|B I1|_DFF_B|Q1 I1|_DFF_B|I_6|MID  2e-12
II1|_DFF_B|I_6|B 0 I1|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_B|1|1 I1|_DFF_B|A1 I1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|1|P I1|_DFF_B|1|MID_SERIES 0  2e-13
RI1|_DFF_B|1|B I1|_DFF_B|A1 I1|_DFF_B|1|MID_SHUNT  2.7439617672
LI1|_DFF_B|1|RB I1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|23|1 I1|_DFF_B|A2 I1|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|23|B I1|_DFF_B|A2 I1|_DFF_B|23|MID_SHUNT  3.84154647408
LI1|_DFF_B|23|RB I1|_DFF_B|23|MID_SHUNT I1|_DFF_B|A3  2.1704737578552e-12
BI1|_DFF_B|3|1 I1|_DFF_B|A3 I1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|3|P I1|_DFF_B|3|MID_SERIES 0  2e-13
RI1|_DFF_B|3|B I1|_DFF_B|A3 I1|_DFF_B|3|MID_SHUNT  2.7439617672
LI1|_DFF_B|3|RB I1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|4|1 I1|_DFF_B|A4 I1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|4|P I1|_DFF_B|4|MID_SERIES 0  2e-13
RI1|_DFF_B|4|B I1|_DFF_B|A4 I1|_DFF_B|4|MID_SHUNT  2.7439617672
LI1|_DFF_B|4|RB I1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|T|1 I1|_DFF_B|T1 I1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|T|P I1|_DFF_B|T|MID_SERIES 0  2e-13
RI1|_DFF_B|T|B I1|_DFF_B|T1 I1|_DFF_B|T|MID_SHUNT  2.7439617672
LI1|_DFF_B|T|RB I1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|45|1 I1|_DFF_B|T2 I1|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|45|B I1|_DFF_B|T2 I1|_DFF_B|45|MID_SHUNT  3.84154647408
LI1|_DFF_B|45|RB I1|_DFF_B|45|MID_SHUNT I1|_DFF_B|A4  2.1704737578552e-12
BI1|_DFF_B|6|1 I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|6|P I1|_DFF_B|6|MID_SERIES 0  2e-13
RI1|_DFF_B|6|B I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SHUNT  2.7439617672
LI1|_DFF_B|6|RB I1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI1|_XOR|I_A1|B I1|_XOR|A1 I1|_XOR|I_A1|MID  2e-12
II1|_XOR|I_A1|B 0 I1|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_A3|B I1|_XOR|A3 I1|_XOR|I_A3|MID  2e-12
II1|_XOR|I_A3|B 0 I1|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B1|B I1|_XOR|B1 I1|_XOR|I_B1|MID  2e-12
II1|_XOR|I_B1|B 0 I1|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B3|B I1|_XOR|B3 I1|_XOR|I_B3|MID  2e-12
II1|_XOR|I_B3|B 0 I1|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_Q1|B I1|_XOR|Q1 I1|_XOR|I_Q1|MID  2e-12
II1|_XOR|I_Q1|B 0 I1|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_XOR|A1|1 I1|_XOR|A1 I1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A1|P I1|_XOR|A1|MID_SERIES 0  5e-13
RI1|_XOR|A1|B I1|_XOR|A1 I1|_XOR|A1|MID_SHUNT  2.7439617672
LI1|_XOR|A1|RB I1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A2|1 I1|_XOR|A2 I1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A2|P I1|_XOR|A2|MID_SERIES 0  5e-13
RI1|_XOR|A2|B I1|_XOR|A2 I1|_XOR|A2|MID_SHUNT  2.7439617672
LI1|_XOR|A2|RB I1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A3|1 I1|_XOR|A2 I1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A3|P I1|_XOR|A3|MID_SERIES I1|_XOR|A3  1.2e-12
RI1|_XOR|A3|B I1|_XOR|A2 I1|_XOR|A3|MID_SHUNT  2.7439617672
LI1|_XOR|A3|RB I1|_XOR|A3|MID_SHUNT I1|_XOR|A3  2.050338398468e-12
BI1|_XOR|B1|1 I1|_XOR|B1 I1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B1|P I1|_XOR|B1|MID_SERIES 0  5e-13
RI1|_XOR|B1|B I1|_XOR|B1 I1|_XOR|B1|MID_SHUNT  2.7439617672
LI1|_XOR|B1|RB I1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B2|1 I1|_XOR|B2 I1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B2|P I1|_XOR|B2|MID_SERIES 0  5e-13
RI1|_XOR|B2|B I1|_XOR|B2 I1|_XOR|B2|MID_SHUNT  2.7439617672
LI1|_XOR|B2|RB I1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B3|1 I1|_XOR|B2 I1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B3|P I1|_XOR|B3|MID_SERIES I1|_XOR|B3  1.2e-12
RI1|_XOR|B3|B I1|_XOR|B2 I1|_XOR|B3|MID_SHUNT  2.7439617672
LI1|_XOR|B3|RB I1|_XOR|B3|MID_SHUNT I1|_XOR|B3  2.050338398468e-12
BI1|_XOR|T1|1 I1|_XOR|T1 I1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|T1|P I1|_XOR|T1|MID_SERIES 0  5e-13
RI1|_XOR|T1|B I1|_XOR|T1 I1|_XOR|T1|MID_SHUNT  2.7439617672
LI1|_XOR|T1|RB I1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|T2|1 I1|_XOR|T2 I1|_XOR|ABTQ JJMIT AREA=2.0
RI1|_XOR|T2|B I1|_XOR|T2 I1|_XOR|T2|MID_SHUNT  3.429952209
LI1|_XOR|T2|RB I1|_XOR|T2|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|AB|1 I1|_XOR|AB I1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI1|_XOR|AB|P I1|_XOR|AB|MID_SERIES I1|_XOR|ABTQ  1.2e-12
RI1|_XOR|AB|B I1|_XOR|AB I1|_XOR|AB|MID_SHUNT  3.429952209
LI1|_XOR|AB|RB I1|_XOR|AB|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|ABTQ|1 I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|ABTQ|P I1|_XOR|ABTQ|MID_SERIES 0  5e-13
RI1|_XOR|ABTQ|B I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI1|_XOR|ABTQ|RB I1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|Q1|1 I1|_XOR|Q1 I1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|Q1|P I1|_XOR|Q1|MID_SERIES 0  5e-13
RI1|_XOR|Q1|B I1|_XOR|Q1 I1|_XOR|Q1|MID_SHUNT  2.7439617672
LI1|_XOR|Q1|RB I1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI1|_AND|I_A1|B I1|_AND|A1 I1|_AND|I_A1|MID  2e-12
II1|_AND|I_A1|B 0 I1|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_B1|B I1|_AND|B1 I1|_AND|I_B1|MID  2e-12
II1|_AND|I_B1|B 0 I1|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q3|B I1|_AND|Q3 I1|_AND|I_Q3|MID  2e-12
II1|_AND|I_Q3|B 0 I1|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1|_AND|I_Q2|B I1|_AND|Q2 I1|_AND|I_Q2|MID  2e-12
II1|_AND|I_Q2|B 0 I1|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q1|B I1|_AND|Q1 I1|_AND|I_Q1|MID  2e-12
II1|_AND|I_Q1|B 0 I1|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_AND|A1|1 I1|_AND|A1 I1|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A1|P I1|_AND|A1|MID_SERIES 0  2e-13
RI1|_AND|A1|B I1|_AND|A1 I1|_AND|A1|MID_SHUNT  2.7439617672
LI1|_AND|A1|RB I1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A2|1 I1|_AND|A2 I1|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A2|P I1|_AND|A2|MID_SERIES 0  2e-13
RI1|_AND|A2|B I1|_AND|A2 I1|_AND|A2|MID_SHUNT  2.7439617672
LI1|_AND|A2|RB I1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A12|1 I1|_AND|A2 I1|_AND|A3 JJMIT AREA=1.7857142857142858
RI1|_AND|A12|B I1|_AND|A2 I1|_AND|A12|MID_SHUNT  3.84154647408
LI1|_AND|A12|RB I1|_AND|A12|MID_SHUNT I1|_AND|A3  2.1704737578552e-12
BI1|_AND|B1|1 I1|_AND|B1 I1|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B1|P I1|_AND|B1|MID_SERIES 0  2e-13
RI1|_AND|B1|B I1|_AND|B1 I1|_AND|B1|MID_SHUNT  2.7439617672
LI1|_AND|B1|RB I1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B2|1 I1|_AND|B2 I1|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B2|P I1|_AND|B2|MID_SERIES 0  2e-13
RI1|_AND|B2|B I1|_AND|B2 I1|_AND|B2|MID_SHUNT  2.7439617672
LI1|_AND|B2|RB I1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B12|1 I1|_AND|B2 I1|_AND|B3 JJMIT AREA=1.7857142857142858
RI1|_AND|B12|B I1|_AND|B2 I1|_AND|B12|MID_SHUNT  3.84154647408
LI1|_AND|B12|RB I1|_AND|B12|MID_SHUNT I1|_AND|B3  2.1704737578552e-12
BI1|_AND|Q2|1 I1|_AND|Q2 I1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q2|P I1|_AND|Q2|MID_SERIES 0  2e-13
RI1|_AND|Q2|B I1|_AND|Q2 I1|_AND|Q2|MID_SHUNT  2.7439617672
LI1|_AND|Q2|RB I1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|Q1|1 I1|_AND|Q1 I1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q1|P I1|_AND|Q1|MID_SERIES 0  2e-13
RI1|_AND|Q1|B I1|_AND|Q1 I1|_AND|Q1|MID_SHUNT  2.7439617672
LI1|_AND|Q1|RB I1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_A|I_D1|B I2|_SPL_A|D1 I2|_SPL_A|I_D1|MID  2e-12
II2|_SPL_A|I_D1|B 0 I2|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_D2|B I2|_SPL_A|D2 I2|_SPL_A|I_D2|MID  2e-12
II2|_SPL_A|I_D2|B 0 I2|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_A|I_Q1|B I2|_SPL_A|QA1 I2|_SPL_A|I_Q1|MID  2e-12
II2|_SPL_A|I_Q1|B 0 I2|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_Q2|B I2|_SPL_A|QB1 I2|_SPL_A|I_Q2|MID  2e-12
II2|_SPL_A|I_Q2|B 0 I2|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_A|1|1 I2|_SPL_A|D1 I2|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|1|P I2|_SPL_A|1|MID_SERIES 0  2e-13
RI2|_SPL_A|1|B I2|_SPL_A|D1 I2|_SPL_A|1|MID_SHUNT  2.7439617672
LI2|_SPL_A|1|RB I2|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|2|1 I2|_SPL_A|D2 I2|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|2|P I2|_SPL_A|2|MID_SERIES 0  2e-13
RI2|_SPL_A|2|B I2|_SPL_A|D2 I2|_SPL_A|2|MID_SHUNT  2.7439617672
LI2|_SPL_A|2|RB I2|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|A|1 I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|A|P I2|_SPL_A|A|MID_SERIES 0  2e-13
RI2|_SPL_A|A|B I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SHUNT  2.7439617672
LI2|_SPL_A|A|RB I2|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|B|1 I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|B|P I2|_SPL_A|B|MID_SERIES 0  2e-13
RI2|_SPL_A|B|B I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SHUNT  2.7439617672
LI2|_SPL_A|B|RB I2|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_B|I_D1|B I2|_SPL_B|D1 I2|_SPL_B|I_D1|MID  2e-12
II2|_SPL_B|I_D1|B 0 I2|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_D2|B I2|_SPL_B|D2 I2|_SPL_B|I_D2|MID  2e-12
II2|_SPL_B|I_D2|B 0 I2|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_B|I_Q1|B I2|_SPL_B|QA1 I2|_SPL_B|I_Q1|MID  2e-12
II2|_SPL_B|I_Q1|B 0 I2|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_Q2|B I2|_SPL_B|QB1 I2|_SPL_B|I_Q2|MID  2e-12
II2|_SPL_B|I_Q2|B 0 I2|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_B|1|1 I2|_SPL_B|D1 I2|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|1|P I2|_SPL_B|1|MID_SERIES 0  2e-13
RI2|_SPL_B|1|B I2|_SPL_B|D1 I2|_SPL_B|1|MID_SHUNT  2.7439617672
LI2|_SPL_B|1|RB I2|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|2|1 I2|_SPL_B|D2 I2|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|2|P I2|_SPL_B|2|MID_SERIES 0  2e-13
RI2|_SPL_B|2|B I2|_SPL_B|D2 I2|_SPL_B|2|MID_SHUNT  2.7439617672
LI2|_SPL_B|2|RB I2|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|A|1 I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|A|P I2|_SPL_B|A|MID_SERIES 0  2e-13
RI2|_SPL_B|A|B I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SHUNT  2.7439617672
LI2|_SPL_B|A|RB I2|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|B|1 I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|B|P I2|_SPL_B|B|MID_SERIES 0  2e-13
RI2|_SPL_B|B|B I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SHUNT  2.7439617672
LI2|_SPL_B|B|RB I2|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_A|I_1|B I2|_DFF_A|A1 I2|_DFF_A|I_1|MID  2e-12
II2|_DFF_A|I_1|B 0 I2|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_3|B I2|_DFF_A|A3 I2|_DFF_A|I_3|MID  2e-12
II2|_DFF_A|I_3|B 0 I2|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_A|I_T|B I2|_DFF_A|T1 I2|_DFF_A|I_T|MID  2e-12
II2|_DFF_A|I_T|B 0 I2|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_6|B I2|_DFF_A|Q1 I2|_DFF_A|I_6|MID  2e-12
II2|_DFF_A|I_6|B 0 I2|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_A|1|1 I2|_DFF_A|A1 I2|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|1|P I2|_DFF_A|1|MID_SERIES 0  2e-13
RI2|_DFF_A|1|B I2|_DFF_A|A1 I2|_DFF_A|1|MID_SHUNT  2.7439617672
LI2|_DFF_A|1|RB I2|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|23|1 I2|_DFF_A|A2 I2|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|23|B I2|_DFF_A|A2 I2|_DFF_A|23|MID_SHUNT  3.84154647408
LI2|_DFF_A|23|RB I2|_DFF_A|23|MID_SHUNT I2|_DFF_A|A3  2.1704737578552e-12
BI2|_DFF_A|3|1 I2|_DFF_A|A3 I2|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|3|P I2|_DFF_A|3|MID_SERIES 0  2e-13
RI2|_DFF_A|3|B I2|_DFF_A|A3 I2|_DFF_A|3|MID_SHUNT  2.7439617672
LI2|_DFF_A|3|RB I2|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|4|1 I2|_DFF_A|A4 I2|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|4|P I2|_DFF_A|4|MID_SERIES 0  2e-13
RI2|_DFF_A|4|B I2|_DFF_A|A4 I2|_DFF_A|4|MID_SHUNT  2.7439617672
LI2|_DFF_A|4|RB I2|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|T|1 I2|_DFF_A|T1 I2|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|T|P I2|_DFF_A|T|MID_SERIES 0  2e-13
RI2|_DFF_A|T|B I2|_DFF_A|T1 I2|_DFF_A|T|MID_SHUNT  2.7439617672
LI2|_DFF_A|T|RB I2|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|45|1 I2|_DFF_A|T2 I2|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|45|B I2|_DFF_A|T2 I2|_DFF_A|45|MID_SHUNT  3.84154647408
LI2|_DFF_A|45|RB I2|_DFF_A|45|MID_SHUNT I2|_DFF_A|A4  2.1704737578552e-12
BI2|_DFF_A|6|1 I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|6|P I2|_DFF_A|6|MID_SERIES 0  2e-13
RI2|_DFF_A|6|B I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SHUNT  2.7439617672
LI2|_DFF_A|6|RB I2|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_B|I_1|B I2|_DFF_B|A1 I2|_DFF_B|I_1|MID  2e-12
II2|_DFF_B|I_1|B 0 I2|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_3|B I2|_DFF_B|A3 I2|_DFF_B|I_3|MID  2e-12
II2|_DFF_B|I_3|B 0 I2|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_B|I_T|B I2|_DFF_B|T1 I2|_DFF_B|I_T|MID  2e-12
II2|_DFF_B|I_T|B 0 I2|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_6|B I2|_DFF_B|Q1 I2|_DFF_B|I_6|MID  2e-12
II2|_DFF_B|I_6|B 0 I2|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_B|1|1 I2|_DFF_B|A1 I2|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|1|P I2|_DFF_B|1|MID_SERIES 0  2e-13
RI2|_DFF_B|1|B I2|_DFF_B|A1 I2|_DFF_B|1|MID_SHUNT  2.7439617672
LI2|_DFF_B|1|RB I2|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|23|1 I2|_DFF_B|A2 I2|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|23|B I2|_DFF_B|A2 I2|_DFF_B|23|MID_SHUNT  3.84154647408
LI2|_DFF_B|23|RB I2|_DFF_B|23|MID_SHUNT I2|_DFF_B|A3  2.1704737578552e-12
BI2|_DFF_B|3|1 I2|_DFF_B|A3 I2|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|3|P I2|_DFF_B|3|MID_SERIES 0  2e-13
RI2|_DFF_B|3|B I2|_DFF_B|A3 I2|_DFF_B|3|MID_SHUNT  2.7439617672
LI2|_DFF_B|3|RB I2|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|4|1 I2|_DFF_B|A4 I2|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|4|P I2|_DFF_B|4|MID_SERIES 0  2e-13
RI2|_DFF_B|4|B I2|_DFF_B|A4 I2|_DFF_B|4|MID_SHUNT  2.7439617672
LI2|_DFF_B|4|RB I2|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|T|1 I2|_DFF_B|T1 I2|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|T|P I2|_DFF_B|T|MID_SERIES 0  2e-13
RI2|_DFF_B|T|B I2|_DFF_B|T1 I2|_DFF_B|T|MID_SHUNT  2.7439617672
LI2|_DFF_B|T|RB I2|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|45|1 I2|_DFF_B|T2 I2|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|45|B I2|_DFF_B|T2 I2|_DFF_B|45|MID_SHUNT  3.84154647408
LI2|_DFF_B|45|RB I2|_DFF_B|45|MID_SHUNT I2|_DFF_B|A4  2.1704737578552e-12
BI2|_DFF_B|6|1 I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|6|P I2|_DFF_B|6|MID_SERIES 0  2e-13
RI2|_DFF_B|6|B I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SHUNT  2.7439617672
LI2|_DFF_B|6|RB I2|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI2|_XOR|I_A1|B I2|_XOR|A1 I2|_XOR|I_A1|MID  2e-12
II2|_XOR|I_A1|B 0 I2|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_A3|B I2|_XOR|A3 I2|_XOR|I_A3|MID  2e-12
II2|_XOR|I_A3|B 0 I2|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B1|B I2|_XOR|B1 I2|_XOR|I_B1|MID  2e-12
II2|_XOR|I_B1|B 0 I2|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B3|B I2|_XOR|B3 I2|_XOR|I_B3|MID  2e-12
II2|_XOR|I_B3|B 0 I2|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_Q1|B I2|_XOR|Q1 I2|_XOR|I_Q1|MID  2e-12
II2|_XOR|I_Q1|B 0 I2|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_XOR|A1|1 I2|_XOR|A1 I2|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A1|P I2|_XOR|A1|MID_SERIES 0  5e-13
RI2|_XOR|A1|B I2|_XOR|A1 I2|_XOR|A1|MID_SHUNT  2.7439617672
LI2|_XOR|A1|RB I2|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A2|1 I2|_XOR|A2 I2|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A2|P I2|_XOR|A2|MID_SERIES 0  5e-13
RI2|_XOR|A2|B I2|_XOR|A2 I2|_XOR|A2|MID_SHUNT  2.7439617672
LI2|_XOR|A2|RB I2|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A3|1 I2|_XOR|A2 I2|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A3|P I2|_XOR|A3|MID_SERIES I2|_XOR|A3  1.2e-12
RI2|_XOR|A3|B I2|_XOR|A2 I2|_XOR|A3|MID_SHUNT  2.7439617672
LI2|_XOR|A3|RB I2|_XOR|A3|MID_SHUNT I2|_XOR|A3  2.050338398468e-12
BI2|_XOR|B1|1 I2|_XOR|B1 I2|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B1|P I2|_XOR|B1|MID_SERIES 0  5e-13
RI2|_XOR|B1|B I2|_XOR|B1 I2|_XOR|B1|MID_SHUNT  2.7439617672
LI2|_XOR|B1|RB I2|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B2|1 I2|_XOR|B2 I2|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B2|P I2|_XOR|B2|MID_SERIES 0  5e-13
RI2|_XOR|B2|B I2|_XOR|B2 I2|_XOR|B2|MID_SHUNT  2.7439617672
LI2|_XOR|B2|RB I2|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B3|1 I2|_XOR|B2 I2|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B3|P I2|_XOR|B3|MID_SERIES I2|_XOR|B3  1.2e-12
RI2|_XOR|B3|B I2|_XOR|B2 I2|_XOR|B3|MID_SHUNT  2.7439617672
LI2|_XOR|B3|RB I2|_XOR|B3|MID_SHUNT I2|_XOR|B3  2.050338398468e-12
BI2|_XOR|T1|1 I2|_XOR|T1 I2|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|T1|P I2|_XOR|T1|MID_SERIES 0  5e-13
RI2|_XOR|T1|B I2|_XOR|T1 I2|_XOR|T1|MID_SHUNT  2.7439617672
LI2|_XOR|T1|RB I2|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|T2|1 I2|_XOR|T2 I2|_XOR|ABTQ JJMIT AREA=2.0
RI2|_XOR|T2|B I2|_XOR|T2 I2|_XOR|T2|MID_SHUNT  3.429952209
LI2|_XOR|T2|RB I2|_XOR|T2|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|AB|1 I2|_XOR|AB I2|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI2|_XOR|AB|P I2|_XOR|AB|MID_SERIES I2|_XOR|ABTQ  1.2e-12
RI2|_XOR|AB|B I2|_XOR|AB I2|_XOR|AB|MID_SHUNT  3.429952209
LI2|_XOR|AB|RB I2|_XOR|AB|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|ABTQ|1 I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|ABTQ|P I2|_XOR|ABTQ|MID_SERIES 0  5e-13
RI2|_XOR|ABTQ|B I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI2|_XOR|ABTQ|RB I2|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|Q1|1 I2|_XOR|Q1 I2|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|Q1|P I2|_XOR|Q1|MID_SERIES 0  5e-13
RI2|_XOR|Q1|B I2|_XOR|Q1 I2|_XOR|Q1|MID_SHUNT  2.7439617672
LI2|_XOR|Q1|RB I2|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI2|_AND|I_A1|B I2|_AND|A1 I2|_AND|I_A1|MID  2e-12
II2|_AND|I_A1|B 0 I2|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_B1|B I2|_AND|B1 I2|_AND|I_B1|MID  2e-12
II2|_AND|I_B1|B 0 I2|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q3|B I2|_AND|Q3 I2|_AND|I_Q3|MID  2e-12
II2|_AND|I_Q3|B 0 I2|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2|_AND|I_Q2|B I2|_AND|Q2 I2|_AND|I_Q2|MID  2e-12
II2|_AND|I_Q2|B 0 I2|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q1|B I2|_AND|Q1 I2|_AND|I_Q1|MID  2e-12
II2|_AND|I_Q1|B 0 I2|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_AND|A1|1 I2|_AND|A1 I2|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A1|P I2|_AND|A1|MID_SERIES 0  2e-13
RI2|_AND|A1|B I2|_AND|A1 I2|_AND|A1|MID_SHUNT  2.7439617672
LI2|_AND|A1|RB I2|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A2|1 I2|_AND|A2 I2|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A2|P I2|_AND|A2|MID_SERIES 0  2e-13
RI2|_AND|A2|B I2|_AND|A2 I2|_AND|A2|MID_SHUNT  2.7439617672
LI2|_AND|A2|RB I2|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A12|1 I2|_AND|A2 I2|_AND|A3 JJMIT AREA=1.7857142857142858
RI2|_AND|A12|B I2|_AND|A2 I2|_AND|A12|MID_SHUNT  3.84154647408
LI2|_AND|A12|RB I2|_AND|A12|MID_SHUNT I2|_AND|A3  2.1704737578552e-12
BI2|_AND|B1|1 I2|_AND|B1 I2|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B1|P I2|_AND|B1|MID_SERIES 0  2e-13
RI2|_AND|B1|B I2|_AND|B1 I2|_AND|B1|MID_SHUNT  2.7439617672
LI2|_AND|B1|RB I2|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B2|1 I2|_AND|B2 I2|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B2|P I2|_AND|B2|MID_SERIES 0  2e-13
RI2|_AND|B2|B I2|_AND|B2 I2|_AND|B2|MID_SHUNT  2.7439617672
LI2|_AND|B2|RB I2|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B12|1 I2|_AND|B2 I2|_AND|B3 JJMIT AREA=1.7857142857142858
RI2|_AND|B12|B I2|_AND|B2 I2|_AND|B12|MID_SHUNT  3.84154647408
LI2|_AND|B12|RB I2|_AND|B12|MID_SHUNT I2|_AND|B3  2.1704737578552e-12
BI2|_AND|Q2|1 I2|_AND|Q2 I2|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q2|P I2|_AND|Q2|MID_SERIES 0  2e-13
RI2|_AND|Q2|B I2|_AND|Q2 I2|_AND|Q2|MID_SHUNT  2.7439617672
LI2|_AND|Q2|RB I2|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|Q1|1 I2|_AND|Q1 I2|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q1|P I2|_AND|Q1|MID_SERIES 0  2e-13
RI2|_AND|Q1|B I2|_AND|Q1 I2|_AND|Q1|MID_SHUNT  2.7439617672
LI2|_AND|Q1|RB I2|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_A|I_D1|B I3|_SPL_A|D1 I3|_SPL_A|I_D1|MID  2e-12
II3|_SPL_A|I_D1|B 0 I3|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_D2|B I3|_SPL_A|D2 I3|_SPL_A|I_D2|MID  2e-12
II3|_SPL_A|I_D2|B 0 I3|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_A|I_Q1|B I3|_SPL_A|QA1 I3|_SPL_A|I_Q1|MID  2e-12
II3|_SPL_A|I_Q1|B 0 I3|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_Q2|B I3|_SPL_A|QB1 I3|_SPL_A|I_Q2|MID  2e-12
II3|_SPL_A|I_Q2|B 0 I3|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_A|1|1 I3|_SPL_A|D1 I3|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|1|P I3|_SPL_A|1|MID_SERIES 0  2e-13
RI3|_SPL_A|1|B I3|_SPL_A|D1 I3|_SPL_A|1|MID_SHUNT  2.7439617672
LI3|_SPL_A|1|RB I3|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|2|1 I3|_SPL_A|D2 I3|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|2|P I3|_SPL_A|2|MID_SERIES 0  2e-13
RI3|_SPL_A|2|B I3|_SPL_A|D2 I3|_SPL_A|2|MID_SHUNT  2.7439617672
LI3|_SPL_A|2|RB I3|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|A|1 I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|A|P I3|_SPL_A|A|MID_SERIES 0  2e-13
RI3|_SPL_A|A|B I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SHUNT  2.7439617672
LI3|_SPL_A|A|RB I3|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|B|1 I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|B|P I3|_SPL_A|B|MID_SERIES 0  2e-13
RI3|_SPL_A|B|B I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SHUNT  2.7439617672
LI3|_SPL_A|B|RB I3|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_B|I_D1|B I3|_SPL_B|D1 I3|_SPL_B|I_D1|MID  2e-12
II3|_SPL_B|I_D1|B 0 I3|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_D2|B I3|_SPL_B|D2 I3|_SPL_B|I_D2|MID  2e-12
II3|_SPL_B|I_D2|B 0 I3|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_B|I_Q1|B I3|_SPL_B|QA1 I3|_SPL_B|I_Q1|MID  2e-12
II3|_SPL_B|I_Q1|B 0 I3|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_Q2|B I3|_SPL_B|QB1 I3|_SPL_B|I_Q2|MID  2e-12
II3|_SPL_B|I_Q2|B 0 I3|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_B|1|1 I3|_SPL_B|D1 I3|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|1|P I3|_SPL_B|1|MID_SERIES 0  2e-13
RI3|_SPL_B|1|B I3|_SPL_B|D1 I3|_SPL_B|1|MID_SHUNT  2.7439617672
LI3|_SPL_B|1|RB I3|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|2|1 I3|_SPL_B|D2 I3|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|2|P I3|_SPL_B|2|MID_SERIES 0  2e-13
RI3|_SPL_B|2|B I3|_SPL_B|D2 I3|_SPL_B|2|MID_SHUNT  2.7439617672
LI3|_SPL_B|2|RB I3|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|A|1 I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|A|P I3|_SPL_B|A|MID_SERIES 0  2e-13
RI3|_SPL_B|A|B I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SHUNT  2.7439617672
LI3|_SPL_B|A|RB I3|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|B|1 I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|B|P I3|_SPL_B|B|MID_SERIES 0  2e-13
RI3|_SPL_B|B|B I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SHUNT  2.7439617672
LI3|_SPL_B|B|RB I3|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_A|I_1|B I3|_DFF_A|A1 I3|_DFF_A|I_1|MID  2e-12
II3|_DFF_A|I_1|B 0 I3|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_3|B I3|_DFF_A|A3 I3|_DFF_A|I_3|MID  2e-12
II3|_DFF_A|I_3|B 0 I3|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_A|I_T|B I3|_DFF_A|T1 I3|_DFF_A|I_T|MID  2e-12
II3|_DFF_A|I_T|B 0 I3|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_6|B I3|_DFF_A|Q1 I3|_DFF_A|I_6|MID  2e-12
II3|_DFF_A|I_6|B 0 I3|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_A|1|1 I3|_DFF_A|A1 I3|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|1|P I3|_DFF_A|1|MID_SERIES 0  2e-13
RI3|_DFF_A|1|B I3|_DFF_A|A1 I3|_DFF_A|1|MID_SHUNT  2.7439617672
LI3|_DFF_A|1|RB I3|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|23|1 I3|_DFF_A|A2 I3|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|23|B I3|_DFF_A|A2 I3|_DFF_A|23|MID_SHUNT  3.84154647408
LI3|_DFF_A|23|RB I3|_DFF_A|23|MID_SHUNT I3|_DFF_A|A3  2.1704737578552e-12
BI3|_DFF_A|3|1 I3|_DFF_A|A3 I3|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|3|P I3|_DFF_A|3|MID_SERIES 0  2e-13
RI3|_DFF_A|3|B I3|_DFF_A|A3 I3|_DFF_A|3|MID_SHUNT  2.7439617672
LI3|_DFF_A|3|RB I3|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|4|1 I3|_DFF_A|A4 I3|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|4|P I3|_DFF_A|4|MID_SERIES 0  2e-13
RI3|_DFF_A|4|B I3|_DFF_A|A4 I3|_DFF_A|4|MID_SHUNT  2.7439617672
LI3|_DFF_A|4|RB I3|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|T|1 I3|_DFF_A|T1 I3|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|T|P I3|_DFF_A|T|MID_SERIES 0  2e-13
RI3|_DFF_A|T|B I3|_DFF_A|T1 I3|_DFF_A|T|MID_SHUNT  2.7439617672
LI3|_DFF_A|T|RB I3|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|45|1 I3|_DFF_A|T2 I3|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|45|B I3|_DFF_A|T2 I3|_DFF_A|45|MID_SHUNT  3.84154647408
LI3|_DFF_A|45|RB I3|_DFF_A|45|MID_SHUNT I3|_DFF_A|A4  2.1704737578552e-12
BI3|_DFF_A|6|1 I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|6|P I3|_DFF_A|6|MID_SERIES 0  2e-13
RI3|_DFF_A|6|B I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SHUNT  2.7439617672
LI3|_DFF_A|6|RB I3|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_B|I_1|B I3|_DFF_B|A1 I3|_DFF_B|I_1|MID  2e-12
II3|_DFF_B|I_1|B 0 I3|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_3|B I3|_DFF_B|A3 I3|_DFF_B|I_3|MID  2e-12
II3|_DFF_B|I_3|B 0 I3|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_B|I_T|B I3|_DFF_B|T1 I3|_DFF_B|I_T|MID  2e-12
II3|_DFF_B|I_T|B 0 I3|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_6|B I3|_DFF_B|Q1 I3|_DFF_B|I_6|MID  2e-12
II3|_DFF_B|I_6|B 0 I3|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_B|1|1 I3|_DFF_B|A1 I3|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|1|P I3|_DFF_B|1|MID_SERIES 0  2e-13
RI3|_DFF_B|1|B I3|_DFF_B|A1 I3|_DFF_B|1|MID_SHUNT  2.7439617672
LI3|_DFF_B|1|RB I3|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|23|1 I3|_DFF_B|A2 I3|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|23|B I3|_DFF_B|A2 I3|_DFF_B|23|MID_SHUNT  3.84154647408
LI3|_DFF_B|23|RB I3|_DFF_B|23|MID_SHUNT I3|_DFF_B|A3  2.1704737578552e-12
BI3|_DFF_B|3|1 I3|_DFF_B|A3 I3|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|3|P I3|_DFF_B|3|MID_SERIES 0  2e-13
RI3|_DFF_B|3|B I3|_DFF_B|A3 I3|_DFF_B|3|MID_SHUNT  2.7439617672
LI3|_DFF_B|3|RB I3|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|4|1 I3|_DFF_B|A4 I3|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|4|P I3|_DFF_B|4|MID_SERIES 0  2e-13
RI3|_DFF_B|4|B I3|_DFF_B|A4 I3|_DFF_B|4|MID_SHUNT  2.7439617672
LI3|_DFF_B|4|RB I3|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|T|1 I3|_DFF_B|T1 I3|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|T|P I3|_DFF_B|T|MID_SERIES 0  2e-13
RI3|_DFF_B|T|B I3|_DFF_B|T1 I3|_DFF_B|T|MID_SHUNT  2.7439617672
LI3|_DFF_B|T|RB I3|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|45|1 I3|_DFF_B|T2 I3|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|45|B I3|_DFF_B|T2 I3|_DFF_B|45|MID_SHUNT  3.84154647408
LI3|_DFF_B|45|RB I3|_DFF_B|45|MID_SHUNT I3|_DFF_B|A4  2.1704737578552e-12
BI3|_DFF_B|6|1 I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|6|P I3|_DFF_B|6|MID_SERIES 0  2e-13
RI3|_DFF_B|6|B I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SHUNT  2.7439617672
LI3|_DFF_B|6|RB I3|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI3|_XOR|I_A1|B I3|_XOR|A1 I3|_XOR|I_A1|MID  2e-12
II3|_XOR|I_A1|B 0 I3|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_A3|B I3|_XOR|A3 I3|_XOR|I_A3|MID  2e-12
II3|_XOR|I_A3|B 0 I3|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B1|B I3|_XOR|B1 I3|_XOR|I_B1|MID  2e-12
II3|_XOR|I_B1|B 0 I3|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B3|B I3|_XOR|B3 I3|_XOR|I_B3|MID  2e-12
II3|_XOR|I_B3|B 0 I3|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_Q1|B I3|_XOR|Q1 I3|_XOR|I_Q1|MID  2e-12
II3|_XOR|I_Q1|B 0 I3|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_XOR|A1|1 I3|_XOR|A1 I3|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A1|P I3|_XOR|A1|MID_SERIES 0  5e-13
RI3|_XOR|A1|B I3|_XOR|A1 I3|_XOR|A1|MID_SHUNT  2.7439617672
LI3|_XOR|A1|RB I3|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A2|1 I3|_XOR|A2 I3|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A2|P I3|_XOR|A2|MID_SERIES 0  5e-13
RI3|_XOR|A2|B I3|_XOR|A2 I3|_XOR|A2|MID_SHUNT  2.7439617672
LI3|_XOR|A2|RB I3|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A3|1 I3|_XOR|A2 I3|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A3|P I3|_XOR|A3|MID_SERIES I3|_XOR|A3  1.2e-12
RI3|_XOR|A3|B I3|_XOR|A2 I3|_XOR|A3|MID_SHUNT  2.7439617672
LI3|_XOR|A3|RB I3|_XOR|A3|MID_SHUNT I3|_XOR|A3  2.050338398468e-12
BI3|_XOR|B1|1 I3|_XOR|B1 I3|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B1|P I3|_XOR|B1|MID_SERIES 0  5e-13
RI3|_XOR|B1|B I3|_XOR|B1 I3|_XOR|B1|MID_SHUNT  2.7439617672
LI3|_XOR|B1|RB I3|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B2|1 I3|_XOR|B2 I3|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B2|P I3|_XOR|B2|MID_SERIES 0  5e-13
RI3|_XOR|B2|B I3|_XOR|B2 I3|_XOR|B2|MID_SHUNT  2.7439617672
LI3|_XOR|B2|RB I3|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B3|1 I3|_XOR|B2 I3|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B3|P I3|_XOR|B3|MID_SERIES I3|_XOR|B3  1.2e-12
RI3|_XOR|B3|B I3|_XOR|B2 I3|_XOR|B3|MID_SHUNT  2.7439617672
LI3|_XOR|B3|RB I3|_XOR|B3|MID_SHUNT I3|_XOR|B3  2.050338398468e-12
BI3|_XOR|T1|1 I3|_XOR|T1 I3|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|T1|P I3|_XOR|T1|MID_SERIES 0  5e-13
RI3|_XOR|T1|B I3|_XOR|T1 I3|_XOR|T1|MID_SHUNT  2.7439617672
LI3|_XOR|T1|RB I3|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|T2|1 I3|_XOR|T2 I3|_XOR|ABTQ JJMIT AREA=2.0
RI3|_XOR|T2|B I3|_XOR|T2 I3|_XOR|T2|MID_SHUNT  3.429952209
LI3|_XOR|T2|RB I3|_XOR|T2|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|AB|1 I3|_XOR|AB I3|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI3|_XOR|AB|P I3|_XOR|AB|MID_SERIES I3|_XOR|ABTQ  1.2e-12
RI3|_XOR|AB|B I3|_XOR|AB I3|_XOR|AB|MID_SHUNT  3.429952209
LI3|_XOR|AB|RB I3|_XOR|AB|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|ABTQ|1 I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|ABTQ|P I3|_XOR|ABTQ|MID_SERIES 0  5e-13
RI3|_XOR|ABTQ|B I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI3|_XOR|ABTQ|RB I3|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|Q1|1 I3|_XOR|Q1 I3|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|Q1|P I3|_XOR|Q1|MID_SERIES 0  5e-13
RI3|_XOR|Q1|B I3|_XOR|Q1 I3|_XOR|Q1|MID_SHUNT  2.7439617672
LI3|_XOR|Q1|RB I3|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI3|_AND|I_A1|B I3|_AND|A1 I3|_AND|I_A1|MID  2e-12
II3|_AND|I_A1|B 0 I3|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_B1|B I3|_AND|B1 I3|_AND|I_B1|MID  2e-12
II3|_AND|I_B1|B 0 I3|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q3|B I3|_AND|Q3 I3|_AND|I_Q3|MID  2e-12
II3|_AND|I_Q3|B 0 I3|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3|_AND|I_Q2|B I3|_AND|Q2 I3|_AND|I_Q2|MID  2e-12
II3|_AND|I_Q2|B 0 I3|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q1|B I3|_AND|Q1 I3|_AND|I_Q1|MID  2e-12
II3|_AND|I_Q1|B 0 I3|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_AND|A1|1 I3|_AND|A1 I3|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A1|P I3|_AND|A1|MID_SERIES 0  2e-13
RI3|_AND|A1|B I3|_AND|A1 I3|_AND|A1|MID_SHUNT  2.7439617672
LI3|_AND|A1|RB I3|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A2|1 I3|_AND|A2 I3|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A2|P I3|_AND|A2|MID_SERIES 0  2e-13
RI3|_AND|A2|B I3|_AND|A2 I3|_AND|A2|MID_SHUNT  2.7439617672
LI3|_AND|A2|RB I3|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A12|1 I3|_AND|A2 I3|_AND|A3 JJMIT AREA=1.7857142857142858
RI3|_AND|A12|B I3|_AND|A2 I3|_AND|A12|MID_SHUNT  3.84154647408
LI3|_AND|A12|RB I3|_AND|A12|MID_SHUNT I3|_AND|A3  2.1704737578552e-12
BI3|_AND|B1|1 I3|_AND|B1 I3|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B1|P I3|_AND|B1|MID_SERIES 0  2e-13
RI3|_AND|B1|B I3|_AND|B1 I3|_AND|B1|MID_SHUNT  2.7439617672
LI3|_AND|B1|RB I3|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B2|1 I3|_AND|B2 I3|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B2|P I3|_AND|B2|MID_SERIES 0  2e-13
RI3|_AND|B2|B I3|_AND|B2 I3|_AND|B2|MID_SHUNT  2.7439617672
LI3|_AND|B2|RB I3|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B12|1 I3|_AND|B2 I3|_AND|B3 JJMIT AREA=1.7857142857142858
RI3|_AND|B12|B I3|_AND|B2 I3|_AND|B12|MID_SHUNT  3.84154647408
LI3|_AND|B12|RB I3|_AND|B12|MID_SHUNT I3|_AND|B3  2.1704737578552e-12
BI3|_AND|Q2|1 I3|_AND|Q2 I3|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q2|P I3|_AND|Q2|MID_SERIES 0  2e-13
RI3|_AND|Q2|B I3|_AND|Q2 I3|_AND|Q2|MID_SHUNT  2.7439617672
LI3|_AND|Q2|RB I3|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|Q1|1 I3|_AND|Q1 I3|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q1|P I3|_AND|Q1|MID_SERIES 0  2e-13
RI3|_AND|Q1|B I3|_AND|Q1 I3|_AND|Q1|MID_SHUNT  2.7439617672
LI3|_AND|Q1|RB I3|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|I_D1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|I_D1|MID  2e-12
ISPL_IP2_0|SPL1|I_D1|B 0 SPL_IP2_0|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL1|I_D2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|I_D2|MID  2e-12
ISPL_IP2_0|SPL1|I_D2|B 0 SPL_IP2_0|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_IP2_0|SPL1|I_Q1|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|I_Q1|MID  2e-12
ISPL_IP2_0|SPL1|I_Q1|B 0 SPL_IP2_0|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL1|I_Q2|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|I_Q2|MID  2e-12
ISPL_IP2_0|SPL1|I_Q2|B 0 SPL_IP2_0|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_IP2_0|SPL1|1|1 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|1|P SPL_IP2_0|SPL1|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|1|RB SPL_IP2_0|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|2|1 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|2|P SPL_IP2_0|SPL1|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|2|RB SPL_IP2_0|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|A|1 SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|A|P SPL_IP2_0|SPL1|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|A|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|A|RB SPL_IP2_0|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|B|1 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|B|P SPL_IP2_0|SPL1|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|B|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|B|RB SPL_IP2_0|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL2|I_D1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|I_D1|MID  2e-12
ISPL_IP2_0|SPL2|I_D1|B 0 SPL_IP2_0|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL2|I_D2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|I_D2|MID  2e-12
ISPL_IP2_0|SPL2|I_D2|B 0 SPL_IP2_0|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_IP2_0|SPL2|I_Q1|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|I_Q1|MID  2e-12
ISPL_IP2_0|SPL2|I_Q1|B 0 SPL_IP2_0|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL2|I_Q2|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|I_Q2|MID  2e-12
ISPL_IP2_0|SPL2|I_Q2|B 0 SPL_IP2_0|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_IP2_0|SPL2|1|1 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|1|P SPL_IP2_0|SPL2|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|1|RB SPL_IP2_0|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|2|1 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|2|P SPL_IP2_0|SPL2|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|2|RB SPL_IP2_0|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|A|1 SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|A|P SPL_IP2_0|SPL2|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|A|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|A|RB SPL_IP2_0|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|B|1 SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|B|P SPL_IP2_0|SPL2|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|B|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|B|RB SPL_IP2_0|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|I_1|B _PG0_01|P|A1 _PG0_01|P|I_1|MID  2e-12
I_PG0_01|P|I_1|B 0 _PG0_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_3|B _PG0_01|P|A3 _PG0_01|P|I_3|MID  2e-12
I_PG0_01|P|I_3|B 0 _PG0_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|P|I_T|B _PG0_01|P|T1 _PG0_01|P|I_T|MID  2e-12
I_PG0_01|P|I_T|B 0 _PG0_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_6|B _PG0_01|P|Q1 _PG0_01|P|I_6|MID  2e-12
I_PG0_01|P|I_6|B 0 _PG0_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|P|1|1 _PG0_01|P|A1 _PG0_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|1|P _PG0_01|P|1|MID_SERIES 0  2e-13
R_PG0_01|P|1|B _PG0_01|P|A1 _PG0_01|P|1|MID_SHUNT  2.7439617672
L_PG0_01|P|1|RB _PG0_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|23|1 _PG0_01|P|A2 _PG0_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|P|23|B _PG0_01|P|A2 _PG0_01|P|23|MID_SHUNT  3.84154647408
L_PG0_01|P|23|RB _PG0_01|P|23|MID_SHUNT _PG0_01|P|A3  2.1704737578552e-12
B_PG0_01|P|3|1 _PG0_01|P|A3 _PG0_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|3|P _PG0_01|P|3|MID_SERIES 0  2e-13
R_PG0_01|P|3|B _PG0_01|P|A3 _PG0_01|P|3|MID_SHUNT  2.7439617672
L_PG0_01|P|3|RB _PG0_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|4|1 _PG0_01|P|A4 _PG0_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|4|P _PG0_01|P|4|MID_SERIES 0  2e-13
R_PG0_01|P|4|B _PG0_01|P|A4 _PG0_01|P|4|MID_SHUNT  2.7439617672
L_PG0_01|P|4|RB _PG0_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|T|1 _PG0_01|P|T1 _PG0_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|T|P _PG0_01|P|T|MID_SERIES 0  2e-13
R_PG0_01|P|T|B _PG0_01|P|T1 _PG0_01|P|T|MID_SHUNT  2.7439617672
L_PG0_01|P|T|RB _PG0_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|45|1 _PG0_01|P|T2 _PG0_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|P|45|B _PG0_01|P|T2 _PG0_01|P|45|MID_SHUNT  3.84154647408
L_PG0_01|P|45|RB _PG0_01|P|45|MID_SHUNT _PG0_01|P|A4  2.1704737578552e-12
B_PG0_01|P|6|1 _PG0_01|P|Q1 _PG0_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|6|P _PG0_01|P|6|MID_SERIES 0  2e-13
R_PG0_01|P|6|B _PG0_01|P|Q1 _PG0_01|P|6|MID_SHUNT  2.7439617672
L_PG0_01|P|6|RB _PG0_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|G|I_1|B _PG0_01|G|A1 _PG0_01|G|I_1|MID  2e-12
I_PG0_01|G|I_1|B 0 _PG0_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_3|B _PG0_01|G|A3 _PG0_01|G|I_3|MID  2e-12
I_PG0_01|G|I_3|B 0 _PG0_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|G|I_T|B _PG0_01|G|T1 _PG0_01|G|I_T|MID  2e-12
I_PG0_01|G|I_T|B 0 _PG0_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_6|B _PG0_01|G|Q1 _PG0_01|G|I_6|MID  2e-12
I_PG0_01|G|I_6|B 0 _PG0_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|G|1|1 _PG0_01|G|A1 _PG0_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|1|P _PG0_01|G|1|MID_SERIES 0  2e-13
R_PG0_01|G|1|B _PG0_01|G|A1 _PG0_01|G|1|MID_SHUNT  2.7439617672
L_PG0_01|G|1|RB _PG0_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|23|1 _PG0_01|G|A2 _PG0_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|G|23|B _PG0_01|G|A2 _PG0_01|G|23|MID_SHUNT  3.84154647408
L_PG0_01|G|23|RB _PG0_01|G|23|MID_SHUNT _PG0_01|G|A3  2.1704737578552e-12
B_PG0_01|G|3|1 _PG0_01|G|A3 _PG0_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|3|P _PG0_01|G|3|MID_SERIES 0  2e-13
R_PG0_01|G|3|B _PG0_01|G|A3 _PG0_01|G|3|MID_SHUNT  2.7439617672
L_PG0_01|G|3|RB _PG0_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|4|1 _PG0_01|G|A4 _PG0_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|4|P _PG0_01|G|4|MID_SERIES 0  2e-13
R_PG0_01|G|4|B _PG0_01|G|A4 _PG0_01|G|4|MID_SHUNT  2.7439617672
L_PG0_01|G|4|RB _PG0_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|T|1 _PG0_01|G|T1 _PG0_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|T|P _PG0_01|G|T|MID_SERIES 0  2e-13
R_PG0_01|G|T|B _PG0_01|G|T1 _PG0_01|G|T|MID_SHUNT  2.7439617672
L_PG0_01|G|T|RB _PG0_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|45|1 _PG0_01|G|T2 _PG0_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|G|45|B _PG0_01|G|T2 _PG0_01|G|45|MID_SHUNT  3.84154647408
L_PG0_01|G|45|RB _PG0_01|G|45|MID_SHUNT _PG0_01|G|A4  2.1704737578552e-12
B_PG0_01|G|6|1 _PG0_01|G|Q1 _PG0_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|6|P _PG0_01|G|6|MID_SERIES 0  2e-13
R_PG0_01|G|6|B _PG0_01|G|Q1 _PG0_01|G|6|MID_SHUNT  2.7439617672
L_PG0_01|G|6|RB _PG0_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_SPL_G1|I_D1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|I_D1|MID  2e-12
I_PG1_01|_SPL_G1|I_D1|B 0 _PG1_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_D2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|I_D2|MID  2e-12
I_PG1_01|_SPL_G1|I_D2|B 0 _PG1_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG1_01|_SPL_G1|I_Q1|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|I_Q1|MID  2e-12
I_PG1_01|_SPL_G1|I_Q1|B 0 _PG1_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_Q2|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|I_Q2|MID  2e-12
I_PG1_01|_SPL_G1|I_Q2|B 0 _PG1_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG1_01|_SPL_G1|1|1 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|1|P _PG1_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|1|RB _PG1_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|2|1 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|2|P _PG1_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|2|RB _PG1_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|A|1 _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|A|P _PG1_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|A|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|A|RB _PG1_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|B|1 _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|B|P _PG1_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|B|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|B|RB _PG1_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_PG|I_A1|B _PG1_01|_PG|A1 _PG1_01|_PG|I_A1|MID  2e-12
I_PG1_01|_PG|I_A1|B 0 _PG1_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_B1|B _PG1_01|_PG|B1 _PG1_01|_PG|I_B1|MID  2e-12
I_PG1_01|_PG|I_B1|B 0 _PG1_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q3|B _PG1_01|_PG|Q3 _PG1_01|_PG|I_Q3|MID  2e-12
I_PG1_01|_PG|I_Q3|B 0 _PG1_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_PG|I_Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|I_Q2|MID  2e-12
I_PG1_01|_PG|I_Q2|B 0 _PG1_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|I_Q1|MID  2e-12
I_PG1_01|_PG|I_Q1|B 0 _PG1_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_PG|A1|1 _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A1|P _PG1_01|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01|_PG|A1|B _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A1|RB _PG1_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A2|1 _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A2|P _PG1_01|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01|_PG|A2|B _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A2|RB _PG1_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A12|1 _PG1_01|_PG|A2 _PG1_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|A12|B _PG1_01|_PG|A2 _PG1_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|A12|RB _PG1_01|_PG|A12|MID_SHUNT _PG1_01|_PG|A3  2.1704737578552e-12
B_PG1_01|_PG|B1|1 _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B1|P _PG1_01|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01|_PG|B1|B _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B1|RB _PG1_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B2|1 _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B2|P _PG1_01|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01|_PG|B2|B _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B2|RB _PG1_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B12|1 _PG1_01|_PG|B2 _PG1_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|B12|B _PG1_01|_PG|B2 _PG1_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|B12|RB _PG1_01|_PG|B12|MID_SHUNT _PG1_01|_PG|B3  2.1704737578552e-12
B_PG1_01|_PG|Q2|1 _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q2|P _PG1_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q2|RB _PG1_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|Q1|1 _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q1|P _PG1_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q1|RB _PG1_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_GG|I_A1|B _PG1_01|_GG|A1 _PG1_01|_GG|I_A1|MID  2e-12
I_PG1_01|_GG|I_A1|B 0 _PG1_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_B1|B _PG1_01|_GG|B1 _PG1_01|_GG|I_B1|MID  2e-12
I_PG1_01|_GG|I_B1|B 0 _PG1_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q3|B _PG1_01|_GG|Q3 _PG1_01|_GG|I_Q3|MID  2e-12
I_PG1_01|_GG|I_Q3|B 0 _PG1_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_GG|I_Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|I_Q2|MID  2e-12
I_PG1_01|_GG|I_Q2|B 0 _PG1_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|I_Q1|MID  2e-12
I_PG1_01|_GG|I_Q1|B 0 _PG1_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_GG|A1|1 _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A1|P _PG1_01|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01|_GG|A1|B _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A1|RB _PG1_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A2|1 _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A2|P _PG1_01|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01|_GG|A2|B _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A2|RB _PG1_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A12|1 _PG1_01|_GG|A2 _PG1_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|A12|B _PG1_01|_GG|A2 _PG1_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|A12|RB _PG1_01|_GG|A12|MID_SHUNT _PG1_01|_GG|A3  2.1704737578552e-12
B_PG1_01|_GG|B1|1 _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B1|P _PG1_01|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01|_GG|B1|B _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B1|RB _PG1_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B2|1 _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B2|P _PG1_01|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01|_GG|B2|B _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B2|RB _PG1_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B12|1 _PG1_01|_GG|B2 _PG1_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|B12|B _PG1_01|_GG|B2 _PG1_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|B12|RB _PG1_01|_GG|B12|MID_SHUNT _PG1_01|_GG|B3  2.1704737578552e-12
B_PG1_01|_GG|Q2|1 _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q2|P _PG1_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q2|RB _PG1_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|Q1|1 _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q1|P _PG1_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q1|RB _PG1_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_PG|I_1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|I_1|MID  2e-12
I_PG1_01|_DFF_PG|I_1|B 0 _PG1_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|I_3|MID  2e-12
I_PG1_01|_DFF_PG|I_3|B 0 _PG1_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_PG|I_T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|I_T|MID  2e-12
I_PG1_01|_DFF_PG|I_T|B 0 _PG1_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|I_6|MID  2e-12
I_PG1_01|_DFF_PG|I_6|B 0 _PG1_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_PG|1|1 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|1|P _PG1_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|1|RB _PG1_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|23|1 _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|23|B _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|23|RB _PG1_01|_DFF_PG|23|MID_SHUNT _PG1_01|_DFF_PG|A3  2.1704737578552e-12
B_PG1_01|_DFF_PG|3|1 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|3|P _PG1_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|3|RB _PG1_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|4|1 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|4|P _PG1_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|4|B _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|4|RB _PG1_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|T|1 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|T|P _PG1_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|T|RB _PG1_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|45|1 _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|45|B _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|45|RB _PG1_01|_DFF_PG|45|MID_SHUNT _PG1_01|_DFF_PG|A4  2.1704737578552e-12
B_PG1_01|_DFF_PG|6|1 _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|6|P _PG1_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|6|RB _PG1_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_GG|I_1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|I_1|MID  2e-12
I_PG1_01|_DFF_GG|I_1|B 0 _PG1_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|I_3|MID  2e-12
I_PG1_01|_DFF_GG|I_3|B 0 _PG1_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_GG|I_T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|I_T|MID  2e-12
I_PG1_01|_DFF_GG|I_T|B 0 _PG1_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|I_6|MID  2e-12
I_PG1_01|_DFF_GG|I_6|B 0 _PG1_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_GG|1|1 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|1|P _PG1_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|1|RB _PG1_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|23|1 _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|23|B _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|23|RB _PG1_01|_DFF_GG|23|MID_SHUNT _PG1_01|_DFF_GG|A3  2.1704737578552e-12
B_PG1_01|_DFF_GG|3|1 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|3|P _PG1_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|3|RB _PG1_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|4|1 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|4|P _PG1_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|4|B _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|4|RB _PG1_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|T|1 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|T|P _PG1_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|T|RB _PG1_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|45|1 _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|45|B _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|45|RB _PG1_01|_DFF_GG|45|MID_SHUNT _PG1_01|_DFF_GG|A4  2.1704737578552e-12
B_PG1_01|_DFF_GG|6|1 _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|6|P _PG1_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|6|RB _PG1_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_G|I_A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|I_A1|MID  2e-12
I_PG1_01|_AND_G|I_A1|B 0 _PG1_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|I_B1|MID  2e-12
I_PG1_01|_AND_G|I_B1|B 0 _PG1_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q3|B _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|I_Q3|MID  2e-12
I_PG1_01|_AND_G|I_Q3|B 0 _PG1_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_G|I_Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|I_Q2|MID  2e-12
I_PG1_01|_AND_G|I_Q2|B 0 _PG1_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|I_Q1|MID  2e-12
I_PG1_01|_AND_G|I_Q1|B 0 _PG1_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_G|A1|1 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A1|P _PG1_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A1|RB _PG1_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A2|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A2|P _PG1_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A2|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A2|RB _PG1_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A12|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|A12|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|A12|RB _PG1_01|_AND_G|A12|MID_SHUNT _PG1_01|_AND_G|A3  2.1704737578552e-12
B_PG1_01|_AND_G|B1|1 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B1|P _PG1_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B1|RB _PG1_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B2|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B2|P _PG1_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B2|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B2|RB _PG1_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B12|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|B12|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|B12|RB _PG1_01|_AND_G|B12|MID_SHUNT _PG1_01|_AND_G|B3  2.1704737578552e-12
B_PG1_01|_AND_G|Q2|1 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q2|P _PG1_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q2|RB _PG1_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|Q1|1 _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q1|P _PG1_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q1|RB _PG1_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|P|I_1|B _PG2_01|P|A1 _PG2_01|P|I_1|MID  2e-12
I_PG2_01|P|I_1|B 0 _PG2_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_3|B _PG2_01|P|A3 _PG2_01|P|I_3|MID  2e-12
I_PG2_01|P|I_3|B 0 _PG2_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|P|I_T|B _PG2_01|P|T1 _PG2_01|P|I_T|MID  2e-12
I_PG2_01|P|I_T|B 0 _PG2_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_6|B _PG2_01|P|Q1 _PG2_01|P|I_6|MID  2e-12
I_PG2_01|P|I_6|B 0 _PG2_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|P|1|1 _PG2_01|P|A1 _PG2_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|1|P _PG2_01|P|1|MID_SERIES 0  2e-13
R_PG2_01|P|1|B _PG2_01|P|A1 _PG2_01|P|1|MID_SHUNT  2.7439617672
L_PG2_01|P|1|RB _PG2_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|23|1 _PG2_01|P|A2 _PG2_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|P|23|B _PG2_01|P|A2 _PG2_01|P|23|MID_SHUNT  3.84154647408
L_PG2_01|P|23|RB _PG2_01|P|23|MID_SHUNT _PG2_01|P|A3  2.1704737578552e-12
B_PG2_01|P|3|1 _PG2_01|P|A3 _PG2_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|3|P _PG2_01|P|3|MID_SERIES 0  2e-13
R_PG2_01|P|3|B _PG2_01|P|A3 _PG2_01|P|3|MID_SHUNT  2.7439617672
L_PG2_01|P|3|RB _PG2_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|4|1 _PG2_01|P|A4 _PG2_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|4|P _PG2_01|P|4|MID_SERIES 0  2e-13
R_PG2_01|P|4|B _PG2_01|P|A4 _PG2_01|P|4|MID_SHUNT  2.7439617672
L_PG2_01|P|4|RB _PG2_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|T|1 _PG2_01|P|T1 _PG2_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|T|P _PG2_01|P|T|MID_SERIES 0  2e-13
R_PG2_01|P|T|B _PG2_01|P|T1 _PG2_01|P|T|MID_SHUNT  2.7439617672
L_PG2_01|P|T|RB _PG2_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|45|1 _PG2_01|P|T2 _PG2_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|P|45|B _PG2_01|P|T2 _PG2_01|P|45|MID_SHUNT  3.84154647408
L_PG2_01|P|45|RB _PG2_01|P|45|MID_SHUNT _PG2_01|P|A4  2.1704737578552e-12
B_PG2_01|P|6|1 _PG2_01|P|Q1 _PG2_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|6|P _PG2_01|P|6|MID_SERIES 0  2e-13
R_PG2_01|P|6|B _PG2_01|P|Q1 _PG2_01|P|6|MID_SHUNT  2.7439617672
L_PG2_01|P|6|RB _PG2_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|G|I_1|B _PG2_01|G|A1 _PG2_01|G|I_1|MID  2e-12
I_PG2_01|G|I_1|B 0 _PG2_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_3|B _PG2_01|G|A3 _PG2_01|G|I_3|MID  2e-12
I_PG2_01|G|I_3|B 0 _PG2_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|G|I_T|B _PG2_01|G|T1 _PG2_01|G|I_T|MID  2e-12
I_PG2_01|G|I_T|B 0 _PG2_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_6|B _PG2_01|G|Q1 _PG2_01|G|I_6|MID  2e-12
I_PG2_01|G|I_6|B 0 _PG2_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|G|1|1 _PG2_01|G|A1 _PG2_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|1|P _PG2_01|G|1|MID_SERIES 0  2e-13
R_PG2_01|G|1|B _PG2_01|G|A1 _PG2_01|G|1|MID_SHUNT  2.7439617672
L_PG2_01|G|1|RB _PG2_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|23|1 _PG2_01|G|A2 _PG2_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|G|23|B _PG2_01|G|A2 _PG2_01|G|23|MID_SHUNT  3.84154647408
L_PG2_01|G|23|RB _PG2_01|G|23|MID_SHUNT _PG2_01|G|A3  2.1704737578552e-12
B_PG2_01|G|3|1 _PG2_01|G|A3 _PG2_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|3|P _PG2_01|G|3|MID_SERIES 0  2e-13
R_PG2_01|G|3|B _PG2_01|G|A3 _PG2_01|G|3|MID_SHUNT  2.7439617672
L_PG2_01|G|3|RB _PG2_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|4|1 _PG2_01|G|A4 _PG2_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|4|P _PG2_01|G|4|MID_SERIES 0  2e-13
R_PG2_01|G|4|B _PG2_01|G|A4 _PG2_01|G|4|MID_SHUNT  2.7439617672
L_PG2_01|G|4|RB _PG2_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|T|1 _PG2_01|G|T1 _PG2_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|T|P _PG2_01|G|T|MID_SERIES 0  2e-13
R_PG2_01|G|T|B _PG2_01|G|T1 _PG2_01|G|T|MID_SHUNT  2.7439617672
L_PG2_01|G|T|RB _PG2_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|45|1 _PG2_01|G|T2 _PG2_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|G|45|B _PG2_01|G|T2 _PG2_01|G|45|MID_SHUNT  3.84154647408
L_PG2_01|G|45|RB _PG2_01|G|45|MID_SHUNT _PG2_01|G|A4  2.1704737578552e-12
B_PG2_01|G|6|1 _PG2_01|G|Q1 _PG2_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|6|P _PG2_01|G|6|MID_SERIES 0  2e-13
R_PG2_01|G|6|B _PG2_01|G|Q1 _PG2_01|G|6|MID_SHUNT  2.7439617672
L_PG2_01|G|6|RB _PG2_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_G1|I_D1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|I_D1|MID  2e-12
I_PG3_01|_SPL_G1|I_D1|B 0 _PG3_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_D2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|I_D2|MID  2e-12
I_PG3_01|_SPL_G1|I_D2|B 0 _PG3_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_G1|I_Q1|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|I_Q1|MID  2e-12
I_PG3_01|_SPL_G1|I_Q1|B 0 _PG3_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_Q2|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|I_Q2|MID  2e-12
I_PG3_01|_SPL_G1|I_Q2|B 0 _PG3_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_G1|1|1 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|1|P _PG3_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|1|RB _PG3_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|2|1 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|2|P _PG3_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|2|RB _PG3_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|A|1 _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|A|P _PG3_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|A|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|A|RB _PG3_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|B|1 _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|B|P _PG3_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|B|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|B|RB _PG3_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_P1|I_D1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|I_D1|MID  2e-12
I_PG3_01|_SPL_P1|I_D1|B 0 _PG3_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_D2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|I_D2|MID  2e-12
I_PG3_01|_SPL_P1|I_D2|B 0 _PG3_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_P1|I_Q1|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|I_Q1|MID  2e-12
I_PG3_01|_SPL_P1|I_Q1|B 0 _PG3_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_Q2|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|I_Q2|MID  2e-12
I_PG3_01|_SPL_P1|I_Q2|B 0 _PG3_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_P1|1|1 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|1|P _PG3_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|1|RB _PG3_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|2|1 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|2|P _PG3_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|2|RB _PG3_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|A|1 _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|A|P _PG3_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|A|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|A|RB _PG3_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|B|1 _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|B|P _PG3_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|B|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|B|RB _PG3_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_PG|I_A1|B _PG3_01|_PG|A1 _PG3_01|_PG|I_A1|MID  2e-12
I_PG3_01|_PG|I_A1|B 0 _PG3_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_B1|B _PG3_01|_PG|B1 _PG3_01|_PG|I_B1|MID  2e-12
I_PG3_01|_PG|I_B1|B 0 _PG3_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q3|B _PG3_01|_PG|Q3 _PG3_01|_PG|I_Q3|MID  2e-12
I_PG3_01|_PG|I_Q3|B 0 _PG3_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_PG|I_Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|I_Q2|MID  2e-12
I_PG3_01|_PG|I_Q2|B 0 _PG3_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|I_Q1|MID  2e-12
I_PG3_01|_PG|I_Q1|B 0 _PG3_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_PG|A1|1 _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A1|P _PG3_01|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01|_PG|A1|B _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A1|RB _PG3_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A2|1 _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A2|P _PG3_01|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01|_PG|A2|B _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A2|RB _PG3_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A12|1 _PG3_01|_PG|A2 _PG3_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|A12|B _PG3_01|_PG|A2 _PG3_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|A12|RB _PG3_01|_PG|A12|MID_SHUNT _PG3_01|_PG|A3  2.1704737578552e-12
B_PG3_01|_PG|B1|1 _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B1|P _PG3_01|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01|_PG|B1|B _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B1|RB _PG3_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B2|1 _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B2|P _PG3_01|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01|_PG|B2|B _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B2|RB _PG3_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B12|1 _PG3_01|_PG|B2 _PG3_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|B12|B _PG3_01|_PG|B2 _PG3_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|B12|RB _PG3_01|_PG|B12|MID_SHUNT _PG3_01|_PG|B3  2.1704737578552e-12
B_PG3_01|_PG|Q2|1 _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q2|P _PG3_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q2|RB _PG3_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|Q1|1 _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q1|P _PG3_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q1|RB _PG3_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_GG|I_A1|B _PG3_01|_GG|A1 _PG3_01|_GG|I_A1|MID  2e-12
I_PG3_01|_GG|I_A1|B 0 _PG3_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_B1|B _PG3_01|_GG|B1 _PG3_01|_GG|I_B1|MID  2e-12
I_PG3_01|_GG|I_B1|B 0 _PG3_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q3|B _PG3_01|_GG|Q3 _PG3_01|_GG|I_Q3|MID  2e-12
I_PG3_01|_GG|I_Q3|B 0 _PG3_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_GG|I_Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|I_Q2|MID  2e-12
I_PG3_01|_GG|I_Q2|B 0 _PG3_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|I_Q1|MID  2e-12
I_PG3_01|_GG|I_Q1|B 0 _PG3_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_GG|A1|1 _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A1|P _PG3_01|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01|_GG|A1|B _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A1|RB _PG3_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A2|1 _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A2|P _PG3_01|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01|_GG|A2|B _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A2|RB _PG3_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A12|1 _PG3_01|_GG|A2 _PG3_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|A12|B _PG3_01|_GG|A2 _PG3_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|A12|RB _PG3_01|_GG|A12|MID_SHUNT _PG3_01|_GG|A3  2.1704737578552e-12
B_PG3_01|_GG|B1|1 _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B1|P _PG3_01|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01|_GG|B1|B _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B1|RB _PG3_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B2|1 _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B2|P _PG3_01|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01|_GG|B2|B _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B2|RB _PG3_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B12|1 _PG3_01|_GG|B2 _PG3_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|B12|B _PG3_01|_GG|B2 _PG3_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|B12|RB _PG3_01|_GG|B12|MID_SHUNT _PG3_01|_GG|B3  2.1704737578552e-12
B_PG3_01|_GG|Q2|1 _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q2|P _PG3_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q2|RB _PG3_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|Q1|1 _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q1|P _PG3_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q1|RB _PG3_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P0|I_1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|I_1|MID  2e-12
I_PG3_01|_DFF_P0|I_1|B 0 _PG3_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|I_3|MID  2e-12
I_PG3_01|_DFF_P0|I_3|B 0 _PG3_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P0|I_T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|I_T|MID  2e-12
I_PG3_01|_DFF_P0|I_T|B 0 _PG3_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|I_6|MID  2e-12
I_PG3_01|_DFF_P0|I_6|B 0 _PG3_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P0|1|1 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|1|P _PG3_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|1|RB _PG3_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|23|1 _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|23|B _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|23|RB _PG3_01|_DFF_P0|23|MID_SHUNT _PG3_01|_DFF_P0|A3  2.1704737578552e-12
B_PG3_01|_DFF_P0|3|1 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|3|P _PG3_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|3|RB _PG3_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|4|1 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|4|P _PG3_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|4|B _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|4|RB _PG3_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|T|1 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|T|P _PG3_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|T|RB _PG3_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|45|1 _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|45|B _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|45|RB _PG3_01|_DFF_P0|45|MID_SHUNT _PG3_01|_DFF_P0|A4  2.1704737578552e-12
B_PG3_01|_DFF_P0|6|1 _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|6|P _PG3_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|6|RB _PG3_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P1|I_1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|I_1|MID  2e-12
I_PG3_01|_DFF_P1|I_1|B 0 _PG3_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|I_3|MID  2e-12
I_PG3_01|_DFF_P1|I_3|B 0 _PG3_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P1|I_T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|I_T|MID  2e-12
I_PG3_01|_DFF_P1|I_T|B 0 _PG3_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|I_6|MID  2e-12
I_PG3_01|_DFF_P1|I_6|B 0 _PG3_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P1|1|1 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|1|P _PG3_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|1|RB _PG3_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|23|1 _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|23|B _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|23|RB _PG3_01|_DFF_P1|23|MID_SHUNT _PG3_01|_DFF_P1|A3  2.1704737578552e-12
B_PG3_01|_DFF_P1|3|1 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|3|P _PG3_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|3|RB _PG3_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|4|1 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|4|P _PG3_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|4|B _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|4|RB _PG3_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|T|1 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|T|P _PG3_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|T|RB _PG3_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|45|1 _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|45|B _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|45|RB _PG3_01|_DFF_P1|45|MID_SHUNT _PG3_01|_DFF_P1|A4  2.1704737578552e-12
B_PG3_01|_DFF_P1|6|1 _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|6|P _PG3_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|6|RB _PG3_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_PG|I_1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|I_1|MID  2e-12
I_PG3_01|_DFF_PG|I_1|B 0 _PG3_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|I_3|MID  2e-12
I_PG3_01|_DFF_PG|I_3|B 0 _PG3_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_PG|I_T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|I_T|MID  2e-12
I_PG3_01|_DFF_PG|I_T|B 0 _PG3_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|I_6|MID  2e-12
I_PG3_01|_DFF_PG|I_6|B 0 _PG3_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_PG|1|1 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|1|P _PG3_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|1|RB _PG3_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|23|1 _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|23|B _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|23|RB _PG3_01|_DFF_PG|23|MID_SHUNT _PG3_01|_DFF_PG|A3  2.1704737578552e-12
B_PG3_01|_DFF_PG|3|1 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|3|P _PG3_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|3|RB _PG3_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|4|1 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|4|P _PG3_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|4|B _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|4|RB _PG3_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|T|1 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|T|P _PG3_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|T|RB _PG3_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|45|1 _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|45|B _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|45|RB _PG3_01|_DFF_PG|45|MID_SHUNT _PG3_01|_DFF_PG|A4  2.1704737578552e-12
B_PG3_01|_DFF_PG|6|1 _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|6|P _PG3_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|6|RB _PG3_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_GG|I_1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|I_1|MID  2e-12
I_PG3_01|_DFF_GG|I_1|B 0 _PG3_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|I_3|MID  2e-12
I_PG3_01|_DFF_GG|I_3|B 0 _PG3_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_GG|I_T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|I_T|MID  2e-12
I_PG3_01|_DFF_GG|I_T|B 0 _PG3_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|I_6|MID  2e-12
I_PG3_01|_DFF_GG|I_6|B 0 _PG3_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_GG|1|1 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|1|P _PG3_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|1|RB _PG3_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|23|1 _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|23|B _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|23|RB _PG3_01|_DFF_GG|23|MID_SHUNT _PG3_01|_DFF_GG|A3  2.1704737578552e-12
B_PG3_01|_DFF_GG|3|1 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|3|P _PG3_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|3|RB _PG3_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|4|1 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|4|P _PG3_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|4|B _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|4|RB _PG3_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|T|1 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|T|P _PG3_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|T|RB _PG3_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|45|1 _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|45|B _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|45|RB _PG3_01|_DFF_GG|45|MID_SHUNT _PG3_01|_DFF_GG|A4  2.1704737578552e-12
B_PG3_01|_DFF_GG|6|1 _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|6|P _PG3_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|6|RB _PG3_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_G|I_A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|I_A1|MID  2e-12
I_PG3_01|_AND_G|I_A1|B 0 _PG3_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|I_B1|MID  2e-12
I_PG3_01|_AND_G|I_B1|B 0 _PG3_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q3|B _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|I_Q3|MID  2e-12
I_PG3_01|_AND_G|I_Q3|B 0 _PG3_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_G|I_Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|I_Q2|MID  2e-12
I_PG3_01|_AND_G|I_Q2|B 0 _PG3_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|I_Q1|MID  2e-12
I_PG3_01|_AND_G|I_Q1|B 0 _PG3_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_G|A1|1 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A1|P _PG3_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A1|RB _PG3_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A2|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A2|P _PG3_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A2|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A2|RB _PG3_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A12|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|A12|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|A12|RB _PG3_01|_AND_G|A12|MID_SHUNT _PG3_01|_AND_G|A3  2.1704737578552e-12
B_PG3_01|_AND_G|B1|1 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B1|P _PG3_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B1|RB _PG3_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B2|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B2|P _PG3_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B2|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B2|RB _PG3_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B12|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|B12|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|B12|RB _PG3_01|_AND_G|B12|MID_SHUNT _PG3_01|_AND_G|B3  2.1704737578552e-12
B_PG3_01|_AND_G|Q2|1 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q2|P _PG3_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q2|RB _PG3_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|Q1|1 _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q1|P _PG3_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q1|RB _PG3_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_P|I_A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|I_A1|MID  2e-12
I_PG3_01|_AND_P|I_A1|B 0 _PG3_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|I_B1|MID  2e-12
I_PG3_01|_AND_P|I_B1|B 0 _PG3_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q3|B _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|I_Q3|MID  2e-12
I_PG3_01|_AND_P|I_Q3|B 0 _PG3_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_P|I_Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|I_Q2|MID  2e-12
I_PG3_01|_AND_P|I_Q2|B 0 _PG3_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|I_Q1|MID  2e-12
I_PG3_01|_AND_P|I_Q1|B 0 _PG3_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_P|A1|1 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A1|P _PG3_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A1|RB _PG3_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A2|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A2|P _PG3_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A2|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A2|RB _PG3_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A12|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|A12|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|A12|RB _PG3_01|_AND_P|A12|MID_SHUNT _PG3_01|_AND_P|A3  2.1704737578552e-12
B_PG3_01|_AND_P|B1|1 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B1|P _PG3_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B1|RB _PG3_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B2|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B2|P _PG3_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B2|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B2|RB _PG3_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B12|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|B12|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|B12|RB _PG3_01|_AND_P|B12|MID_SHUNT _PG3_01|_AND_P|B3  2.1704737578552e-12
B_PG3_01|_AND_P|Q2|1 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q2|P _PG3_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q2|RB _PG3_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|Q1|1 _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q1|P _PG3_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q1|RB _PG3_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL1|I_D1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|I_D1|MID  2e-12
ISPL_G1_1|SPL1|I_D1|B 0 SPL_G1_1|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_D2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|I_D2|MID  2e-12
ISPL_G1_1|SPL1|I_D2|B 0 SPL_G1_1|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL1|I_Q1|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|I_Q1|MID  2e-12
ISPL_G1_1|SPL1|I_Q1|B 0 SPL_G1_1|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_Q2|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|I_Q2|MID  2e-12
ISPL_G1_1|SPL1|I_Q2|B 0 SPL_G1_1|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL1|1|1 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|1|P SPL_G1_1|SPL1|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|1|RB SPL_G1_1|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|2|1 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|2|P SPL_G1_1|SPL1|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|2|RB SPL_G1_1|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|A|1 SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|A|P SPL_G1_1|SPL1|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|A|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|A|RB SPL_G1_1|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|B|1 SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|B|P SPL_G1_1|SPL1|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|B|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|B|RB SPL_G1_1|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL2|I_D1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|I_D1|MID  2e-12
ISPL_G1_1|SPL2|I_D1|B 0 SPL_G1_1|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_D2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|I_D2|MID  2e-12
ISPL_G1_1|SPL2|I_D2|B 0 SPL_G1_1|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL2|I_Q1|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|I_Q1|MID  2e-12
ISPL_G1_1|SPL2|I_Q1|B 0 SPL_G1_1|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_Q2|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|I_Q2|MID  2e-12
ISPL_G1_1|SPL2|I_Q2|B 0 SPL_G1_1|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL2|1|1 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|1|P SPL_G1_1|SPL2|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|1|RB SPL_G1_1|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|2|1 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|2|P SPL_G1_1|SPL2|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|2|RB SPL_G1_1|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|A|1 SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|A|P SPL_G1_1|SPL2|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|A|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|A|RB SPL_G1_1|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|B|1 SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|B|P SPL_G1_1|SPL2|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|B|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|B|RB SPL_G1_1|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|P|I_1|B _PG0_12|P|A1 _PG0_12|P|I_1|MID  2e-12
I_PG0_12|P|I_1|B 0 _PG0_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_3|B _PG0_12|P|A3 _PG0_12|P|I_3|MID  2e-12
I_PG0_12|P|I_3|B 0 _PG0_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|P|I_T|B _PG0_12|P|T1 _PG0_12|P|I_T|MID  2e-12
I_PG0_12|P|I_T|B 0 _PG0_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_6|B _PG0_12|P|Q1 _PG0_12|P|I_6|MID  2e-12
I_PG0_12|P|I_6|B 0 _PG0_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|P|1|1 _PG0_12|P|A1 _PG0_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|1|P _PG0_12|P|1|MID_SERIES 0  2e-13
R_PG0_12|P|1|B _PG0_12|P|A1 _PG0_12|P|1|MID_SHUNT  2.7439617672
L_PG0_12|P|1|RB _PG0_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|23|1 _PG0_12|P|A2 _PG0_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|P|23|B _PG0_12|P|A2 _PG0_12|P|23|MID_SHUNT  3.84154647408
L_PG0_12|P|23|RB _PG0_12|P|23|MID_SHUNT _PG0_12|P|A3  2.1704737578552e-12
B_PG0_12|P|3|1 _PG0_12|P|A3 _PG0_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|3|P _PG0_12|P|3|MID_SERIES 0  2e-13
R_PG0_12|P|3|B _PG0_12|P|A3 _PG0_12|P|3|MID_SHUNT  2.7439617672
L_PG0_12|P|3|RB _PG0_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|4|1 _PG0_12|P|A4 _PG0_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|4|P _PG0_12|P|4|MID_SERIES 0  2e-13
R_PG0_12|P|4|B _PG0_12|P|A4 _PG0_12|P|4|MID_SHUNT  2.7439617672
L_PG0_12|P|4|RB _PG0_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|T|1 _PG0_12|P|T1 _PG0_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|T|P _PG0_12|P|T|MID_SERIES 0  2e-13
R_PG0_12|P|T|B _PG0_12|P|T1 _PG0_12|P|T|MID_SHUNT  2.7439617672
L_PG0_12|P|T|RB _PG0_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|45|1 _PG0_12|P|T2 _PG0_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|P|45|B _PG0_12|P|T2 _PG0_12|P|45|MID_SHUNT  3.84154647408
L_PG0_12|P|45|RB _PG0_12|P|45|MID_SHUNT _PG0_12|P|A4  2.1704737578552e-12
B_PG0_12|P|6|1 _PG0_12|P|Q1 _PG0_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|6|P _PG0_12|P|6|MID_SERIES 0  2e-13
R_PG0_12|P|6|B _PG0_12|P|Q1 _PG0_12|P|6|MID_SHUNT  2.7439617672
L_PG0_12|P|6|RB _PG0_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|G|I_1|B _PG0_12|G|A1 _PG0_12|G|I_1|MID  2e-12
I_PG0_12|G|I_1|B 0 _PG0_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_3|B _PG0_12|G|A3 _PG0_12|G|I_3|MID  2e-12
I_PG0_12|G|I_3|B 0 _PG0_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|G|I_T|B _PG0_12|G|T1 _PG0_12|G|I_T|MID  2e-12
I_PG0_12|G|I_T|B 0 _PG0_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_6|B _PG0_12|G|Q1 _PG0_12|G|I_6|MID  2e-12
I_PG0_12|G|I_6|B 0 _PG0_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|G|1|1 _PG0_12|G|A1 _PG0_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|1|P _PG0_12|G|1|MID_SERIES 0  2e-13
R_PG0_12|G|1|B _PG0_12|G|A1 _PG0_12|G|1|MID_SHUNT  2.7439617672
L_PG0_12|G|1|RB _PG0_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|23|1 _PG0_12|G|A2 _PG0_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|G|23|B _PG0_12|G|A2 _PG0_12|G|23|MID_SHUNT  3.84154647408
L_PG0_12|G|23|RB _PG0_12|G|23|MID_SHUNT _PG0_12|G|A3  2.1704737578552e-12
B_PG0_12|G|3|1 _PG0_12|G|A3 _PG0_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|3|P _PG0_12|G|3|MID_SERIES 0  2e-13
R_PG0_12|G|3|B _PG0_12|G|A3 _PG0_12|G|3|MID_SHUNT  2.7439617672
L_PG0_12|G|3|RB _PG0_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|4|1 _PG0_12|G|A4 _PG0_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|4|P _PG0_12|G|4|MID_SERIES 0  2e-13
R_PG0_12|G|4|B _PG0_12|G|A4 _PG0_12|G|4|MID_SHUNT  2.7439617672
L_PG0_12|G|4|RB _PG0_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|T|1 _PG0_12|G|T1 _PG0_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|T|P _PG0_12|G|T|MID_SERIES 0  2e-13
R_PG0_12|G|T|B _PG0_12|G|T1 _PG0_12|G|T|MID_SHUNT  2.7439617672
L_PG0_12|G|T|RB _PG0_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|45|1 _PG0_12|G|T2 _PG0_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|G|45|B _PG0_12|G|T2 _PG0_12|G|45|MID_SHUNT  3.84154647408
L_PG0_12|G|45|RB _PG0_12|G|45|MID_SHUNT _PG0_12|G|A4  2.1704737578552e-12
B_PG0_12|G|6|1 _PG0_12|G|Q1 _PG0_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|6|P _PG0_12|G|6|MID_SERIES 0  2e-13
R_PG0_12|G|6|B _PG0_12|G|Q1 _PG0_12|G|6|MID_SHUNT  2.7439617672
L_PG0_12|G|6|RB _PG0_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|I_D1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|I_D1|MID  2e-12
I_PG2_12|_SPL_G1|I_D1|B 0 _PG2_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_D2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|I_D2|MID  2e-12
I_PG2_12|_SPL_G1|I_D2|B 0 _PG2_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG2_12|_SPL_G1|I_Q1|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|I_Q1|MID  2e-12
I_PG2_12|_SPL_G1|I_Q1|B 0 _PG2_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_Q2|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|I_Q2|MID  2e-12
I_PG2_12|_SPL_G1|I_Q2|B 0 _PG2_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG2_12|_SPL_G1|1|1 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|1|P _PG2_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|1|RB _PG2_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|2|1 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|2|P _PG2_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|2|RB _PG2_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|A|1 _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|A|P _PG2_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|A|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|A|RB _PG2_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|B|1 _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|B|P _PG2_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|B|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|B|RB _PG2_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_PG|I_A1|B _PG2_12|_PG|A1 _PG2_12|_PG|I_A1|MID  2e-12
I_PG2_12|_PG|I_A1|B 0 _PG2_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_B1|B _PG2_12|_PG|B1 _PG2_12|_PG|I_B1|MID  2e-12
I_PG2_12|_PG|I_B1|B 0 _PG2_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q3|B _PG2_12|_PG|Q3 _PG2_12|_PG|I_Q3|MID  2e-12
I_PG2_12|_PG|I_Q3|B 0 _PG2_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_PG|I_Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|I_Q2|MID  2e-12
I_PG2_12|_PG|I_Q2|B 0 _PG2_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|I_Q1|MID  2e-12
I_PG2_12|_PG|I_Q1|B 0 _PG2_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_PG|A1|1 _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A1|P _PG2_12|_PG|A1|MID_SERIES 0  2e-13
R_PG2_12|_PG|A1|B _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A1|RB _PG2_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A2|1 _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A2|P _PG2_12|_PG|A2|MID_SERIES 0  2e-13
R_PG2_12|_PG|A2|B _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A2|RB _PG2_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A12|1 _PG2_12|_PG|A2 _PG2_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|A12|B _PG2_12|_PG|A2 _PG2_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|A12|RB _PG2_12|_PG|A12|MID_SHUNT _PG2_12|_PG|A3  2.1704737578552e-12
B_PG2_12|_PG|B1|1 _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B1|P _PG2_12|_PG|B1|MID_SERIES 0  2e-13
R_PG2_12|_PG|B1|B _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B1|RB _PG2_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B2|1 _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B2|P _PG2_12|_PG|B2|MID_SERIES 0  2e-13
R_PG2_12|_PG|B2|B _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B2|RB _PG2_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B12|1 _PG2_12|_PG|B2 _PG2_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|B12|B _PG2_12|_PG|B2 _PG2_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|B12|RB _PG2_12|_PG|B12|MID_SHUNT _PG2_12|_PG|B3  2.1704737578552e-12
B_PG2_12|_PG|Q2|1 _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q2|P _PG2_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q2|RB _PG2_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|Q1|1 _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q1|P _PG2_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q1|RB _PG2_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_GG|I_A1|B _PG2_12|_GG|A1 _PG2_12|_GG|I_A1|MID  2e-12
I_PG2_12|_GG|I_A1|B 0 _PG2_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_B1|B _PG2_12|_GG|B1 _PG2_12|_GG|I_B1|MID  2e-12
I_PG2_12|_GG|I_B1|B 0 _PG2_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q3|B _PG2_12|_GG|Q3 _PG2_12|_GG|I_Q3|MID  2e-12
I_PG2_12|_GG|I_Q3|B 0 _PG2_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_GG|I_Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|I_Q2|MID  2e-12
I_PG2_12|_GG|I_Q2|B 0 _PG2_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|I_Q1|MID  2e-12
I_PG2_12|_GG|I_Q1|B 0 _PG2_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_GG|A1|1 _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A1|P _PG2_12|_GG|A1|MID_SERIES 0  2e-13
R_PG2_12|_GG|A1|B _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A1|RB _PG2_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A2|1 _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A2|P _PG2_12|_GG|A2|MID_SERIES 0  2e-13
R_PG2_12|_GG|A2|B _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A2|RB _PG2_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A12|1 _PG2_12|_GG|A2 _PG2_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|A12|B _PG2_12|_GG|A2 _PG2_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|A12|RB _PG2_12|_GG|A12|MID_SHUNT _PG2_12|_GG|A3  2.1704737578552e-12
B_PG2_12|_GG|B1|1 _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B1|P _PG2_12|_GG|B1|MID_SERIES 0  2e-13
R_PG2_12|_GG|B1|B _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B1|RB _PG2_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B2|1 _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B2|P _PG2_12|_GG|B2|MID_SERIES 0  2e-13
R_PG2_12|_GG|B2|B _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B2|RB _PG2_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B12|1 _PG2_12|_GG|B2 _PG2_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|B12|B _PG2_12|_GG|B2 _PG2_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|B12|RB _PG2_12|_GG|B12|MID_SHUNT _PG2_12|_GG|B3  2.1704737578552e-12
B_PG2_12|_GG|Q2|1 _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q2|P _PG2_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q2|RB _PG2_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|Q1|1 _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q1|P _PG2_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q1|RB _PG2_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_PG|I_1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|I_1|MID  2e-12
I_PG2_12|_DFF_PG|I_1|B 0 _PG2_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|I_3|MID  2e-12
I_PG2_12|_DFF_PG|I_3|B 0 _PG2_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_PG|I_T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|I_T|MID  2e-12
I_PG2_12|_DFF_PG|I_T|B 0 _PG2_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|I_6|MID  2e-12
I_PG2_12|_DFF_PG|I_6|B 0 _PG2_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_PG|1|1 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|1|P _PG2_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|1|RB _PG2_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|23|1 _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|23|B _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|23|RB _PG2_12|_DFF_PG|23|MID_SHUNT _PG2_12|_DFF_PG|A3  2.1704737578552e-12
B_PG2_12|_DFF_PG|3|1 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|3|P _PG2_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|3|RB _PG2_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|4|1 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|4|P _PG2_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|4|B _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|4|RB _PG2_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|T|1 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|T|P _PG2_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|T|RB _PG2_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|45|1 _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|45|B _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|45|RB _PG2_12|_DFF_PG|45|MID_SHUNT _PG2_12|_DFF_PG|A4  2.1704737578552e-12
B_PG2_12|_DFF_PG|6|1 _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|6|P _PG2_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|6|RB _PG2_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_GG|I_1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|I_1|MID  2e-12
I_PG2_12|_DFF_GG|I_1|B 0 _PG2_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|I_3|MID  2e-12
I_PG2_12|_DFF_GG|I_3|B 0 _PG2_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_GG|I_T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|I_T|MID  2e-12
I_PG2_12|_DFF_GG|I_T|B 0 _PG2_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|I_6|MID  2e-12
I_PG2_12|_DFF_GG|I_6|B 0 _PG2_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_GG|1|1 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|1|P _PG2_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|1|RB _PG2_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|23|1 _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|23|B _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|23|RB _PG2_12|_DFF_GG|23|MID_SHUNT _PG2_12|_DFF_GG|A3  2.1704737578552e-12
B_PG2_12|_DFF_GG|3|1 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|3|P _PG2_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|3|RB _PG2_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|4|1 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|4|P _PG2_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|4|B _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|4|RB _PG2_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|T|1 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|T|P _PG2_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|T|RB _PG2_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|45|1 _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|45|B _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|45|RB _PG2_12|_DFF_GG|45|MID_SHUNT _PG2_12|_DFF_GG|A4  2.1704737578552e-12
B_PG2_12|_DFF_GG|6|1 _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|6|P _PG2_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|6|RB _PG2_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_G|I_A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|I_A1|MID  2e-12
I_PG2_12|_AND_G|I_A1|B 0 _PG2_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|I_B1|MID  2e-12
I_PG2_12|_AND_G|I_B1|B 0 _PG2_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q3|B _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|I_Q3|MID  2e-12
I_PG2_12|_AND_G|I_Q3|B 0 _PG2_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_G|I_Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|I_Q2|MID  2e-12
I_PG2_12|_AND_G|I_Q2|B 0 _PG2_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|I_Q1|MID  2e-12
I_PG2_12|_AND_G|I_Q1|B 0 _PG2_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_G|A1|1 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A1|P _PG2_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A1|RB _PG2_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A2|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A2|P _PG2_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A2|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A2|RB _PG2_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A12|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|A12|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|A12|RB _PG2_12|_AND_G|A12|MID_SHUNT _PG2_12|_AND_G|A3  2.1704737578552e-12
B_PG2_12|_AND_G|B1|1 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B1|P _PG2_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B1|RB _PG2_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B2|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B2|P _PG2_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B2|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B2|RB _PG2_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B12|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|B12|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|B12|RB _PG2_12|_AND_G|B12|MID_SHUNT _PG2_12|_AND_G|B3  2.1704737578552e-12
B_PG2_12|_AND_G|Q2|1 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q2|P _PG2_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q2|RB _PG2_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|Q1|1 _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q1|P _PG2_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q1|RB _PG2_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_SPL_G1|I_D1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|I_D1|MID  2e-12
I_PG3_12|_SPL_G1|I_D1|B 0 _PG3_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_D2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|I_D2|MID  2e-12
I_PG3_12|_SPL_G1|I_D2|B 0 _PG3_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_12|_SPL_G1|I_Q1|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|I_Q1|MID  2e-12
I_PG3_12|_SPL_G1|I_Q1|B 0 _PG3_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_Q2|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|I_Q2|MID  2e-12
I_PG3_12|_SPL_G1|I_Q2|B 0 _PG3_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_12|_SPL_G1|1|1 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|1|P _PG3_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|1|RB _PG3_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|2|1 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|2|P _PG3_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|2|RB _PG3_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|A|1 _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|A|P _PG3_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|A|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|A|RB _PG3_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|B|1 _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|B|P _PG3_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|B|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|B|RB _PG3_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_PG|I_A1|B _PG3_12|_PG|A1 _PG3_12|_PG|I_A1|MID  2e-12
I_PG3_12|_PG|I_A1|B 0 _PG3_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_B1|B _PG3_12|_PG|B1 _PG3_12|_PG|I_B1|MID  2e-12
I_PG3_12|_PG|I_B1|B 0 _PG3_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q3|B _PG3_12|_PG|Q3 _PG3_12|_PG|I_Q3|MID  2e-12
I_PG3_12|_PG|I_Q3|B 0 _PG3_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_PG|I_Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|I_Q2|MID  2e-12
I_PG3_12|_PG|I_Q2|B 0 _PG3_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|I_Q1|MID  2e-12
I_PG3_12|_PG|I_Q1|B 0 _PG3_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_PG|A1|1 _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A1|P _PG3_12|_PG|A1|MID_SERIES 0  2e-13
R_PG3_12|_PG|A1|B _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A1|RB _PG3_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A2|1 _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A2|P _PG3_12|_PG|A2|MID_SERIES 0  2e-13
R_PG3_12|_PG|A2|B _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A2|RB _PG3_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A12|1 _PG3_12|_PG|A2 _PG3_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|A12|B _PG3_12|_PG|A2 _PG3_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|A12|RB _PG3_12|_PG|A12|MID_SHUNT _PG3_12|_PG|A3  2.1704737578552e-12
B_PG3_12|_PG|B1|1 _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B1|P _PG3_12|_PG|B1|MID_SERIES 0  2e-13
R_PG3_12|_PG|B1|B _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B1|RB _PG3_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B2|1 _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B2|P _PG3_12|_PG|B2|MID_SERIES 0  2e-13
R_PG3_12|_PG|B2|B _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B2|RB _PG3_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B12|1 _PG3_12|_PG|B2 _PG3_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|B12|B _PG3_12|_PG|B2 _PG3_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|B12|RB _PG3_12|_PG|B12|MID_SHUNT _PG3_12|_PG|B3  2.1704737578552e-12
B_PG3_12|_PG|Q2|1 _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q2|P _PG3_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q2|RB _PG3_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|Q1|1 _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q1|P _PG3_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q1|RB _PG3_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_GG|I_A1|B _PG3_12|_GG|A1 _PG3_12|_GG|I_A1|MID  2e-12
I_PG3_12|_GG|I_A1|B 0 _PG3_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_B1|B _PG3_12|_GG|B1 _PG3_12|_GG|I_B1|MID  2e-12
I_PG3_12|_GG|I_B1|B 0 _PG3_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q3|B _PG3_12|_GG|Q3 _PG3_12|_GG|I_Q3|MID  2e-12
I_PG3_12|_GG|I_Q3|B 0 _PG3_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_GG|I_Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|I_Q2|MID  2e-12
I_PG3_12|_GG|I_Q2|B 0 _PG3_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|I_Q1|MID  2e-12
I_PG3_12|_GG|I_Q1|B 0 _PG3_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_GG|A1|1 _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A1|P _PG3_12|_GG|A1|MID_SERIES 0  2e-13
R_PG3_12|_GG|A1|B _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A1|RB _PG3_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A2|1 _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A2|P _PG3_12|_GG|A2|MID_SERIES 0  2e-13
R_PG3_12|_GG|A2|B _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A2|RB _PG3_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A12|1 _PG3_12|_GG|A2 _PG3_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|A12|B _PG3_12|_GG|A2 _PG3_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|A12|RB _PG3_12|_GG|A12|MID_SHUNT _PG3_12|_GG|A3  2.1704737578552e-12
B_PG3_12|_GG|B1|1 _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B1|P _PG3_12|_GG|B1|MID_SERIES 0  2e-13
R_PG3_12|_GG|B1|B _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B1|RB _PG3_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B2|1 _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B2|P _PG3_12|_GG|B2|MID_SERIES 0  2e-13
R_PG3_12|_GG|B2|B _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B2|RB _PG3_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B12|1 _PG3_12|_GG|B2 _PG3_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|B12|B _PG3_12|_GG|B2 _PG3_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|B12|RB _PG3_12|_GG|B12|MID_SHUNT _PG3_12|_GG|B3  2.1704737578552e-12
B_PG3_12|_GG|Q2|1 _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q2|P _PG3_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q2|RB _PG3_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|Q1|1 _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q1|P _PG3_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q1|RB _PG3_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_PG|I_1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|I_1|MID  2e-12
I_PG3_12|_DFF_PG|I_1|B 0 _PG3_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|I_3|MID  2e-12
I_PG3_12|_DFF_PG|I_3|B 0 _PG3_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_PG|I_T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|I_T|MID  2e-12
I_PG3_12|_DFF_PG|I_T|B 0 _PG3_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|I_6|MID  2e-12
I_PG3_12|_DFF_PG|I_6|B 0 _PG3_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_PG|1|1 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|1|P _PG3_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|1|RB _PG3_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|23|1 _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|23|B _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|23|RB _PG3_12|_DFF_PG|23|MID_SHUNT _PG3_12|_DFF_PG|A3  2.1704737578552e-12
B_PG3_12|_DFF_PG|3|1 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|3|P _PG3_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|3|RB _PG3_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|4|1 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|4|P _PG3_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|4|B _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|4|RB _PG3_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|T|1 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|T|P _PG3_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|T|RB _PG3_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|45|1 _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|45|B _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|45|RB _PG3_12|_DFF_PG|45|MID_SHUNT _PG3_12|_DFF_PG|A4  2.1704737578552e-12
B_PG3_12|_DFF_PG|6|1 _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|6|P _PG3_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|6|RB _PG3_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_GG|I_1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|I_1|MID  2e-12
I_PG3_12|_DFF_GG|I_1|B 0 _PG3_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|I_3|MID  2e-12
I_PG3_12|_DFF_GG|I_3|B 0 _PG3_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_GG|I_T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|I_T|MID  2e-12
I_PG3_12|_DFF_GG|I_T|B 0 _PG3_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|I_6|MID  2e-12
I_PG3_12|_DFF_GG|I_6|B 0 _PG3_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_GG|1|1 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|1|P _PG3_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|1|RB _PG3_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|23|1 _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|23|B _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|23|RB _PG3_12|_DFF_GG|23|MID_SHUNT _PG3_12|_DFF_GG|A3  2.1704737578552e-12
B_PG3_12|_DFF_GG|3|1 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|3|P _PG3_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|3|RB _PG3_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|4|1 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|4|P _PG3_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|4|B _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|4|RB _PG3_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|T|1 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|T|P _PG3_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|T|RB _PG3_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|45|1 _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|45|B _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|45|RB _PG3_12|_DFF_GG|45|MID_SHUNT _PG3_12|_DFF_GG|A4  2.1704737578552e-12
B_PG3_12|_DFF_GG|6|1 _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|6|P _PG3_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|6|RB _PG3_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_G|I_A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|I_A1|MID  2e-12
I_PG3_12|_AND_G|I_A1|B 0 _PG3_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|I_B1|MID  2e-12
I_PG3_12|_AND_G|I_B1|B 0 _PG3_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q3|B _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|I_Q3|MID  2e-12
I_PG3_12|_AND_G|I_Q3|B 0 _PG3_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_G|I_Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|I_Q2|MID  2e-12
I_PG3_12|_AND_G|I_Q2|B 0 _PG3_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|I_Q1|MID  2e-12
I_PG3_12|_AND_G|I_Q1|B 0 _PG3_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_G|A1|1 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A1|P _PG3_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A1|RB _PG3_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A2|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A2|P _PG3_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A2|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A2|RB _PG3_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A12|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|A12|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|A12|RB _PG3_12|_AND_G|A12|MID_SHUNT _PG3_12|_AND_G|A3  2.1704737578552e-12
B_PG3_12|_AND_G|B1|1 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B1|P _PG3_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B1|RB _PG3_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B2|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B2|P _PG3_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B2|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B2|RB _PG3_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B12|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|B12|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|B12|RB _PG3_12|_AND_G|B12|MID_SHUNT _PG3_12|_AND_G|B3  2.1704737578552e-12
B_PG3_12|_AND_G|Q2|1 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q2|P _PG3_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q2|RB _PG3_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|Q1|1 _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q1|P _PG3_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q1|RB _PG3_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_S0
.print DEVI R_S1
.print DEVI R_S2
.print DEVI R_S3
.print DEVI R_S4
.print DEVI IA0|A
.print DEVI IB0|B
.print DEVI IA1|C
.print DEVI IB1|D
.print DEVI IA2|E
.print DEVI IB2|F
.print DEVI IA3|G
.print DEVI IB3|H
.print DEVI IT00|T
.print DEVI IT01|T
.print DEVI IT02|T
.print DEVI IT03|T
.print DEVI LSPL_IG0_0|1
.print DEVI LSPL_IG0_0|2
.print DEVI LSPL_IG0_0|3
.print DEVI LSPL_IG0_0|4
.print DEVI LSPL_IG0_0|5
.print DEVI LSPL_IG0_0|6
.print DEVI LSPL_IG0_0|7
.print DEVI LSPL_IP1_0|1
.print DEVI LSPL_IP1_0|2
.print DEVI LSPL_IP1_0|3
.print DEVI LSPL_IP1_0|4
.print DEVI LSPL_IP1_0|5
.print DEVI LSPL_IP1_0|6
.print DEVI LSPL_IP1_0|7
.print DEVI LSPL_IG2_0|1
.print DEVI LSPL_IG2_0|2
.print DEVI LSPL_IG2_0|3
.print DEVI LSPL_IG2_0|4
.print DEVI LSPL_IG2_0|5
.print DEVI LSPL_IG2_0|6
.print DEVI LSPL_IG2_0|7
.print DEVI LSPL_IP3_0|1
.print DEVI LSPL_IP3_0|2
.print DEVI LSPL_IP3_0|3
.print DEVI LSPL_IP3_0|4
.print DEVI LSPL_IP3_0|5
.print DEVI LSPL_IP3_0|6
.print DEVI LSPL_IP3_0|7
.print DEVI IT04|T
.print DEVI IT05|T
.print DEVI IT06|T
.print DEVI IT07|T
.print DEVI ID01|T
.print DEVI L_DFF_IP1_01|1
.print DEVI L_DFF_IP1_01|2
.print DEVI L_DFF_IP1_01|3
.print DEVI L_DFF_IP1_01|T
.print DEVI L_DFF_IP1_01|4
.print DEVI L_DFF_IP1_01|5
.print DEVI L_DFF_IP1_01|6
.print DEVI ID02|T
.print DEVI L_DFF_IP2_01|1
.print DEVI L_DFF_IP2_01|2
.print DEVI L_DFF_IP2_01|3
.print DEVI L_DFF_IP2_01|T
.print DEVI L_DFF_IP2_01|4
.print DEVI L_DFF_IP2_01|5
.print DEVI L_DFF_IP2_01|6
.print DEVI ID03|T
.print DEVI L_DFF_IP3_01|1
.print DEVI L_DFF_IP3_01|2
.print DEVI L_DFF_IP3_01|3
.print DEVI L_DFF_IP3_01|T
.print DEVI L_DFF_IP3_01|4
.print DEVI L_DFF_IP3_01|5
.print DEVI L_DFF_IP3_01|6
.print DEVI IT08|T
.print DEVI IT09|T
.print DEVI L_PG1_12|1
.print DEVI L_PG1_12|2
.print DEVI L_PG1_12|3
.print DEVI L_PG1_12|T
.print DEVI L_PG1_12|4
.print DEVI L_PG1_12|5
.print DEVI L_PG1_12|6
.print DEVI IT10|T
.print DEVI IT11|T
.print DEVI ID11|T
.print DEVI L_DFF_IP1_12|1
.print DEVI L_DFF_IP1_12|2
.print DEVI L_DFF_IP1_12|3
.print DEVI L_DFF_IP1_12|T
.print DEVI L_DFF_IP1_12|4
.print DEVI L_DFF_IP1_12|5
.print DEVI L_DFF_IP1_12|6
.print DEVI ID12|T
.print DEVI L_DFF_IP2_12|1
.print DEVI L_DFF_IP2_12|2
.print DEVI L_DFF_IP2_12|3
.print DEVI L_DFF_IP2_12|T
.print DEVI L_DFF_IP2_12|4
.print DEVI L_DFF_IP2_12|5
.print DEVI L_DFF_IP2_12|6
.print DEVI ID13|T
.print DEVI L_DFF_IP3_12|1
.print DEVI L_DFF_IP3_12|2
.print DEVI L_DFF_IP3_12|3
.print DEVI L_DFF_IP3_12|T
.print DEVI L_DFF_IP3_12|4
.print DEVI L_DFF_IP3_12|5
.print DEVI L_DFF_IP3_12|6
.print DEVI IT12|T
.print DEVI L_S0|1
.print DEVI L_S0|2
.print DEVI L_S0|3
.print DEVI L_S0|T
.print DEVI L_S0|4
.print DEVI L_S0|5
.print DEVI L_S0|6
.print DEVI IT13|T
.print DEVI L_S1|A1
.print DEVI L_S1|A2
.print DEVI L_S1|A3
.print DEVI L_S1|B1
.print DEVI L_S1|B2
.print DEVI L_S1|B3
.print DEVI L_S1|T1
.print DEVI L_S1|T2
.print DEVI L_S1|Q2
.print DEVI L_S1|Q1
.print DEVI IT14|T
.print DEVI L_S2|A1
.print DEVI L_S2|A2
.print DEVI L_S2|A3
.print DEVI L_S2|B1
.print DEVI L_S2|B2
.print DEVI L_S2|B3
.print DEVI L_S2|T1
.print DEVI L_S2|T2
.print DEVI L_S2|Q2
.print DEVI L_S2|Q1
.print DEVI IT15|T
.print DEVI L_S3|A1
.print DEVI L_S3|A2
.print DEVI L_S3|A3
.print DEVI L_S3|B1
.print DEVI L_S3|B2
.print DEVI L_S3|B3
.print DEVI L_S3|T1
.print DEVI L_S3|T2
.print DEVI L_S3|Q2
.print DEVI L_S3|Q1
.print DEVI IT16|T
.print DEVI L_S4|1
.print DEVI L_S4|2
.print DEVI L_S4|3
.print DEVI L_S4|T
.print DEVI L_S4|4
.print DEVI L_S4|5
.print DEVI L_S4|6
.print V I1|A1
.print V T01
.print V B0_TX
.print V _PG3_12|PG_SYNC
.print V _DFF_IP1_12|T1
.print V _S3|T2
.print V _S3|B3
.print V _S0|Q1
.print V _S0|T2
.print V T12
.print V _PG1_01|GG
.print V A2_RX
.print V _DFF_IP3_01|Q1
.print V _PTL_IP3_0|A_PTL
.print V A3_TX
.print V SPL_IP1_0|D1
.print V G0_2
.print V P0_1
.print V _PTL_B0|A_PTL
.print V T16
.print V _S2|A3
.print V P3_1
.print V B2_TX
.print V _PTL_G1_2|A_PTL_RX
.print V _PTL_IP2_1|A_PTL
.print V _DFF_IP3_12|A1
.print V SPL_IP1_0|QA1
.print V IP2_0_RX
.print V IP3_0_OUT
.print V _PG3_01|G1_COPY_1
.print V _PG3_12|G1_COPY_2
.print V B0_RX
.print V _PTL_G0_2|A_PTL
.print V _DFF_IP3_01|T2
.print V _PG1_12|T1
.print V B1_RX
.print V _PG2_12|G1_COPY_2
.print V G1_1_RX
.print V T15
.print V IG2_0_RX
.print V IG0_0_RX
.print V I0|B1_SYNC
.print V I0|A2
.print V _PG1_01|PG
.print V _PTL_G0_1|A_PTL
.print V _S2|T2
.print V _S3|B1
.print V _PTL_P3_1|A_PTL
.print V _PG3_12|GG
.print V _DFF_IP2_12|Q1
.print V S2
.print V _DFF_IP3_12|T2
.print V IP3_2_OUT_RX
.print V _PTL_IP1_2|A_PTL
.print V A1_RX
.print V _DFF_IP2_01|A4
.print V _PTL_B2|A_PTL
.print V _PTL_G1_1|A_PTL
.print V D03
.print V _DFF_IP2_01|T1
.print V _S0|A2
.print V I2|A2
.print V _PTL_A3|A_PTL
.print V _PTL_IP2_0|A_PTL
.print V SPL_IP3_0|D2
.print V IP2_0_TO3
.print V _PTL_G3_2|A_PTL
.print V _PG1_01|PG_SYNC
.print V B1_TX
.print V _DFF_IP3_01|T1
.print V IP2_1_OUT
.print V _DFF_IP1_12|A2
.print V T14
.print V _PTL_IP3_2|A_PTL_RX
.print V IG1_0
.print V P0_2
.print V _S4|A2
.print V _PTL_G2_2|A_PTL
.print V SPL_IG0_0|QB1
.print V P3_1_RX
.print V I3|B2
.print V G3_2_RX
.print V _DFF_IP3_01|A1
.print V A0_TX
.print V I3|B1_SYNC
.print V _PG2_12|PG
.print V SPL_IG2_0|JCT
.print V _PTL_IP1_0|A_PTL
.print V G3_1
.print V T05
.print V T13
.print V _S4|T1
.print V _PG3_01|PG_SYNC
.print V _S1|ABTQ
.print V _PG3_12|GG_SYNC
.print V IG0_0_TO1
.print V SPL_IP1_0|JCT
.print V G1_1
.print V _PTL_A0|A_PTL
.print V _S3|ABTQ
.print V _DFF_IP1_01|T1
.print V _DFF_IP2_12|A1
.print V _S0|A3
.print V _PTL_G2_1|A_PTL
.print V _S3|A3
.print V _S4|T2
.print V _PTL_G2_2|A_PTL_RX
.print V _PTL_IP0_0|A_PTL
.print V _DFF_IP3_01|A4
.print V _S2|B3
.print V _S4|Q1
.print V I0|B2
.print V _S2|ABTQ
.print V _S0|T1
.print V I1|B2
.print V P0_1_RX
.print V IP2_1_OUT_RX
.print V A2_TX
.print V D02
.print V D01
.print V I3|A2
.print V _DFF_IP3_12|A2
.print V _S3|B2
.print V _S2|Q1
.print V IG2_0_TO2
.print V G2_2
.print V SPL_G1_1|QTMP
.print V _DFF_IP1_01|T2
.print V T09
.print V _DFF_IP3_12|Q1
.print V _PTL_IG1_0|A_PTL
.print V _DFF_IP2_01|Q1
.print V I3|A1_SYNC
.print V IP3_0_RX
.print V _S3|Q1
.print V SPL_IG2_0|QA1
.print V _S1|A2
.print V _PG3_01|P1_COPY_2
.print V P2_1
.print V _DFF_IP2_12|A2
.print V _DFF_IP1_12|Q1
.print V SPL_IG2_0|QB1
.print V IP1_1_OUT
.print V S1
.print V I0|A1
.print V _S3|A1
.print V SPL_IG0_0|QA1
.print V IP2_2_OUT_RX
.print V _S1|T2
.print V D13
.print V SPL_IP1_0|QB1
.print V T03
.print V SPL_IG2_0|D1
.print V G1_2_RX
.print V _S2|AB
.print V T08
.print V SPL_IG0_0|JCT
.print V _PG1_01|G1_COPY_2
.print V IP2_0_TO2
.print V IP3_0_TO1
.print V _S2|A2
.print V SPL_IP3_0|QA1
.print V I0|B1
.print V _PG3_01|P0_SYNC
.print V IP3_0
.print V _PTL_IP3_1|A_PTL
.print V _PG1_12|A3
.print V IP1_0
.print V IP3_1_OUT_RX
.print V IP1_0_RX
.print V SPL_IG0_0|D1
.print V SPL_IG2_0|D2
.print V _PTL_IG0_0|A_PTL
.print V _PG1_12|Q1
.print V T06
.print V _PTL_P0_1|A_PTL
.print V _PG1_01|G1_COPY_1
.print V IP2_0_OUT
.print V IP1_2_OUT_RX
.print V _DFF_IP2_12|A4
.print V I1|A2
.print V _PG1_12|T2
.print V _PTL_IP2_2|A_PTL
.print V _S2|A1
.print V I3|B1
.print V _PTL_P0_2|A_PTL
.print V _PTL_IP1_1|A_PTL
.print V _PTL_IP3_2|A_PTL
.print V SPL_IP3_0|QB1
.print V SPL_IP2_0|QTMP
.print V _DFF_IP3_12|A3
.print V IP1_0_OUT
.print V _PG2_12|PG_SYNC
.print V _DFF_IP1_01|A4
.print V _PG1_12|A2
.print V SPL_IP3_0|D1
.print V G1_2
.print V _DFF_IP1_01|Q1
.print V IG3_0_RX
.print V G0_1
.print V _DFF_IP1_01|A3
.print V _PG3_01|GG_SYNC
.print V _PG3_01|P1_COPY_1
.print V _S0|A4
.print V I2|A1
.print V _PG1_12|A4
.print V _PTL_IP2_2|A_PTL_RX
.print V _PG2_12|G1_COPY_1
.print V _PTL_P0_2|A_PTL_RX
.print V _S4|A1
.print V G0_1_RX
.print V D11
.print V I2|B1_SYNC
.print V G1_1_TO2
.print V _DFF_IP1_12|A3
.print V _PTL_IG3_0|A_PTL
.print V _PG3_01|P1_SYNC
.print V _DFF_IP2_01|A2
.print V _S3|T1
.print V IG0_0
.print V IG3_0
.print V B3_TX
.print V _S1|AB
.print V IG1_0_RX
.print V I2|B1
.print V _PTL_G3_2|A_PTL_RX
.print V SPL_IG0_0|D2
.print V _S1|B2
.print V IG2_0
.print V T10
.print V _DFF_IP3_01|A2
.print V _S1|Q1
.print V IP0_0_RX
.print V S4
.print V T02
.print V B3_RX
.print V S0
.print V G3_2
.print V SPL_IP1_0|D2
.print V _PG2_12|GG
.print V SPL_IP3_0|JCT
.print V _PG3_12|PG
.print V _PG1_12|A1
.print V _S1|B1
.print V D12
.print V _PG1_01|GG_SYNC
.print V G2_1_RX
.print V _DFF_IP3_12|T1
.print V _PG3_12|G1_COPY_1
.print V _PG3_01|GG
.print V _S1|A3
.print V I0|A1_SYNC
.print V B2_RX
.print V _S3|AB
.print V _DFF_IP1_01|A1
.print V _S4|A4
.print V _S3|A2
.print V _DFF_IP2_12|T1
.print V S3
.print V G2_2_RX
.print V _S1|T1
.print V IP3_2_OUT
.print V _S4|A3
.print V G3_1_RX
.print V _PTL_A2|A_PTL
.print V _S1|B3
.print V I1|B1
.print V IG0_0_TO0
.print V _S2|T1
.print V T04
.print V T00
.print V IP2_2_OUT
.print V _DFF_IP1_12|T2
.print V _PG3_01|PG
.print V _PTL_B1|A_PTL
.print V A0_RX
.print V _PTL_G3_1|A_PTL
.print V _DFF_IP1_12|A1
.print V IG2_0_TO3
.print V _PTL_IG2_0|A_PTL
.print V T07
.print V _PG3_01|G1_COPY_2
.print V IP2_0
.print V _DFF_IP2_01|A3
.print V A1_TX
.print V I1|A1_SYNC
.print V _DFF_IP2_01|T2
.print V _PTL_G1_2|A_PTL
.print V _DFF_IP3_01|A3
.print V I3|A1
.print V IP0_0
.print V _PTL_A1|A_PTL
.print V IP3_1_OUT
.print V _PTL_P2_1|A_PTL
.print V I1|B1_SYNC
.print V IP1_1_OUT_RX
.print V G1_1_TO1
.print V _DFF_IP2_12|A3
.print V G0_2_RX
.print V T11
.print V G2_1
.print V _PTL_IP1_2|A_PTL_RX
.print V IP1_2_OUT
.print V _DFF_IP2_12|T2
.print V P0_2_RX
.print V G1_1_TO3
.print V _DFF_IP1_01|A2
.print V _S1|A1
.print V _DFF_IP2_01|A1
.print V _DFF_IP1_12|A4
.print V A3_RX
.print V _PTL_B3|A_PTL
.print V _S2|B1
.print V _S0|A1
.print V _PG2_12|GG_SYNC
.print V _DFF_IP3_12|A4
.print V I2|B2
.print V _S2|B2
.print V IP1_0_TO1
.print V _PTL_G0_2|A_PTL_RX
.print V I2|A1_SYNC
.print V P2_1_RX
