*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM IU=1.25e-05
.PARAM VU=0.0006857
.PARAM LU=2.632e-12
.PARAM JCRIT=5e-05
.PARAM OFFSET1=5e-11
.PARAM TCLOCK=4e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT_ADJ JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 4E-9
LINPUT CLK0 CLK  PHI0/(4*IC*IC0)
LSUM SUM0 SUM1  PHI0/(4*IC*IC0)
RSUM SUM 0  1
LCARRY CARRY0 CARRY1  PHI0/(4*IC*IC0)
RCARRY CARRY 0  1
RCBAR CBAR 0  1
IDATA|H 0 A  PWL(0 0 -5.3e-11 0 -5e-11 0 -4.7e-11 0 4.7e-11 0 5e-11 0 5.3e-11 0 1.47e-10 0 1.5e-10 0 1.53e-10 0 2.47e-10 0 2.5e-10 0 2.53e-10 0 3.47e-10 0 3.5e-10 0 3.53e-10 0 4.47e-10 0 4.5e-10 0 4.53e-10 0 5.47e-10 0 5.5e-10 0 5.53e-10 0 6.47e-10 0 6.5e-10 0 6.53e-10 0 7.47e-10 0 7.5e-10 0.0007 7.53e-10 0 8.47e-10 0 8.5e-10 0 8.53e-10 0 9.47e-10 0 9.5e-10 0 9.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.147e-09 0 1.15e-09 0 1.153e-09 0 1.247e-09 0 1.25e-09 0 1.253e-09 0 1.347e-09 0 1.35e-09 0.0007 1.353e-09 0 1.447e-09 0 1.45e-09 0 1.453e-09 0 1.547e-09 0 1.55e-09 0 1.553e-09 0 1.647e-09 0 1.65e-09 0 1.653e-09 0 1.747e-09 0 1.75e-09 0 1.753e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 1.947e-09 0 1.95e-09 0.0007 1.953e-09 0 2.047e-09 0 2.05e-09 0 2.053e-09 0 2.147e-09 0 2.15e-09 0.0007 2.153e-09 0 2.247e-09 0 2.25e-09 0 2.253e-09 0 2.347e-09 0 2.35e-09 0.0007 2.353e-09 0 2.447e-09 0 2.45e-09 0 2.453e-09 0 2.547e-09 0 2.55e-09 0.0007 2.553e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.747e-09 0 2.75e-09 0 2.753e-09 0 2.847e-09 0 2.85e-09 0 2.853e-09 0 2.947e-09 0 2.95e-09 0.0007 2.953e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.147e-09 0 3.15e-09 0.0007 3.153e-09 0 3.247e-09 0 3.25e-09 0 3.253e-09 0 3.347e-09 0 3.35e-09 0 3.353e-09 0 3.447e-09 0 3.45e-09 0.0014 3.453e-09 0 3.547e-09 0 3.55e-09 0 3.553e-09 0 3.647e-09 0 3.65e-09 0 3.653e-09 0 3.747e-09 0 3.75e-09 0 3.753e-09 0 3.847e-09 0 3.85e-09 0 3.853e-09 0 3.947e-09 0 3.95e-09 0 3.953e-09 0 4.047e-09 0 4.05e-09 0 4.053e-09 0 4.147e-09 0 4.15e-09 0 4.153e-09 0 4.247e-09 0 4.25e-09 0 4.253e-09 0 4.347e-09 0 4.35e-09 0 4.353e-09 0 4.447e-09 0 4.45e-09 0 4.453e-09 0 4.547e-09 0 4.55e-09 0 4.553e-09 0 4.647e-09 0 4.65e-09 0 4.653e-09 0 4.747e-09 0 4.75e-09 0 4.753e-09 0 4.847e-09 0 4.85e-09 0 4.853e-09 0 4.947e-09 0 4.95e-09 0 4.953e-09 0 5.047e-09 0 5.05e-09 0 5.053e-09 0 5.147e-09 0 5.15e-09 0 5.153e-09 0 5.247e-09 0 5.25e-09 0 5.253e-09 0 5.347e-09 0 5.35e-09 0 5.353e-09 0 5.447e-09 0 5.45e-09 0 5.453e-09 0 5.547e-09 0 5.55e-09 0 5.553e-09 0 5.647e-09 0 5.65e-09 0 5.653e-09 0 5.747e-09 0 5.75e-09 0 5.753e-09 0 5.847e-09 0 5.85e-09 0 5.853e-09 0 5.947e-09 0 5.95e-09 0 5.953e-09 0 6.047e-09 0 6.05e-09 0 6.053e-09 0 6.147e-09 0 6.15e-09 0 6.153e-09 0 6.247e-09 0 6.25e-09 0 6.253e-09 0 6.347e-09 0 6.35e-09 0 6.353e-09 0 6.447e-09 0 6.45e-09 0 6.453e-09 0 6.547e-09 0 6.55e-09 0 6.553e-09 0 6.647e-09 0 6.65e-09 0 6.653e-09 0 6.747e-09 0 6.75e-09 0 6.753e-09 0 6.847e-09 0 6.85e-09 0 6.853e-09 0 6.947e-09 0 6.95e-09 0 6.953e-09 0 7.047e-09 0 7.05e-09 0 7.053e-09 0 7.147e-09 0 7.15e-09 0 7.153e-09 0 7.247e-09 0 7.25e-09 0 7.253e-09 0 7.347e-09 0 7.35e-09 0 7.353e-09 0 7.447e-09 0 7.45e-09 0 7.453e-09 0 7.547e-09 0 7.55e-09 0 7.553e-09 0 7.647e-09 0 7.65e-09 0 7.653e-09 0 7.747e-09 0 7.75e-09 0 7.753e-09 0 7.847e-09 0 7.85e-09 0 7.853e-09 0 7.947e-09 0 7.95e-09 0 7.953e-09 0 8.047e-09 0 8.05e-09 0 8.053e-09 0 8.147e-09 0 8.15e-09 0 8.153e-09 0 8.247e-09 0 8.25e-09 0 8.253e-09 0 8.347e-09 0 8.35e-09 0 8.353e-09 0 8.447e-09 0 8.45e-09 0 8.453e-09 0 8.547e-09 0 8.55e-09 0 8.553e-09 0 8.647e-09 0 8.65e-09 0 8.653e-09 0 8.747e-09 0 8.75e-09 0 8.753e-09 0 8.847e-09 0 8.85e-09 0 8.853e-09 0 8.947e-09 0 8.95e-09 0 8.953e-09 0 9.047e-09 0 9.05e-09 0 9.053e-09 0 9.147e-09 0 9.15e-09 0 9.153e-09 0 9.247e-09 0 9.25e-09 0 9.253e-09 0 9.347e-09 0 9.35e-09 0 9.353e-09 0 9.447e-09 0 9.45e-09 0 9.453e-09 0 9.547e-09 0 9.55e-09 0 9.553e-09 0 9.647e-09 0 9.65e-09 0 9.653e-09 0 9.747e-09 0 9.75e-09 0 9.753e-09 0 9.847e-09 0 9.85e-09 0 9.853e-09 0 9.947e-09 0 9.95e-09 0 9.953e-09 0 1.0047e-08 0 1.005e-08 0 1.0053e-08 0 1.0147e-08 0 1.015e-08 0 1.0153e-08 0 1.0247e-08 0 1.025e-08 0 1.0253e-08 0 1.0347e-08 0 1.035e-08 0 1.0353e-08 0 1.0447e-08 0 1.045e-08 0 1.0453e-08 0 1.0547e-08 0 1.055e-08 0 1.0553e-08 0 1.0647e-08 0 1.065e-08 0 1.0653e-08 0 1.0747e-08 0 1.075e-08 0 1.0753e-08 0 1.0847e-08 0 1.085e-08 0 1.0853e-08 0 1.0947e-08 0 1.095e-08 0 1.0953e-08 0 1.1047e-08 0 1.105e-08 0 1.1053e-08 0 1.1147e-08 0 1.115e-08 0 1.1153e-08 0 1.1247e-08 0 1.125e-08 0 1.1253e-08 0 1.1347e-08 0 1.135e-08 0 1.1353e-08 0 1.1447e-08 0 1.145e-08 0 1.1453e-08 0 1.1547e-08 0 1.155e-08 0 1.1553e-08 0 1.1647e-08 0 1.165e-08 0 1.1653e-08 0 1.1747e-08 0 1.175e-08 0 1.1753e-08 0 1.1847e-08 0 1.185e-08 0 1.1853e-08 0 1.1947e-08 0 1.195e-08 0 1.1953e-08 0 1.2047e-08 0 1.205e-08 0 1.2053e-08 0 1.2147e-08 0 1.215e-08 0 1.2153e-08 0 1.2247e-08 0 1.225e-08 0 1.2253e-08 0 1.2347e-08 0 1.235e-08 0 1.2353e-08 0 1.2447e-08 0 1.245e-08 0 1.2453e-08 0 1.2547e-08 0 1.255e-08 0 1.2553e-08 0 1.2647e-08 0 1.265e-08 0 1.2653e-08 0 1.2747e-08 0 1.275e-08 0 1.2753e-08 0)
IT1|T 0 CLK0  PWL(0 0 4.7e-11 0 5e-11 0.000231 5.3e-11 0 4.47e-10 0 4.5e-10 0.000231 4.53e-10 0 8.47e-10 0 8.5e-10 0.000231 8.53e-10 0 1.247e-09 0 1.25e-09 0.000231 1.253e-09 0 1.647e-09 0 1.65e-09 0.000231 1.653e-09 0 2.047e-09 0 2.05e-09 0.000231 2.053e-09 0 2.447e-09 0 2.45e-09 0.000231 2.453e-09 0 2.847e-09 0 2.85e-09 0.000231 2.853e-09 0 3.247e-09 0 3.25e-09 0.000231 3.253e-09 0 3.647e-09 0 3.65e-09 0.000231 3.653e-09 0 4.047e-09 0 4.05e-09 0.000231 4.053e-09 0 4.447e-09 0 4.45e-09 0.000231 4.453e-09 0 4.847e-09 0 4.85e-09 0.000231 4.853e-09 0 5.247e-09 0 5.25e-09 0.000231 5.253e-09 0 5.647e-09 0 5.65e-09 0.000231 5.653e-09 0 6.047e-09 0 6.05e-09 0.000231 6.053e-09 0 6.447e-09 0 6.45e-09 0.000231 6.453e-09 0 6.847e-09 0 6.85e-09 0.000231 6.853e-09 0 7.247e-09 0 7.25e-09 0.000231 7.253e-09 0 7.647e-09 0 7.65e-09 0.000231 7.653e-09 0 8.047e-09 0 8.05e-09 0.000231 8.053e-09 0 8.447e-09 0 8.45e-09 0.000231 8.453e-09 0 8.847e-09 0 8.85e-09 0.000231 8.853e-09 0 9.247e-09 0 9.25e-09 0.000231 9.253e-09 0 9.647e-09 0 9.65e-09 0.000231 9.653e-09 0 1.0047e-08 0 1.005e-08 0.000231 1.0053e-08 0 1.0447e-08 0 1.045e-08 0.000231 1.0453e-08 0 1.0847e-08 0 1.085e-08 0.000231 1.0853e-08 0 1.1247e-08 0 1.125e-08 0.000231 1.1253e-08 0 1.1647e-08 0 1.165e-08 0.000231 1.1653e-08 0 1.2047e-08 0 1.205e-08 0.000231 1.2053e-08 0 1.2447e-08 0 1.245e-08 0.000231 1.2453e-08 0 1.2847e-08 0 1.285e-08 0.000231 1.2853e-08 0 1.3247e-08 0 1.325e-08 0.000231 1.3253e-08 0 1.3647e-08 0 1.365e-08 0.000231 1.3653e-08 0 1.4047e-08 0 1.405e-08 0.000231 1.4053e-08 0 1.4447e-08 0 1.445e-08 0.000231 1.4453e-08 0 1.4847e-08 0 1.485e-08 0.000231 1.4853e-08 0 1.5247e-08 0 1.525e-08 0.000231 1.5253e-08 0 1.5647e-08 0 1.565e-08 0.000231 1.5653e-08 0 1.6047e-08 0 1.605e-08 0.000231 1.6053e-08 0 1.6447e-08 0 1.645e-08 0.000231 1.6453e-08 0 1.6847e-08 0 1.685e-08 0.000231 1.6853e-08 0 1.7247e-08 0 1.725e-08 0.000231 1.7253e-08 0 1.7647e-08 0 1.765e-08 0.000231 1.7653e-08 0 1.8047e-08 0 1.805e-08 0.000231 1.8053e-08 0 1.8447e-08 0 1.845e-08 0.000231 1.8453e-08 0 1.8847e-08 0 1.885e-08 0.000231 1.8853e-08 0 1.9247e-08 0 1.925e-08 0.000231 1.9253e-08 0 1.9647e-08 0 1.965e-08 0.000231 1.9653e-08 0 2.0047e-08 0 2.005e-08 0.000231 2.0053e-08 0 2.0447e-08 0 2.045e-08 0.000231 2.0453e-08 0 2.0847e-08 0 2.085e-08 0.000231 2.0853e-08 0 2.1247e-08 0 2.125e-08 0.000231 2.1253e-08 0 2.1647e-08 0 2.165e-08 0.000231 2.1653e-08 0 2.2047e-08 0 2.205e-08 0.000231 2.2053e-08 0 2.2447e-08 0 2.245e-08 0.000231 2.2453e-08 0 2.2847e-08 0 2.285e-08 0.000231 2.2853e-08 0 2.3247e-08 0 2.325e-08 0.000231 2.3253e-08 0 2.3647e-08 0 2.365e-08 0.000231 2.3653e-08 0 2.4047e-08 0 2.405e-08 0.000231 2.4053e-08 0 2.4447e-08 0 2.445e-08 0.000231 2.4453e-08 0 2.4847e-08 0 2.485e-08 0.000231 2.4853e-08 0 2.5247e-08 0 2.525e-08 0.000231 2.5253e-08 0 2.5647e-08 0 2.565e-08 0.000231 2.5653e-08 0 2.6047e-08 0 2.605e-08 0.000231 2.6053e-08 0 2.6447e-08 0 2.645e-08 0.000231 2.6453e-08 0 2.6847e-08 0 2.685e-08 0.000231 2.6853e-08 0 2.7247e-08 0 2.725e-08 0.000231 2.7253e-08 0 2.7647e-08 0 2.765e-08 0.000231 2.7653e-08 0 2.8047e-08 0 2.805e-08 0.000231 2.8053e-08 0 2.8447e-08 0 2.845e-08 0.000231 2.8453e-08 0 2.8847e-08 0 2.885e-08 0.000231 2.8853e-08 0 2.9247e-08 0 2.925e-08 0.000231 2.9253e-08 0 2.9647e-08 0 2.965e-08 0.000231 2.9653e-08 0 3.0047e-08 0 3.005e-08 0.000231 3.0053e-08 0 3.0447e-08 0 3.045e-08 0.000231 3.0453e-08 0 3.0847e-08 0 3.085e-08 0.000231 3.0853e-08 0 3.1247e-08 0 3.125e-08 0.000231 3.1253e-08 0 3.1647e-08 0 3.165e-08 0.000231 3.1653e-08 0 3.2047e-08 0 3.205e-08 0.000231 3.2053e-08 0 3.2447e-08 0 3.245e-08 0.000231 3.2453e-08 0 3.2847e-08 0 3.285e-08 0.000231 3.2853e-08 0 3.3247e-08 0 3.325e-08 0.000231 3.3253e-08 0 3.3647e-08 0 3.365e-08 0.000231 3.3653e-08 0 3.4047e-08 0 3.405e-08 0.000231 3.4053e-08 0 3.4447e-08 0 3.445e-08 0.000231 3.4453e-08 0 3.4847e-08 0 3.485e-08 0.000231 3.4853e-08 0 3.5247e-08 0 3.525e-08 0.000231 3.5253e-08 0 3.5647e-08 0 3.565e-08 0.000231 3.5653e-08 0 3.6047e-08 0 3.605e-08 0.000231 3.6053e-08 0 3.6447e-08 0 3.645e-08 0.000231 3.6453e-08 0 3.6847e-08 0 3.685e-08 0.000231 3.6853e-08 0 3.7247e-08 0 3.725e-08 0.000231 3.7253e-08 0 3.7647e-08 0 3.765e-08 0.000231 3.7653e-08 0 3.8047e-08 0 3.805e-08 0.000231 3.8053e-08 0 3.8447e-08 0 3.845e-08 0.000231 3.8453e-08 0 3.8847e-08 0 3.885e-08 0.000231 3.8853e-08 0 3.9247e-08 0 3.925e-08 0.000231 3.9253e-08 0 3.9647e-08 0 3.965e-08 0.000231 3.9653e-08 0 4.0047e-08 0 4.005e-08 0.000231 4.0053e-08 0 4.0447e-08 0 4.045e-08 0.000231 4.0453e-08 0 4.0847e-08 0 4.085e-08 0.000231 4.0853e-08 0 4.1247e-08 0 4.125e-08 0.000231 4.1253e-08 0 4.1647e-08 0 4.165e-08 0.000231 4.1653e-08 0 4.2047e-08 0 4.205e-08 0.000231 4.2053e-08 0 4.2447e-08 0 4.245e-08 0.000231 4.2453e-08 0 4.2847e-08 0 4.285e-08 0.000231 4.2853e-08 0 4.3247e-08 0 4.325e-08 0.000231 4.3253e-08 0 4.3647e-08 0 4.365e-08 0.000231 4.3653e-08 0 4.4047e-08 0 4.405e-08 0.000231 4.4053e-08 0 4.4447e-08 0 4.445e-08 0.000231 4.4453e-08 0 4.4847e-08 0 4.485e-08 0.000231 4.4853e-08 0 4.5247e-08 0 4.525e-08 0.000231 4.5253e-08 0 4.5647e-08 0 4.565e-08 0.000231 4.5653e-08 0 4.6047e-08 0 4.605e-08 0.000231 4.6053e-08 0 4.6447e-08 0 4.645e-08 0.000231 4.6453e-08 0 4.6847e-08 0 4.685e-08 0.000231 4.6853e-08 0 4.7247e-08 0 4.725e-08 0.000231 4.7253e-08 0 4.7647e-08 0 4.765e-08 0.000231 4.7653e-08 0 4.8047e-08 0 4.805e-08 0.000231 4.8053e-08 0 4.8447e-08 0 4.845e-08 0.000231 4.8453e-08 0 4.8847e-08 0 4.885e-08 0.000231 4.8853e-08 0 4.9247e-08 0 4.925e-08 0.000231 4.9253e-08 0 4.9647e-08 0 4.965e-08 0.000231 4.9653e-08 0 5.0047e-08 0 5.005e-08 0.000231 5.0053e-08 0 5.0447e-08 0 5.045e-08 0.000231 5.0453e-08 0 5.0847e-08 0 5.085e-08 0.000231 5.0853e-08 0 5.1247e-08 0 5.125e-08 0.000231 5.1253e-08 0 5.1647e-08 0 5.165e-08 0.000231 5.1653e-08 0 5.2047e-08 0 5.205e-08 0.000231 5.2053e-08 0 5.2447e-08 0 5.245e-08 0.000231 5.2453e-08 0 5.2847e-08 0 5.285e-08 0.000231 5.2853e-08 0 5.3247e-08 0 5.325e-08 0.000231 5.3253e-08 0 5.3647e-08 0 5.365e-08 0.000231 5.3653e-08 0 5.4047e-08 0 5.405e-08 0.000231 5.4053e-08 0 5.4447e-08 0 5.445e-08 0.000231 5.4453e-08 0 5.4847e-08 0 5.485e-08 0.000231 5.4853e-08 0 5.5247e-08 0 5.525e-08 0.000231 5.5253e-08 0 5.5647e-08 0 5.565e-08 0.000231 5.5653e-08 0 5.6047e-08 0 5.605e-08 0.000231 5.6053e-08 0 5.6447e-08 0 5.645e-08 0.000231 5.6453e-08 0 5.6847e-08 0 5.685e-08 0.000231 5.6853e-08 0 5.7247e-08 0 5.725e-08 0.000231 5.7253e-08 0 5.7647e-08 0 5.765e-08 0.000231 5.7653e-08 0 5.8047e-08 0 5.805e-08 0.000231 5.8053e-08 0 5.8447e-08 0 5.845e-08 0.000231 5.8453e-08 0 5.8847e-08 0 5.885e-08 0.000231 5.8853e-08 0 5.9247e-08 0 5.925e-08 0.000231 5.9253e-08 0 5.9647e-08 0 5.965e-08 0.000231 5.9653e-08 0 6.0047e-08 0 6.005e-08 0.000231 6.0053e-08 0 6.0447e-08 0 6.045e-08 0.000231 6.0453e-08 0 6.0847e-08 0 6.085e-08 0.000231 6.0853e-08 0 6.1247e-08 0 6.125e-08 0.000231 6.1253e-08 0 6.1647e-08 0 6.165e-08 0.000231 6.1653e-08 0 6.2047e-08 0 6.205e-08 0.000231 6.2053e-08 0 6.2447e-08 0 6.245e-08 0.000231 6.2453e-08 0 6.2847e-08 0 6.285e-08 0.000231 6.2853e-08 0 6.3247e-08 0 6.325e-08 0.000231 6.3253e-08 0 6.3647e-08 0 6.365e-08 0.000231 6.3653e-08 0 6.4047e-08 0 6.405e-08 0.000231 6.4053e-08 0 6.4447e-08 0 6.445e-08 0.000231 6.4453e-08 0 6.4847e-08 0 6.485e-08 0.000231 6.4853e-08 0 6.5247e-08 0 6.525e-08 0.000231 6.5253e-08 0 6.5647e-08 0 6.565e-08 0.000231 6.5653e-08 0 6.6047e-08 0 6.605e-08 0.000231 6.6053e-08 0 6.6447e-08 0 6.645e-08 0.000231 6.6453e-08 0 6.6847e-08 0 6.685e-08 0.000231 6.6853e-08 0 6.7247e-08 0 6.725e-08 0.000231 6.7253e-08 0 6.7647e-08 0 6.765e-08 0.000231 6.7653e-08 0 6.8047e-08 0 6.805e-08 0.000231 6.8053e-08 0 6.8447e-08 0 6.845e-08 0.000231 6.8453e-08 0 6.8847e-08 0 6.885e-08 0.000231 6.8853e-08 0 6.9247e-08 0 6.925e-08 0.000231 6.9253e-08 0 6.9647e-08 0 6.965e-08 0.000231 6.9653e-08 0 7.0047e-08 0 7.005e-08 0.000231 7.0053e-08 0 7.0447e-08 0 7.045e-08 0.000231 7.0453e-08 0 7.0847e-08 0 7.085e-08 0.000231 7.0853e-08 0 7.1247e-08 0 7.125e-08 0.000231 7.1253e-08 0 7.1647e-08 0 7.165e-08 0.000231 7.1653e-08 0 7.2047e-08 0 7.205e-08 0.000231 7.2053e-08 0 7.2447e-08 0 7.245e-08 0.000231 7.2453e-08 0 7.2847e-08 0 7.285e-08 0.000231 7.2853e-08 0 7.3247e-08 0 7.325e-08 0.000231 7.3253e-08 0 7.3647e-08 0 7.365e-08 0.000231 7.3653e-08 0 7.4047e-08 0 7.405e-08 0.000231 7.4053e-08 0 7.4447e-08 0 7.445e-08 0.000231 7.4453e-08 0 7.4847e-08 0 7.485e-08 0.000231 7.4853e-08 0 7.5247e-08 0 7.525e-08 0.000231 7.5253e-08 0 7.5647e-08 0 7.565e-08 0.000231 7.5653e-08 0 7.6047e-08 0 7.605e-08 0.000231 7.6053e-08 0 7.6447e-08 0 7.645e-08 0.000231 7.6453e-08 0 7.6847e-08 0 7.685e-08 0.000231 7.6853e-08 0 7.7247e-08 0 7.725e-08 0.000231 7.7253e-08 0 7.7647e-08 0 7.765e-08 0.000231 7.7653e-08 0 7.8047e-08 0 7.805e-08 0.000231 7.8053e-08 0 7.8447e-08 0 7.845e-08 0.000231 7.8453e-08 0 7.8847e-08 0 7.885e-08 0.000231 7.8853e-08 0 7.9247e-08 0 7.925e-08 0.000231 7.9253e-08 0 7.9647e-08 0 7.965e-08 0.000231 7.9653e-08 0 8.0047e-08 0 8.005e-08 0.000231 8.0053e-08 0 8.0447e-08 0 8.045e-08 0.000231 8.0453e-08 0 8.0847e-08 0 8.085e-08 0.000231 8.0853e-08 0 8.1247e-08 0 8.125e-08 0.000231 8.1253e-08 0 8.1647e-08 0 8.165e-08 0.000231 8.1653e-08 0 8.2047e-08 0 8.205e-08 0.000231 8.2053e-08 0 8.2447e-08 0 8.245e-08 0.000231 8.2453e-08 0 8.2847e-08 0 8.285e-08 0.000231 8.2853e-08 0 8.3247e-08 0 8.325e-08 0.000231 8.3253e-08 0 8.3647e-08 0 8.365e-08 0.000231 8.3653e-08 0 8.4047e-08 0 8.405e-08 0.000231 8.4053e-08 0 8.4447e-08 0 8.445e-08 0.000231 8.4453e-08 0 8.4847e-08 0 8.485e-08 0.000231 8.4853e-08 0 8.5247e-08 0 8.525e-08 0.000231 8.5253e-08 0 8.5647e-08 0 8.565e-08 0.000231 8.5653e-08 0 8.6047e-08 0 8.605e-08 0.000231 8.6053e-08 0 8.6447e-08 0 8.645e-08 0.000231 8.6453e-08 0 8.6847e-08 0 8.685e-08 0.000231 8.6853e-08 0 8.7247e-08 0 8.725e-08 0.000231 8.7253e-08 0 8.7647e-08 0 8.765e-08 0.000231 8.7653e-08 0 8.8047e-08 0 8.805e-08 0.000231 8.8053e-08 0 8.8447e-08 0 8.845e-08 0.000231 8.8453e-08 0 8.8847e-08 0 8.885e-08 0.000231 8.8853e-08 0 8.9247e-08 0 8.925e-08 0.000231 8.9253e-08 0 8.9647e-08 0 8.965e-08 0.000231 8.9653e-08 0 9.0047e-08 0 9.005e-08 0.000231 9.0053e-08 0 9.0447e-08 0 9.045e-08 0.000231 9.0453e-08 0 9.0847e-08 0 9.085e-08 0.000231 9.0853e-08 0 9.1247e-08 0 9.125e-08 0.000231 9.1253e-08 0 9.1647e-08 0 9.165e-08 0.000231 9.1653e-08 0 9.2047e-08 0 9.205e-08 0.000231 9.2053e-08 0 9.2447e-08 0 9.245e-08 0.000231 9.2453e-08 0 9.2847e-08 0 9.285e-08 0.000231 9.2853e-08 0 9.3247e-08 0 9.325e-08 0.000231 9.3253e-08 0 9.3647e-08 0 9.365e-08 0.000231 9.3653e-08 0 9.4047e-08 0 9.405e-08 0.000231 9.4053e-08 0 9.4447e-08 0 9.445e-08 0.000231 9.4453e-08 0 9.4847e-08 0 9.485e-08 0.000231 9.4853e-08 0 9.5247e-08 0 9.525e-08 0.000231 9.5253e-08 0 9.5647e-08 0 9.565e-08 0.000231 9.5653e-08 0 9.6047e-08 0 9.605e-08 0.000231 9.6053e-08 0 9.6447e-08 0 9.645e-08 0.000231 9.6453e-08 0 9.6847e-08 0 9.685e-08 0.000231 9.6853e-08 0 9.7247e-08 0 9.725e-08 0.000231 9.7253e-08 0 9.7647e-08 0 9.765e-08 0.000231 9.7653e-08 0 9.8047e-08 0 9.805e-08 0.000231 9.8053e-08 0 9.8447e-08 0 9.845e-08 0.000231 9.8453e-08 0 9.8847e-08 0 9.885e-08 0.000231 9.8853e-08 0 9.9247e-08 0 9.925e-08 0.000231 9.9253e-08 0 9.9647e-08 0 9.965e-08 0.000231 9.9653e-08 0 1.00047e-07 0 1.0005e-07 0.000231 1.00053e-07 0 1.00447e-07 0 1.0045e-07 0.000231 1.00453e-07 0 1.00847e-07 0 1.0085e-07 0.000231 1.00853e-07 0 1.01247e-07 0 1.0125e-07 0.000231 1.01253e-07 0 1.01647e-07 0 1.0165e-07 0.000231 1.01653e-07 0 1.02047e-07 0 1.0205e-07 0.000231 1.02053e-07 0 1.02447e-07 0 1.0245e-07 0.000231 1.02453e-07 0 1.02847e-07 0 1.0285e-07 0.000231 1.02853e-07 0 1.03247e-07 0 1.0325e-07 0.000231 1.03253e-07 0 1.03647e-07 0 1.0365e-07 0.000231 1.03653e-07 0 1.04047e-07 0 1.0405e-07 0.000231 1.04053e-07 0 1.04447e-07 0 1.0445e-07 0.000231 1.04453e-07 0 1.04847e-07 0 1.0485e-07 0.000231 1.04853e-07 0 1.05247e-07 0 1.0525e-07 0.000231 1.05253e-07 0 1.05647e-07 0 1.0565e-07 0.000231 1.05653e-07 0 1.06047e-07 0 1.0605e-07 0.000231 1.06053e-07 0 1.06447e-07 0 1.0645e-07 0.000231 1.06453e-07 0 1.06847e-07 0 1.0685e-07 0.000231 1.06853e-07 0 1.07247e-07 0 1.0725e-07 0.000231 1.07253e-07 0 1.07647e-07 0 1.0765e-07 0.000231 1.07653e-07 0 1.08047e-07 0 1.0805e-07 0.000231 1.08053e-07 0 1.08447e-07 0 1.0845e-07 0.000231 1.08453e-07 0 1.08847e-07 0 1.0885e-07 0.000231 1.08853e-07 0 1.09247e-07 0 1.0925e-07 0.000231 1.09253e-07 0 1.09647e-07 0 1.0965e-07 0.000231 1.09653e-07 0 1.10047e-07 0 1.1005e-07 0.000231 1.10053e-07 0 1.10447e-07 0 1.1045e-07 0.000231 1.10453e-07 0 1.10847e-07 0 1.1085e-07 0.000231 1.10853e-07 0 1.11247e-07 0 1.1125e-07 0.000231 1.11253e-07 0 1.11647e-07 0 1.1165e-07 0.000231 1.11653e-07 0 1.12047e-07 0 1.1205e-07 0.000231 1.12053e-07 0 1.12447e-07 0 1.1245e-07 0.000231 1.12453e-07 0 1.12847e-07 0 1.1285e-07 0.000231 1.12853e-07 0 1.13247e-07 0 1.1325e-07 0.000231 1.13253e-07 0 1.13647e-07 0 1.1365e-07 0.000231 1.13653e-07 0 1.14047e-07 0 1.1405e-07 0.000231 1.14053e-07 0 1.14447e-07 0 1.1445e-07 0.000231 1.14453e-07 0 1.14847e-07 0 1.1485e-07 0.000231 1.14853e-07 0 1.15247e-07 0 1.1525e-07 0.000231 1.15253e-07 0 1.15647e-07 0 1.1565e-07 0.000231 1.15653e-07 0 1.16047e-07 0 1.1605e-07 0.000231 1.16053e-07 0 1.16447e-07 0 1.1645e-07 0.000231 1.16453e-07 0 1.16847e-07 0 1.1685e-07 0.000231 1.16853e-07 0 1.17247e-07 0 1.1725e-07 0.000231 1.17253e-07 0 1.17647e-07 0 1.1765e-07 0.000231 1.17653e-07 0 1.18047e-07 0 1.1805e-07 0.000231 1.18053e-07 0 1.18447e-07 0 1.1845e-07 0.000231 1.18453e-07 0 1.18847e-07 0 1.1885e-07 0.000231 1.18853e-07 0 1.19247e-07 0 1.1925e-07 0.000231 1.19253e-07 0 1.19647e-07 0 1.1965e-07 0.000231 1.19653e-07 0 1.20047e-07 0 1.2005e-07 0.000231 1.20053e-07 0 1.20447e-07 0 1.2045e-07 0.000231 1.20453e-07 0 1.20847e-07 0 1.2085e-07 0.000231 1.20853e-07 0 1.21247e-07 0 1.2125e-07 0.000231 1.21253e-07 0 1.21647e-07 0 1.2165e-07 0.000231 1.21653e-07 0 1.22047e-07 0 1.2205e-07 0.000231 1.22053e-07 0 1.22447e-07 0 1.2245e-07 0.000231 1.22453e-07 0 1.22847e-07 0 1.2285e-07 0.000231 1.22853e-07 0 1.23247e-07 0 1.2325e-07 0.000231 1.23253e-07 0 1.23647e-07 0 1.2365e-07 0.000231 1.23653e-07 0 1.24047e-07 0 1.2405e-07 0.000231 1.24053e-07 0 1.24447e-07 0 1.2445e-07 0.000231 1.24453e-07 0 1.24847e-07 0 1.2485e-07 0.000231 1.24853e-07 0 1.25247e-07 0 1.2525e-07 0.000231 1.25253e-07 0 1.25647e-07 0 1.2565e-07 0.000231 1.25653e-07 0 1.26047e-07 0 1.2605e-07 0.000231 1.26053e-07 0 1.26447e-07 0 1.2645e-07 0.000231 1.26453e-07 0 1.26847e-07 0 1.2685e-07 0.000231 1.26853e-07 0 1.27247e-07 0 1.2725e-07 0.000231 1.27253e-07 0 1.27647e-07 0 1.2765e-07 0.000231 1.27653e-07 0 1.28047e-07 0 1.2805e-07 0.000231 1.28053e-07 0 1.28447e-07 0 1.2845e-07 0.000231 1.28453e-07 0 1.28847e-07 0 1.2885e-07 0.000231 1.28853e-07 0 1.29247e-07 0 1.2925e-07 0.000231 1.29253e-07 0 1.29647e-07 0 1.2965e-07 0.000231 1.29653e-07 0 1.30047e-07 0 1.3005e-07 0.000231 1.30053e-07 0 1.30447e-07 0 1.3045e-07 0.000231 1.30453e-07 0 1.30847e-07 0 1.3085e-07 0.000231 1.30853e-07 0 1.31247e-07 0 1.3125e-07 0.000231 1.31253e-07 0 1.31647e-07 0 1.3165e-07 0.000231 1.31653e-07 0 1.32047e-07 0 1.3205e-07 0.000231 1.32053e-07 0 1.32447e-07 0 1.3245e-07 0.000231 1.32453e-07 0 1.32847e-07 0 1.3285e-07 0.000231 1.32853e-07 0 1.33247e-07 0 1.3325e-07 0.000231 1.33253e-07 0 1.33647e-07 0 1.3365e-07 0.000231 1.33653e-07 0 1.34047e-07 0 1.3405e-07 0.000231 1.34053e-07 0 1.34447e-07 0 1.3445e-07 0.000231 1.34453e-07 0 1.34847e-07 0 1.3485e-07 0.000231 1.34853e-07 0 1.35247e-07 0 1.3525e-07 0.000231 1.35253e-07 0 1.35647e-07 0 1.3565e-07 0.000231 1.35653e-07 0 1.36047e-07 0 1.3605e-07 0.000231 1.36053e-07 0 1.36447e-07 0 1.3645e-07 0.000231 1.36453e-07 0 1.36847e-07 0 1.3685e-07 0.000231 1.36853e-07 0 1.37247e-07 0 1.3725e-07 0.000231 1.37253e-07 0 1.37647e-07 0 1.3765e-07 0.000231 1.37653e-07 0 1.38047e-07 0 1.3805e-07 0.000231 1.38053e-07 0 1.38447e-07 0 1.3845e-07 0.000231 1.38453e-07 0 1.38847e-07 0 1.3885e-07 0.000231 1.38853e-07 0 1.39247e-07 0 1.3925e-07 0.000231 1.39253e-07 0 1.39647e-07 0 1.3965e-07 0.000231 1.39653e-07 0 1.40047e-07 0 1.4005e-07 0.000231 1.40053e-07 0 1.40447e-07 0 1.4045e-07 0.000231 1.40453e-07 0 1.40847e-07 0 1.4085e-07 0.000231 1.40853e-07 0 1.41247e-07 0 1.4125e-07 0.000231 1.41253e-07 0 1.41647e-07 0 1.4165e-07 0.000231 1.41653e-07 0 1.42047e-07 0 1.4205e-07 0.000231 1.42053e-07 0 1.42447e-07 0 1.4245e-07 0.000231 1.42453e-07 0 1.42847e-07 0 1.4285e-07 0.000231 1.42853e-07 0 1.43247e-07 0 1.4325e-07 0.000231 1.43253e-07 0 1.43647e-07 0 1.4365e-07 0.000231 1.43653e-07 0 1.44047e-07 0 1.4405e-07 0.000231 1.44053e-07 0 1.44447e-07 0 1.4445e-07 0.000231 1.44453e-07 0 1.44847e-07 0 1.4485e-07 0.000231 1.44853e-07 0 1.45247e-07 0 1.4525e-07 0.000231 1.45253e-07 0 1.45647e-07 0 1.4565e-07 0.000231 1.45653e-07 0 1.46047e-07 0 1.4605e-07 0.000231 1.46053e-07 0 1.46447e-07 0 1.4645e-07 0.000231 1.46453e-07 0 1.46847e-07 0 1.4685e-07 0.000231 1.46853e-07 0 1.47247e-07 0 1.4725e-07 0.000231 1.47253e-07 0 1.47647e-07 0 1.4765e-07 0.000231 1.47653e-07 0 1.48047e-07 0 1.4805e-07 0.000231 1.48053e-07 0 1.48447e-07 0 1.4845e-07 0.000231 1.48453e-07 0 1.48847e-07 0 1.4885e-07 0.000231 1.48853e-07 0 1.49247e-07 0 1.4925e-07 0.000231 1.49253e-07 0 1.49647e-07 0 1.4965e-07 0.000231 1.49653e-07 0 1.50047e-07 0 1.5005e-07 0.000231 1.50053e-07 0 1.50447e-07 0 1.5045e-07 0.000231 1.50453e-07 0 1.50847e-07 0 1.5085e-07 0.000231 1.50853e-07 0 1.51247e-07 0 1.5125e-07 0.000231 1.51253e-07 0 1.51647e-07 0 1.5165e-07 0.000231 1.51653e-07 0 1.52047e-07 0 1.5205e-07 0.000231 1.52053e-07 0 1.52447e-07 0 1.5245e-07 0.000231 1.52453e-07 0 1.52847e-07 0 1.5285e-07 0.000231 1.52853e-07 0 1.53247e-07 0 1.5325e-07 0.000231 1.53253e-07 0 1.53647e-07 0 1.5365e-07 0.000231 1.53653e-07 0 1.54047e-07 0 1.5405e-07 0.000231 1.54053e-07 0 1.54447e-07 0 1.5445e-07 0.000231 1.54453e-07 0 1.54847e-07 0 1.5485e-07 0.000231 1.54853e-07 0 1.55247e-07 0 1.5525e-07 0.000231 1.55253e-07 0 1.55647e-07 0 1.5565e-07 0.000231 1.55653e-07 0 1.56047e-07 0 1.5605e-07 0.000231 1.56053e-07 0 1.56447e-07 0 1.5645e-07 0.000231 1.56453e-07 0 1.56847e-07 0 1.5685e-07 0.000231 1.56853e-07 0 1.57247e-07 0 1.5725e-07 0.000231 1.57253e-07 0 1.57647e-07 0 1.5765e-07 0.000231 1.57653e-07 0 1.58047e-07 0 1.5805e-07 0.000231 1.58053e-07 0 1.58447e-07 0 1.5845e-07 0.000231 1.58453e-07 0 1.58847e-07 0 1.5885e-07 0.000231 1.58853e-07 0 1.59247e-07 0 1.5925e-07 0.000231 1.59253e-07 0)
L_TFF|6 CLK _TFF|1  2.63e-12
B_TFF|11 _TFF|1 _TFF|2 JJMIT_ADJ 
B_TFF|10 _TFF|2 0 JJMIT_ADJ 
L_TFF|8 _TFF|2 SUM0  5.26e-12
B_TFF|12 _TFF|2 _TFF|4 JJMIT_ADJ 
B_TFF|6 _TFF|4 _TFF|6 JJMIT_ADJ AREA=3.8
L_TFF|1 _TFF|3 _TFF|4  5.26e-12
L_TFF|3 _TFF|3 CBAR  5.26e-12
B_TFF|1 _TFF|3 0 JJMIT_ADJ AREA=5.0
B_TFF|2 _TFF|3 _TFF|5 JJMIT_ADJ AREA=5.0
B_TFF|5 _TFF|5 _TFF|6 JJMIT_ADJ AREA=2.5
L_TFF|4 _TFF|6 CARRY0  5.26e-12
B_TFF|4 _TFF|6 0 JJMIT_ADJ AREA=2.5
L_TFF|2 _TFF|5 _TFF|7  1.3e-12
B_TFF|3 _TFF|7 0 JJMIT_ADJ AREA=5.0
L_TFF|7 _TFF|7 A  3.9e-12
BSUM|1 SUM|1 SUM|2 JJMIT AREA=2.5
BSUM|2 SUM|4 SUM|5 JJMIT AREA=2.5
BSUM|3 SUM|7 SUM|8 JJMIT AREA=2.5
BSUM|4 SUM|10 SUM|11 JJMIT AREA=2.5
ISUM|B1 0 SUM|3  PWL(0 0 5e-12 0.000175)
ISUM|B2 0 SUM|6  PWL(0 0 5e-12 0.0002375)
ISUM|B3 0 SUM|9  PWL(0 0 5e-12 0.0002375)
ISUM|B4 0 SUM|12  PWL(0 0 5e-12 0.000175)
LSUM|1 SUM1 SUM|1  2.067833848e-12
LSUM|2 SUM|1 SUM|4  4.135667696e-12
LSUM|3 SUM|4 SUM|7  4.135667696e-12
LSUM|4 SUM|7 SUM|10  4.135667696e-12
LSUM|5 SUM|10 SUM  2.067833848e-12
LSUM|P1 SUM|2 0  5e-13
LSUM|P2 SUM|5 0  5e-13
LSUM|P3 SUM|8 0  5e-13
LSUM|P4 SUM|11 0  5e-13
LSUM|B1 SUM|1 SUM|3  2e-12
LSUM|B2 SUM|4 SUM|6  2e-12
LSUM|B3 SUM|7 SUM|9  2e-12
LSUM|B4 SUM|10 SUM|12  2e-12
RSUM|B1 SUM|1 SUM|101  2.7439617672
RSUM|B2 SUM|4 SUM|104  2.7439617672
RSUM|B3 SUM|7 SUM|107  2.7439617672
RSUM|B4 SUM|10 SUM|110  2.7439617672
LSUM|RB1 SUM|101 0  2.050338398468e-12
LSUM|RB2 SUM|104 0  2.050338398468e-12
LSUM|RB3 SUM|107 0  2.050338398468e-12
LSUM|RB4 SUM|110 0  2.050338398468e-12
BQ|1 Q|1 Q|2 JJMIT AREA=2.5
BQ|2 Q|4 Q|5 JJMIT AREA=2.5
BQ|3 Q|7 Q|8 JJMIT AREA=2.5
BQ|4 Q|10 Q|11 JJMIT AREA=2.5
IQ|B1 0 Q|3  PWL(0 0 5e-12 0.000175)
IQ|B2 0 Q|6  PWL(0 0 5e-12 0.0002375)
IQ|B3 0 Q|9  PWL(0 0 5e-12 0.0002375)
IQ|B4 0 Q|12  PWL(0 0 5e-12 0.000175)
LQ|1 CARRY1 Q|1  2.067833848e-12
LQ|2 Q|1 Q|4  4.135667696e-12
LQ|3 Q|4 Q|7  4.135667696e-12
LQ|4 Q|7 Q|10  4.135667696e-12
LQ|5 Q|10 CARRY  2.067833848e-12
LQ|P1 Q|2 0  5e-13
LQ|P2 Q|5 0  5e-13
LQ|P3 Q|8 0  5e-13
LQ|P4 Q|11 0  5e-13
LQ|B1 Q|1 Q|3  2e-12
LQ|B2 Q|4 Q|6  2e-12
LQ|B3 Q|7 Q|9  2e-12
LQ|B4 Q|10 Q|12  2e-12
RQ|B1 Q|1 Q|101  2.7439617672
RQ|B2 Q|4 Q|104  2.7439617672
RQ|B3 Q|7 Q|107  2.7439617672
RQ|B4 Q|10 Q|110  2.7439617672
LQ|RB1 Q|101 0  2.050338398468e-12
LQ|RB2 Q|104 0  2.050338398468e-12
LQ|RB3 Q|107 0  2.050338398468e-12
LQ|RB4 Q|110 0  2.050338398468e-12
L_TFF|I1|B _TFF|3 _TFF|I1|MID  2e-12
I_TFF|I1|B 0 _TFF|I1|MID  PWL(0 0 5e-12 0.00019)
L_TFF|I2|B _TFF|7 _TFF|I2|MID  2e-12
I_TFF|I2|B 0 _TFF|I2|MID  PWL(0 0 5e-12 0.00019)
.print DEVI LINPUT
.print DEVI LSUM
.print DEVI RSUM
.print DEVI LCARRY
.print DEVI RCARRY
.print DEVI RCBAR
.print DEVI IDATA|H
.print DEVI IT1|T
.print DEVI L_TFF|6
.print DEVI B_TFF|11
.print DEVI B_TFF|10
.print DEVI L_TFF|8
.print DEVI B_TFF|12
.print DEVI B_TFF|6
.print DEVI L_TFF|1
.print DEVI L_TFF|3
.print DEVI B_TFF|1
.print DEVI B_TFF|2
.print DEVI B_TFF|5
.print DEVI L_TFF|4
.print DEVI B_TFF|4
.print DEVI L_TFF|2
.print DEVI B_TFF|3
.print DEVI L_TFF|7
.print DEVI BSUM|1
.print DEVI BSUM|2
.print DEVI BSUM|3
.print DEVI BSUM|4
.print DEVI ISUM|B1
.print DEVI ISUM|B2
.print DEVI ISUM|B3
.print DEVI ISUM|B4
.print DEVI LSUM|1
.print DEVI LSUM|2
.print DEVI LSUM|3
.print DEVI LSUM|4
.print DEVI LSUM|5
.print DEVI LSUM|P1
.print DEVI LSUM|P2
.print DEVI LSUM|P3
.print DEVI LSUM|P4
.print DEVI LSUM|B1
.print DEVI LSUM|B2
.print DEVI LSUM|B3
.print DEVI LSUM|B4
.print DEVI RSUM|B1
.print DEVI RSUM|B2
.print DEVI RSUM|B3
.print DEVI RSUM|B4
.print DEVI LSUM|RB1
.print DEVI LSUM|RB2
.print DEVI LSUM|RB3
.print DEVI LSUM|RB4
.print DEVI BQ|1
.print DEVI BQ|2
.print DEVI BQ|3
.print DEVI BQ|4
.print DEVI IQ|B1
.print DEVI IQ|B2
.print DEVI IQ|B3
.print DEVI IQ|B4
.print DEVI LQ|1
.print DEVI LQ|2
.print DEVI LQ|3
.print DEVI LQ|4
.print DEVI LQ|5
.print DEVI LQ|P1
.print DEVI LQ|P2
.print DEVI LQ|P3
.print DEVI LQ|P4
.print DEVI LQ|B1
.print DEVI LQ|B2
.print DEVI LQ|B3
.print DEVI LQ|B4
.print DEVI RQ|B1
.print DEVI RQ|B2
.print DEVI RQ|B3
.print DEVI RQ|B4
.print DEVI LQ|RB1
.print DEVI LQ|RB2
.print DEVI LQ|RB3
.print DEVI LQ|RB4
.print V SUM|8
.print V Q|7
.print V _TFF|2
.print V Q|110
.print V SUM1
.print V Q|6
.print V Q|5
.print V Q|11
.print V SUM|104
.print V Q|1
.print V CBAR
.print V Q|4
.print V Q|9
.print V Q|104
.print V CARRY
.print V A
.print V SUM|9
.print V SUM|12
.print V Q|2
.print V _TFF|6
.print V SUM|11
.print V SUM0
.print V CLK0
.print V _TFF|5
.print V _TFF|7
.print V _TFF|3
.print V SUM|10
.print V SUM|107
.print V SUM|3
.print V Q|10
.print V Q|101
.print V SUM|6
.print V SUM|1
.print V SUM|7
.print V CARRY1
.print V SUM|5
.print V Q|3
.print V CARRY0
.print V _TFF|1
.print V Q|12
.print V SUM|101
.print V SUM|2
.print V SUM
.print V _TFF|4
.print V SUM|4
.print V Q|107
.print V Q|8
.print V SUM|110
.print V CLK
.print DEVP B_TFF|11
.print DEVP B_TFF|10
.print DEVP B_TFF|12
.print DEVP B_TFF|6
.print DEVP B_TFF|1
.print DEVP B_TFF|2
.print DEVP B_TFF|5
.print DEVP B_TFF|4
.print DEVP B_TFF|3
.print DEVP BSUM|1
.print DEVP BSUM|2
.print DEVP BSUM|3
.print DEVP BSUM|4
.print DEVP BQ|1
.print DEVP BQ|2
.print DEVP BQ|3
.print DEVP BQ|4
