*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM IU=1.25e-05
.PARAM VU=0.0006857
.PARAM LU=2.632e-12
.PARAM JCRIT=0.0001
.PARAM OFFSET1=5e-11
.PARAM TCLOCK=2.5e-10
.PARAM DO=6.25e-11
.PARAM ZED0=2.5
.PARAM IMAX=0.0005
.PARAM TR=9.5e-12
.PARAM TF=9.5e-12
.PARAM PW=1e-12
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMITLL100 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JMITLL JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160OHM, RN=16OHM, ICRIT=0.1MA)
TCLK  CLK_RX 0 CLK 0 LOSSLESS Z0=ZED0 TD=10P
TA  A_RX 0 A 0 LOSSLESS Z0=ZED0 TD=10P
.TRAN 0.25E-12 2.6E-9
ICLK 0 CLK_DC  PULSE(0 IMAX OFFSET1 TR TF PW TCLOCK)
IA1_1 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+1*TCLOCK TR TF PW 8*TCLOCK)
IA1_2 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+3*TCLOCK TR TF PW 8*TCLOCK)
IA1_3 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+5*TCLOCK TR TF PW 8*TCLOCK)
IA1_4 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+7*TCLOCK TR TF PW 8*TCLOCK)
IA2_1 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+2*TCLOCK TR TF PW 8*TCLOCK)
IA2_2 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+3*TCLOCK TR TF PW 8*TCLOCK)
IA2_3 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+6*TCLOCK TR TF PW 8*TCLOCK)
IA2_4 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+7*TCLOCK TR TF PW 8*TCLOCK)
IA3_1 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+4*TCLOCK TR TF PW 8*TCLOCK)
IA3_2 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+5*TCLOCK TR TF PW 8*TCLOCK)
IA3_3 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+6*TCLOCK TR TF PW 8*TCLOCK)
IA3_4 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+7*TCLOCK TR TF PW 8*TCLOCK)
RSUM SUM 0  1
RCARRY CARRY 0  1
RCBAR CBAR 0  1
LDCSFQCLK|1 CLK_DC DCSFQCLK|1  1e-12
RDCSFQCLK|2 DCSFQCLK|1 0  5
LDCSFQCLK|3 DCSFQCLK|1 DCSFQCLK|2  6e-13
BDCSFQCLK|1 DCSFQCLK|2 DCSFQCLK|3 JJMIT AREA=2.25
RDCSFQCLK|B1 DCSFQCLK|2 DCSFQCLK|102  3.048846408
LDCSFQCLK|RB1 DCSFQCLK|102 DCSFQCLK|3  1.7225982205200002e-12
LDCSFQCLK|4 DCSFQCLK|3 DCSFQCLK|5  1.1e-12
BDCSFQCLK|2 DCSFQCLK|5 DCSFQCLK|6 JJMIT AREA=2.25
LDCSFQCLK|P2 DCSFQCLK|6 0  5e-13
RDCSFQCLK|B2 DCSFQCLK|5 DCSFQCLK|105  3.048846408
LDCSFQCLK|RB2 DCSFQCLK|105 0  2.2225982205200003e-12
LDCSFQCLK|5 DCSFQCLK|5 DCSFQCLK|7  4.5e-12
BDCSFQCLK|3 DCSFQCLK|7 DCSFQCLK|8 JJMIT AREA=2.5
LDCSFQCLK|P3 DCSFQCLK|8 0  5e-13
RDCSFQCLK|B3 DCSFQCLK|7 DCSFQCLK|107  2.7439617672
LDCSFQCLK|RB3 DCSFQCLK|107 0  2.050338398468e-12
IDCSFQCLK|B1 0 DCSFQCLK|4  PWL(0 0 5e-12 0.000196429)
LDCSFQCLK|B1 DCSFQCLK|4 DCSFQCLK|3  2e-12
IDCSFQCLK|B2 0 DCSFQCLK|9  PWL(0 0 5e-12 0.000175)
LDCSFQCLK|B2 DCSFQCLK|9 DCSFQCLK|7  2e-12
LDCSFQCLK|6 DCSFQCLK|7 CLK0  2.067833848e-12
BJTLCLK|1 JTLCLK|1 JTLCLK|6 JJMITLL100 AREA=2.5
BJTLCLK|2 JTLCLK|4 JTLCLK|8 JJMITLL100 AREA=2.5
IJTLCLK|B1 0 JTLCLK|3  PWL(0 0 5e-12 0.00035)
LJTLCLK|1 CLK0 JTLCLK|1  2e-12
LJTLCLK|2 JTLCLK|1 JTLCLK|3  2e-12
LJTLCLK|3 JTLCLK|3 JTLCLK|4  2e-12
LJTLCLK|4 JTLCLK|4 JTLCLK|5  2e-12
LJTLCLK|B1 JTLCLK|7 JTLCLK|6  1e-12
LJTLCLK|B2 JTLCLK|9 JTLCLK|8  1e-12
LJTLCLK|P1 JTLCLK|6 0  2e-13
LJTLCLK|P2 JTLCLK|8 0  2e-13
RJTLCLK|B1 JTLCLK|1 JTLCLK|7  3.88
RJTLCLK|B2 JTLCLK|4 JTLCLK|9  3.88
LDCSFQ_1|1 A1_DC DCSFQ_1|1  1e-12
RDCSFQ_1|2 DCSFQ_1|1 0  5
LDCSFQ_1|3 DCSFQ_1|1 DCSFQ_1|2  6e-13
BDCSFQ_1|1 DCSFQ_1|2 DCSFQ_1|3 JJMIT AREA=2.25
RDCSFQ_1|B1 DCSFQ_1|2 DCSFQ_1|102  3.048846408
LDCSFQ_1|RB1 DCSFQ_1|102 DCSFQ_1|3  1.7225982205200002e-12
LDCSFQ_1|4 DCSFQ_1|3 DCSFQ_1|5  1.1e-12
BDCSFQ_1|2 DCSFQ_1|5 DCSFQ_1|6 JJMIT AREA=2.25
LDCSFQ_1|P2 DCSFQ_1|6 0  5e-13
RDCSFQ_1|B2 DCSFQ_1|5 DCSFQ_1|105  3.048846408
LDCSFQ_1|RB2 DCSFQ_1|105 0  2.2225982205200003e-12
LDCSFQ_1|5 DCSFQ_1|5 DCSFQ_1|7  4.5e-12
BDCSFQ_1|3 DCSFQ_1|7 DCSFQ_1|8 JJMIT AREA=2.5
LDCSFQ_1|P3 DCSFQ_1|8 0  5e-13
RDCSFQ_1|B3 DCSFQ_1|7 DCSFQ_1|107  2.7439617672
LDCSFQ_1|RB3 DCSFQ_1|107 0  2.050338398468e-12
IDCSFQ_1|B1 0 DCSFQ_1|4  PWL(0 0 5e-12 0.000196429)
LDCSFQ_1|B1 DCSFQ_1|4 DCSFQ_1|3  2e-12
IDCSFQ_1|B2 0 DCSFQ_1|9  PWL(0 0 5e-12 0.000175)
LDCSFQ_1|B2 DCSFQ_1|9 DCSFQ_1|7  2e-12
LDCSFQ_1|6 DCSFQ_1|7 A1  2.067833848e-12
BJTL_1|1 JTL_1|1 JTL_1|6 JJMITLL100 AREA=2.5
BJTL_1|2 JTL_1|4 JTL_1|8 JJMITLL100 AREA=2.5
IJTL_1|B1 0 JTL_1|3  PWL(0 0 5e-12 0.00035)
LJTL_1|1 A1 JTL_1|1  2e-12
LJTL_1|2 JTL_1|1 JTL_1|3  2e-12
LJTL_1|3 JTL_1|3 JTL_1|4  2e-12
LJTL_1|4 JTL_1|4 JTL_1|5  2e-12
LJTL_1|B1 JTL_1|7 JTL_1|6  1e-12
LJTL_1|B2 JTL_1|9 JTL_1|8  1e-12
LJTL_1|P1 JTL_1|6 0  2e-13
LJTL_1|P2 JTL_1|8 0  2e-13
RJTL_1|B1 JTL_1|1 JTL_1|7  3.88
RJTL_1|B2 JTL_1|4 JTL_1|9  3.88
L_TFF|6 _TFF|READOUT _TFF|1  5.26e-12
B_TFF|11 _TFF|1 _TFF|2 JJMIT AREA=2.2
B_TFF|10 _TFF|2 0 JJMIT AREA=1.4999999999999998
L_TFF|8 _TFF|2 _TFF|SUM_TX  3.9e-12
B_TFF|12 _TFF|2 _TFF|4 JJMIT AREA=1.25
B_TFF|6 _TFF|4 _TFF|6 JJMIT AREA=1.9
L_TFF|1 _TFF|3 _TFF|4  2.104e-11
L_TFF|3 _TFF|3 _TFF|CBAR_TX  5.26e-12
B_TFF|1 _TFF|3 0 JJMIT AREA=2.5
B_TFF|2 _TFF|3 _TFF|5 JJMIT AREA=2.5
B_TFF|5 _TFF|5 _TFF|6 JJMIT AREA=1.25
L_TFF|4 _TFF|6 _TFF|CARRY_TX  5.26e-12
B_TFF|4 _TFF|6 0 JJMIT AREA=1.25
L_TFF|2 _TFF|5 _TFF|7  2.6e-12
B_TFF|3 _TFF|7 0 JJMIT AREA=2.75
L_TFF|7 _TFF|7 _TFF|TOGGLE  2.63e-12
BJTLCLK|POUT|01 JTLCLK|POUT|3 JTLCLK|POUT|7 JMITLL AREA=2
BJTLCLK|POUT|02 JTLCLK|POUT|4 JTLCLK|POUT|6 JMITLL AREA=1.62
IJTLCLK|POUT|B01 0 JTLCLK|POUT|10  PWL(0 0 5e-12 0.00023)
IJTLCLK|POUT|B02 0 JTLCLK|POUT|11  PWL(0 0 5e-12 8.2e-05)
LJTLCLK|POUT|01 JTLCLK|5 JTLCLK|POUT|3  2.5e-12
LJTLCLK|POUT|02 JTLCLK|POUT|3 JTLCLK|POUT|4  3.3e-12
LJTLCLK|POUT|03 JTLCLK|POUT|4 JTLCLK|POUT|5  3.5e-13
LJTLCLK|POUT|P01 0 JTLCLK|POUT|7  5e-14
LJTLCLK|POUT|P02 0 JTLCLK|POUT|6  1.2e-13
LJTLCLK|POUT|PR01 JTLCLK|POUT|3 JTLCLK|POUT|10  2e-13
LJTLCLK|POUT|PR02 JTLCLK|POUT|4 JTLCLK|POUT|11  1.3e-12
LJTLCLK|POUT|RB01 JTLCLK|POUT|7 JTLCLK|POUT|8  1e-12
LJTLCLK|POUT|RB02 JTLCLK|POUT|6 JTLCLK|POUT|9  1e-12
RJTLCLK|POUT|B01 JTLCLK|POUT|8 JTLCLK|POUT|3  4.85
RJTLCLK|POUT|B02 JTLCLK|POUT|9 JTLCLK|POUT|4  6.3
RJTLCLK|POUT|INS JTLCLK|POUT|5 CLK_RX  1.36
BJTL_1|POUT|01 JTL_1|POUT|3 JTL_1|POUT|7 JMITLL AREA=2
BJTL_1|POUT|02 JTL_1|POUT|4 JTL_1|POUT|6 JMITLL AREA=1.62
IJTL_1|POUT|B01 0 JTL_1|POUT|10  PWL(0 0 5e-12 0.00023)
IJTL_1|POUT|B02 0 JTL_1|POUT|11  PWL(0 0 5e-12 8.2e-05)
LJTL_1|POUT|01 JTL_1|5 JTL_1|POUT|3  2.5e-12
LJTL_1|POUT|02 JTL_1|POUT|3 JTL_1|POUT|4  3.3e-12
LJTL_1|POUT|03 JTL_1|POUT|4 JTL_1|POUT|5  3.5e-13
LJTL_1|POUT|P01 0 JTL_1|POUT|7  5e-14
LJTL_1|POUT|P02 0 JTL_1|POUT|6  1.2e-13
LJTL_1|POUT|PR01 JTL_1|POUT|3 JTL_1|POUT|10  2e-13
LJTL_1|POUT|PR02 JTL_1|POUT|4 JTL_1|POUT|11  1.3e-12
LJTL_1|POUT|RB01 JTL_1|POUT|7 JTL_1|POUT|8  1e-12
LJTL_1|POUT|RB02 JTL_1|POUT|6 JTL_1|POUT|9  1e-12
RJTL_1|POUT|B01 JTL_1|POUT|8 JTL_1|POUT|3  4.85
RJTL_1|POUT|B02 JTL_1|POUT|9 JTL_1|POUT|4  6.3
RJTL_1|POUT|INS JTL_1|POUT|5 A_RX  1.36
B_TFF|_READOUT|01 _TFF|_READOUT|1 _TFF|_READOUT|9 JMITLL AREA=1
B_TFF|_READOUT|02 _TFF|_READOUT|4 _TFF|_READOUT|8 JMITLL AREA=1
B_TFF|_READOUT|03 _TFF|_READOUT|5 _TFF|_READOUT|7 JMITLL AREA=1
I_TFF|_READOUT|B01 0 _TFF|_READOUT|10  PWL(0 0 5e-12 0.0002015)
L_TFF|_READOUT|01 CLK _TFF|_READOUT|1  2e-13
L_TFF|_READOUT|02 _TFF|_READOUT|1 _TFF|_READOUT|3  4.3e-12
L_TFF|_READOUT|03 _TFF|_READOUT|3 _TFF|_READOUT|4  4.6e-12
L_TFF|_READOUT|04 _TFF|_READOUT|4 _TFF|_READOUT|5  5e-12
L_TFF|_READOUT|05 _TFF|_READOUT|5 _TFF|READOUT  2.3e-12
L_TFF|_READOUT|P01 0 _TFF|_READOUT|9  3.4e-13
L_TFF|_READOUT|P02 0 _TFF|_READOUT|8  6e-14
L_TFF|_READOUT|P03 0 _TFF|_READOUT|7  3e-14
L_TFF|_READOUT|PR01 _TFF|_READOUT|3 _TFF|_READOUT|10  2e-13
L_TFF|_READOUT|RB01 _TFF|_READOUT|9 _TFF|_READOUT|11  5e-13
L_TFF|_READOUT|RB02 _TFF|_READOUT|8 _TFF|_READOUT|12  1e-12
L_TFF|_READOUT|RB03 _TFF|_READOUT|7 _TFF|_READOUT|13  1e-12
R_TFF|_READOUT|B01 _TFF|_READOUT|11 _TFF|_READOUT|1  9.7
R_TFF|_READOUT|B02 _TFF|_READOUT|12 _TFF|_READOUT|4  9.7
R_TFF|_READOUT|B03 _TFF|_READOUT|13 _TFF|_READOUT|5  9.7
B_TFF|_TOGGLE|01 _TFF|_TOGGLE|1 _TFF|_TOGGLE|9 JMITLL AREA=1
B_TFF|_TOGGLE|02 _TFF|_TOGGLE|4 _TFF|_TOGGLE|8 JMITLL AREA=1
B_TFF|_TOGGLE|03 _TFF|_TOGGLE|5 _TFF|_TOGGLE|7 JMITLL AREA=1
I_TFF|_TOGGLE|B01 0 _TFF|_TOGGLE|10  PWL(0 0 5e-12 0.000155)
L_TFF|_TOGGLE|01 A _TFF|_TOGGLE|1  2e-13
L_TFF|_TOGGLE|02 _TFF|_TOGGLE|1 _TFF|_TOGGLE|3  4.3e-12
L_TFF|_TOGGLE|03 _TFF|_TOGGLE|3 _TFF|_TOGGLE|4  4.6e-12
L_TFF|_TOGGLE|04 _TFF|_TOGGLE|4 _TFF|_TOGGLE|5  5e-12
L_TFF|_TOGGLE|05 _TFF|_TOGGLE|5 _TFF|TOGGLE  2.3e-12
L_TFF|_TOGGLE|P01 0 _TFF|_TOGGLE|9  3.4e-13
L_TFF|_TOGGLE|P02 0 _TFF|_TOGGLE|8  6e-14
L_TFF|_TOGGLE|P03 0 _TFF|_TOGGLE|7  3e-14
L_TFF|_TOGGLE|PR01 _TFF|_TOGGLE|3 _TFF|_TOGGLE|10  2e-13
L_TFF|_TOGGLE|RB01 _TFF|_TOGGLE|9 _TFF|_TOGGLE|11  5e-13
L_TFF|_TOGGLE|RB02 _TFF|_TOGGLE|8 _TFF|_TOGGLE|12  1e-12
L_TFF|_TOGGLE|RB03 _TFF|_TOGGLE|7 _TFF|_TOGGLE|13  1e-12
R_TFF|_TOGGLE|B01 _TFF|_TOGGLE|11 _TFF|_TOGGLE|1  9.7
R_TFF|_TOGGLE|B02 _TFF|_TOGGLE|12 _TFF|_TOGGLE|4  9.7
R_TFF|_TOGGLE|B03 _TFF|_TOGGLE|13 _TFF|_TOGGLE|5  9.7
B_TFF|_SUM|01 _TFF|_SUM|3 _TFF|_SUM|7 JMITLL AREA=2
B_TFF|_SUM|02 _TFF|_SUM|4 _TFF|_SUM|6 JMITLL AREA=1.62
I_TFF|_SUM|B01 0 _TFF|_SUM|10  PWL(0 0 5e-12 0.00023)
I_TFF|_SUM|B02 0 _TFF|_SUM|11  PWL(0 0 5e-12 8.2e-05)
L_TFF|_SUM|01 _TFF|SUM_TX _TFF|_SUM|3  2.5e-12
L_TFF|_SUM|02 _TFF|_SUM|3 _TFF|_SUM|4  3.3e-12
L_TFF|_SUM|03 _TFF|_SUM|4 _TFF|_SUM|5  3.5e-13
L_TFF|_SUM|P01 0 _TFF|_SUM|7  5e-14
L_TFF|_SUM|P02 0 _TFF|_SUM|6  1.2e-13
L_TFF|_SUM|PR01 _TFF|_SUM|3 _TFF|_SUM|10  2e-13
L_TFF|_SUM|PR02 _TFF|_SUM|4 _TFF|_SUM|11  1.3e-12
L_TFF|_SUM|RB01 _TFF|_SUM|7 _TFF|_SUM|8  1e-12
L_TFF|_SUM|RB02 _TFF|_SUM|6 _TFF|_SUM|9  1e-12
R_TFF|_SUM|B01 _TFF|_SUM|8 _TFF|_SUM|3  4.85
R_TFF|_SUM|B02 _TFF|_SUM|9 _TFF|_SUM|4  6.3
R_TFF|_SUM|INS _TFF|_SUM|5 SUM  1.36
B_TFF|_CARRY|01 _TFF|_CARRY|3 _TFF|_CARRY|7 JMITLL AREA=2
B_TFF|_CARRY|02 _TFF|_CARRY|4 _TFF|_CARRY|6 JMITLL AREA=1.62
I_TFF|_CARRY|B01 0 _TFF|_CARRY|10  PWL(0 0 5e-12 0.00023)
I_TFF|_CARRY|B02 0 _TFF|_CARRY|11  PWL(0 0 5e-12 8.2e-05)
L_TFF|_CARRY|01 _TFF|CARRY_TX _TFF|_CARRY|3  2.5e-12
L_TFF|_CARRY|02 _TFF|_CARRY|3 _TFF|_CARRY|4  3.3e-12
L_TFF|_CARRY|03 _TFF|_CARRY|4 _TFF|_CARRY|5  3.5e-13
L_TFF|_CARRY|P01 0 _TFF|_CARRY|7  5e-14
L_TFF|_CARRY|P02 0 _TFF|_CARRY|6  1.2e-13
L_TFF|_CARRY|PR01 _TFF|_CARRY|3 _TFF|_CARRY|10  2e-13
L_TFF|_CARRY|PR02 _TFF|_CARRY|4 _TFF|_CARRY|11  1.3e-12
L_TFF|_CARRY|RB01 _TFF|_CARRY|7 _TFF|_CARRY|8  1e-12
L_TFF|_CARRY|RB02 _TFF|_CARRY|6 _TFF|_CARRY|9  1e-12
R_TFF|_CARRY|B01 _TFF|_CARRY|8 _TFF|_CARRY|3  4.85
R_TFF|_CARRY|B02 _TFF|_CARRY|9 _TFF|_CARRY|4  6.3
R_TFF|_CARRY|INS _TFF|_CARRY|5 CARRY  1.36
B_TFF|_CBAR|01 _TFF|_CBAR|3 _TFF|_CBAR|7 JMITLL AREA=2
B_TFF|_CBAR|02 _TFF|_CBAR|4 _TFF|_CBAR|6 JMITLL AREA=1.62
I_TFF|_CBAR|B01 0 _TFF|_CBAR|10  PWL(0 0 5e-12 0.00023)
I_TFF|_CBAR|B02 0 _TFF|_CBAR|11  PWL(0 0 5e-12 8.2e-05)
L_TFF|_CBAR|01 _TFF|CBAR_TX _TFF|_CBAR|3  2.5e-12
L_TFF|_CBAR|02 _TFF|_CBAR|3 _TFF|_CBAR|4  3.3e-12
L_TFF|_CBAR|03 _TFF|_CBAR|4 _TFF|_CBAR|5  3.5e-13
L_TFF|_CBAR|P01 0 _TFF|_CBAR|7  5e-14
L_TFF|_CBAR|P02 0 _TFF|_CBAR|6  1.2e-13
L_TFF|_CBAR|PR01 _TFF|_CBAR|3 _TFF|_CBAR|10  2e-13
L_TFF|_CBAR|PR02 _TFF|_CBAR|4 _TFF|_CBAR|11  1.3e-12
L_TFF|_CBAR|RB01 _TFF|_CBAR|7 _TFF|_CBAR|8  1e-12
L_TFF|_CBAR|RB02 _TFF|_CBAR|6 _TFF|_CBAR|9  1e-12
R_TFF|_CBAR|B01 _TFF|_CBAR|8 _TFF|_CBAR|3  4.85
R_TFF|_CBAR|B02 _TFF|_CBAR|9 _TFF|_CBAR|4  6.3
R_TFF|_CBAR|INS _TFF|_CBAR|5 CBAR  1.36
L_TFF|I1|B _TFF|3 _TFF|I1|MID  2e-12
I_TFF|I1|B 0 _TFF|I1|MID  PWL(0 0 5e-12 0.000228)
L_TFF|I2|B _TFF|7 _TFF|I2|MID  2e-12
I_TFF|I2|B 0 _TFF|I2|MID  PWL(0 0 5e-12 0.000133)
.print DEVI ICLK
.print DEVI IA1_1
.print DEVI IA1_2
.print DEVI IA1_3
.print DEVI IA1_4
.print DEVI IA2_1
.print DEVI IA2_2
.print DEVI IA2_3
.print DEVI IA2_4
.print DEVI IA3_1
.print DEVI IA3_2
.print DEVI IA3_3
.print DEVI IA3_4
.print DEVI RSUM
.print DEVI RCARRY
.print DEVI RCBAR
.print DEVI LDCSFQCLK|1
.print DEVI RDCSFQCLK|2
.print DEVI LDCSFQCLK|3
.print DEVI BDCSFQCLK|1
.print DEVI RDCSFQCLK|B1
.print DEVI LDCSFQCLK|RB1
.print DEVI LDCSFQCLK|4
.print DEVI BDCSFQCLK|2
.print DEVI LDCSFQCLK|P2
.print DEVI RDCSFQCLK|B2
.print DEVI LDCSFQCLK|RB2
.print DEVI LDCSFQCLK|5
.print DEVI BDCSFQCLK|3
.print DEVI LDCSFQCLK|P3
.print DEVI RDCSFQCLK|B3
.print DEVI LDCSFQCLK|RB3
.print DEVI IDCSFQCLK|B1
.print DEVI LDCSFQCLK|B1
.print DEVI IDCSFQCLK|B2
.print DEVI LDCSFQCLK|B2
.print DEVI LDCSFQCLK|6
.print DEVI BJTLCLK|1
.print DEVI BJTLCLK|2
.print DEVI IJTLCLK|B1
.print DEVI LJTLCLK|1
.print DEVI LJTLCLK|2
.print DEVI LJTLCLK|3
.print DEVI LJTLCLK|4
.print DEVI LJTLCLK|B1
.print DEVI LJTLCLK|B2
.print DEVI LJTLCLK|P1
.print DEVI LJTLCLK|P2
.print DEVI RJTLCLK|B1
.print DEVI RJTLCLK|B2
.print DEVI LDCSFQ_1|1
.print DEVI RDCSFQ_1|2
.print DEVI LDCSFQ_1|3
.print DEVI BDCSFQ_1|1
.print DEVI RDCSFQ_1|B1
.print DEVI LDCSFQ_1|RB1
.print DEVI LDCSFQ_1|4
.print DEVI BDCSFQ_1|2
.print DEVI LDCSFQ_1|P2
.print DEVI RDCSFQ_1|B2
.print DEVI LDCSFQ_1|RB2
.print DEVI LDCSFQ_1|5
.print DEVI BDCSFQ_1|3
.print DEVI LDCSFQ_1|P3
.print DEVI RDCSFQ_1|B3
.print DEVI LDCSFQ_1|RB3
.print DEVI IDCSFQ_1|B1
.print DEVI LDCSFQ_1|B1
.print DEVI IDCSFQ_1|B2
.print DEVI LDCSFQ_1|B2
.print DEVI LDCSFQ_1|6
.print DEVI BJTL_1|1
.print DEVI BJTL_1|2
.print DEVI IJTL_1|B1
.print DEVI LJTL_1|1
.print DEVI LJTL_1|2
.print DEVI LJTL_1|3
.print DEVI LJTL_1|4
.print DEVI LJTL_1|B1
.print DEVI LJTL_1|B2
.print DEVI LJTL_1|P1
.print DEVI LJTL_1|P2
.print DEVI RJTL_1|B1
.print DEVI RJTL_1|B2
.print DEVI L_TFF|6
.print DEVI B_TFF|11
.print DEVI B_TFF|10
.print DEVI L_TFF|8
.print DEVI B_TFF|12
.print DEVI B_TFF|6
.print DEVI L_TFF|1
.print DEVI L_TFF|3
.print DEVI B_TFF|1
.print DEVI B_TFF|2
.print DEVI B_TFF|5
.print DEVI L_TFF|4
.print DEVI B_TFF|4
.print DEVI L_TFF|2
.print DEVI B_TFF|3
.print DEVI L_TFF|7
.print V CLK_RX
.print V JTL_1|4
.print V JTL_1|1
.print V DCSFQ_1|2
.print V _TFF|READOUT
.print V DCSFQCLK|2
.print V _TFF|4
.print V SUM
.print V _TFF|5
.print V JTL_1|7
.print V JTLCLK|1
.print V _TFF|TOGGLE
.print V DCSFQCLK|8
.print V JTLCLK|3
.print V CLK0
.print V JTLCLK|6
.print V JTLCLK|4
.print V A_RX
.print V DCSFQ_1|5
.print V JTL_1|5
.print V DCSFQ_1|102
.print V DCSFQ_1|6
.print V _TFF|SUM_TX
.print V JTLCLK|8
.print V DCSFQ_1|8
.print V JTL_1|6
.print V DCSFQCLK|107
.print V A1
.print V DCSFQCLK|102
.print V DCSFQ_1|107
.print V DCSFQ_1|7
.print V DCSFQCLK|6
.print V _TFF|7
.print V CARRY
.print V _TFF|CBAR_TX
.print V DCSFQCLK|1
.print V JTL_1|3
.print V DCSFQCLK|4
.print V _TFF|6
.print V CLK
.print V DCSFQCLK|105
.print V CBAR
.print V A1_DC
.print V DCSFQ_1|105
.print V DCSFQ_1|9
.print V DCSFQ_1|4
.print V _TFF|CARRY_TX
.print V DCSFQCLK|9
.print V JTLCLK|9
.print V DCSFQ_1|3
.print V _TFF|1
.print V _TFF|3
.print V DCSFQ_1|1
.print V DCSFQCLK|5
.print V JTL_1|9
.print V JTLCLK|5
.print V DCSFQCLK|7
.print V JTLCLK|7
.print V DCSFQCLK|3
.print V A
.print V CLK_DC
.print V _TFF|2
.print V JTL_1|8
.print DEVP BDCSFQCLK|1
.print DEVP BDCSFQCLK|2
.print DEVP BDCSFQCLK|3
.print DEVP BJTLCLK|1
.print DEVP BJTLCLK|2
.print DEVP BDCSFQ_1|1
.print DEVP BDCSFQ_1|2
.print DEVP BDCSFQ_1|3
.print DEVP BJTL_1|1
.print DEVP BJTL_1|2
.print DEVP B_TFF|11
.print DEVP B_TFF|10
.print DEVP B_TFF|12
.print DEVP B_TFF|6
.print DEVP B_TFF|1
.print DEVP B_TFF|2
.print DEVP B_TFF|5
.print DEVP B_TFF|4
.print DEVP B_TFF|3
.print DEVP BJTLCLK|POUT|01
.print DEVP BJTLCLK|POUT|02
.print DEVP BJTL_1|POUT|01
.print DEVP BJTL_1|POUT|02
.print DEVP B_TFF|_READOUT|01
.print DEVP B_TFF|_READOUT|02
.print DEVP B_TFF|_READOUT|03
.print DEVP B_TFF|_TOGGLE|01
.print DEVP B_TFF|_TOGGLE|02
.print DEVP B_TFF|_TOGGLE|03
.print DEVP B_TFF|_SUM|01
.print DEVP B_TFF|_SUM|02
.print DEVP B_TFF|_CARRY|01
.print DEVP B_TFF|_CARRY|02
.print DEVP B_TFF|_CBAR|01
.print DEVP B_TFF|_CBAR|02
