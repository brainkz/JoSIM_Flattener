*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM TCLOCK=6.1e-11
.PARAM OS=3.0499999999999997e-12
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 2000E-12
R_S0 S0 0  1
R_S1 S1 0  1
R_S2 S2 0  1
R_S3 S3 0  1
R_S4 S4 0  1
I_VEC|A0 0 A0  PWL(0 0 1.408e-11 0 1.708e-11 0.0007 2.008e-11 0 1.3608e-10 0 1.3908e-10 0.0007 1.4208e-10 0 1.9708e-10 0 2.0008e-10 0.0007 2.0308e-10 0 2.5808e-10 0 2.6108e-10 0.0007 2.6408e-10 0 3.1908e-10 0 3.2208e-10 0.0007 3.2508e-10 0 4.4108e-10 0 4.4408e-10 0.0007 4.4708e-10 0 5.0208e-10 0 5.0508e-10 0.0007 5.0808e-10 0 6.2408e-10 0 6.2708e-10 0.0007 6.3008e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|A1 0 A1  PWL(0 0 1.9708e-10 0 2.0008e-10 0.0007 2.0308e-10 0 2.5808e-10 0 2.6108e-10 0.0007 2.6408e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|A2 0 A2  PWL(0 0 7.508e-11 0 7.808e-11 0.0007 8.108e-11 0 2.5808e-10 0 2.6108e-10 0.0007 2.6408e-10 0 3.8008e-10 0 3.8308e-10 0.0007 3.8608e-10 0 5.0208e-10 0 5.0508e-10 0.0007 5.0808e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|A3 0 A3  PWL(0 0 3.8008e-10 0 3.8308e-10 0.0007 3.8608e-10 0 5.0208e-10 0 5.0508e-10 0.0007 5.0808e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|B0 0 B0  PWL(0 0 1.408e-11 0 1.708e-11 0.0007 2.008e-11 0 1.3608e-10 0 1.3908e-10 0.0007 1.4208e-10 0 3.1908e-10 0 3.2208e-10 0.0007 3.2508e-10 0 4.4108e-10 0 4.4408e-10 0.0007 4.4708e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|B1 0 B1  PWL(0 0 1.408e-11 0 1.708e-11 0.0007 2.008e-11 0 1.3608e-10 0 1.3908e-10 0.0007 1.4208e-10 0 1.9708e-10 0 2.0008e-10 0.0007 2.0308e-10 0 2.5808e-10 0 2.6108e-10 0.0007 2.6408e-10 0 5.6308e-10 0 5.6608e-10 0.0007 5.6908e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|B2 0 B2  PWL(0 0 1.408e-11 0 1.708e-11 0.0007 2.008e-11 0 7.508e-11 0 7.808e-11 0.0007 8.108e-11 0 1.3608e-10 0 1.3908e-10 0.0007 1.4208e-10 0 2.5808e-10 0 2.6108e-10 0.0007 2.6408e-10 0 3.1908e-10 0 3.2208e-10 0.0007 3.2508e-10 0 4.4108e-10 0 4.4408e-10 0.0007 4.4708e-10 0 5.0208e-10 0 5.0508e-10 0.0007 5.0808e-10 0 5.6308e-10 0 5.6608e-10 0.0007 5.6908e-10 0 6.2408e-10 0 6.2708e-10 0.0007 6.3008e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
I_VEC|B3 0 B3  PWL(0 0 1.408e-11 0 1.708e-11 0.0007 2.008e-11 0 7.508e-11 0 7.808e-11 0.0007 8.108e-11 0 1.9708e-10 0 2.0008e-10 0.0007 2.0308e-10 0 4.4108e-10 0 4.4408e-10 0.0007 4.4708e-10 0 6.2408e-10 0 6.2708e-10 0.0007 6.3008e-10 0 6.8508e-10 0 6.8808e-10 0.0007 6.9108e-10 0)
IT00|T 0 T00  PWL(0 0 9.2e-12 0 1.22e-11 0.0021 1.52e-11 0 7.02e-11 0 7.32e-11 0.0021 7.62e-11 0 1.312e-10 0 1.342e-10 0.0021 1.372e-10 0 1.922e-10 0 1.952e-10 0.0021 1.982e-10 0 2.532e-10 0 2.562e-10 0.0021 2.592e-10 0 3.142e-10 0 3.172e-10 0.0021 3.202e-10 0 3.752e-10 0 3.782e-10 0.0021 3.812e-10 0 4.362e-10 0 4.392e-10 0.0021 4.422e-10 0 4.972e-10 0 5.002e-10 0.0021 5.032e-10 0 5.582e-10 0 5.612e-10 0.0021 5.642e-10 0 6.192e-10 0 6.222e-10 0.0021 6.252e-10 0 6.802e-10 0 6.832e-10 0.0021 6.862e-10 0 7.412e-10 0 7.442e-10 0.0021 7.472e-10 0 8.022e-10 0 8.052e-10 0.0021 8.082e-10 0 8.632e-10 0 8.662e-10 0.0021 8.692e-10 0 9.242e-10 0 9.272e-10 0.0021 9.302e-10 0 9.852e-10 0 9.882e-10 0.0021 9.912e-10 0 1.0462e-09 0 1.0492e-09 0.0021 1.0522e-09 0 1.1072e-09 0 1.1102e-09 0.0021 1.1132e-09 0 1.1682e-09 0 1.1712e-09 0.0021 1.1742e-09 0 1.2292e-09 0 1.2322e-09 0.0021 1.2352e-09 0 1.2902e-09 0 1.2932e-09 0.0021 1.2962e-09 0 1.3512e-09 0 1.3542e-09 0.0021 1.3572e-09 0 1.4122e-09 0 1.4152e-09 0.0021 1.4182e-09 0 1.4732e-09 0 1.4762e-09 0.0021 1.4792e-09 0 1.5342e-09 0 1.5372e-09 0.0021 1.5402e-09 0 1.5952e-09 0 1.5982e-09 0.0021 1.6012e-09 0 1.6562e-09 0 1.6592e-09 0.0021 1.6622e-09 0 1.7172e-09 0 1.7202e-09 0.0021 1.7232e-09 0 1.7782e-09 0 1.7812e-09 0.0021 1.7842e-09 0 1.8392e-09 0 1.8422e-09 0.0021 1.8452e-09 0 1.9002e-09 0 1.9032e-09 0.0021 1.9062e-09 0 1.9612e-09 0 1.9642e-09 0.0021 1.9672e-09 0 2.0222e-09 0 2.0252e-09 0.0021 2.0282e-09 0 2.0832e-09 0 2.0862e-09 0.0021 2.0892e-09 0 2.1442e-09 0 2.1472e-09 0.0021 2.1502e-09 0 2.2052e-09 0 2.2082e-09 0.0021 2.2112e-09 0 2.2662e-09 0 2.2692e-09 0.0021 2.2722e-09 0 2.3272e-09 0 2.3302e-09 0.0021 2.3332e-09 0 2.3882e-09 0 2.3912e-09 0.0021 2.3942e-09 0 2.4492e-09 0 2.4522e-09 0.0021 2.4552e-09 0 2.5102e-09 0 2.5132e-09 0.0021 2.5162e-09 0 2.5712e-09 0 2.5742e-09 0.0021 2.5772e-09 0 2.6322e-09 0 2.6352e-09 0.0021 2.6382e-09 0 2.6932e-09 0 2.6962e-09 0.0021 2.6992e-09 0 2.7542e-09 0 2.7572e-09 0.0021 2.7602e-09 0 2.8152e-09 0 2.8182e-09 0.0021 2.8212e-09 0 2.8762e-09 0 2.8792e-09 0.0021 2.8822e-09 0 2.9372e-09 0 2.9402e-09 0.0021 2.9432e-09 0 2.9982e-09 0 3.0012e-09 0.0021 3.0042e-09 0 3.0592e-09 0 3.0622e-09 0.0021 3.0652e-09 0 3.1202e-09 0 3.1232e-09 0.0021 3.1262e-09 0 3.1812e-09 0 3.1842e-09 0.0021 3.1872e-09 0 3.2422e-09 0 3.2452e-09 0.0021 3.2482e-09 0 3.3032e-09 0 3.3062e-09 0.0021 3.3092e-09 0 3.3642e-09 0 3.3672e-09 0.0021 3.3702e-09 0 3.4252e-09 0 3.4282e-09 0.0021 3.4312e-09 0 3.4862e-09 0 3.4892e-09 0.0021 3.4922e-09 0 3.5472e-09 0 3.5502e-09 0.0021 3.5532e-09 0 3.6082e-09 0 3.6112e-09 0.0021 3.6142e-09 0 3.6692e-09 0 3.6722e-09 0.0021 3.6752e-09 0 3.7302e-09 0 3.7332e-09 0.0021 3.7362e-09 0 3.7912e-09 0 3.7942e-09 0.0021 3.7972e-09 0 3.8522e-09 0 3.8552e-09 0.0021 3.8582e-09 0 3.9132e-09 0 3.9162e-09 0.0021 3.9192e-09 0 3.9742e-09 0 3.9772e-09 0.0021 3.9802e-09 0 4.0352e-09 0 4.0382e-09 0.0021 4.0412e-09 0 4.0962e-09 0 4.0992e-09 0.0021 4.1022e-09 0 4.1572e-09 0 4.1602e-09 0.0021 4.1632e-09 0 4.2182e-09 0 4.2212e-09 0.0021 4.2242e-09 0 4.2792e-09 0 4.2822e-09 0.0021 4.2852e-09 0 4.3402e-09 0 4.3432e-09 0.0021 4.3462e-09 0 4.4012e-09 0 4.4042e-09 0.0021 4.4072e-09 0 4.4622e-09 0 4.4652e-09 0.0021 4.4682e-09 0 4.5232e-09 0 4.5262e-09 0.0021 4.5292e-09 0 4.5842e-09 0 4.5872e-09 0.0021 4.5902e-09 0 4.6452e-09 0 4.6482e-09 0.0021 4.6512e-09 0 4.7062e-09 0 4.7092e-09 0.0021 4.7122e-09 0 4.7672e-09 0 4.7702e-09 0.0021 4.7732e-09 0 4.8282e-09 0 4.8312e-09 0.0021 4.8342e-09 0 4.8892e-09 0 4.8922e-09 0.0021 4.8952e-09 0 4.9502e-09 0 4.9532e-09 0.0021 4.9562e-09 0 5.0112e-09 0 5.0142e-09 0.0021 5.0172e-09 0 5.0722e-09 0 5.0752e-09 0.0021 5.0782e-09 0 5.1332e-09 0 5.1362e-09 0.0021 5.1392e-09 0 5.1942e-09 0 5.1972e-09 0.0021 5.2002e-09 0 5.2552e-09 0 5.2582e-09 0.0021 5.2612e-09 0 5.3162e-09 0 5.3192e-09 0.0021 5.3222e-09 0 5.3772e-09 0 5.3802e-09 0.0021 5.3832e-09 0 5.4382e-09 0 5.4412e-09 0.0021 5.4442e-09 0 5.4992e-09 0 5.5022e-09 0.0021 5.5052e-09 0 5.5602e-09 0 5.5632e-09 0.0021 5.5662e-09 0 5.6212e-09 0 5.6242e-09 0.0021 5.6272e-09 0 5.6822e-09 0 5.6852e-09 0.0021 5.6882e-09 0 5.7432e-09 0 5.7462e-09 0.0021 5.7492e-09 0 5.8042e-09 0 5.8072e-09 0.0021 5.8102e-09 0 5.8652e-09 0 5.8682e-09 0.0021 5.8712e-09 0 5.9262e-09 0 5.9292e-09 0.0021 5.9322e-09 0 5.9872e-09 0 5.9902e-09 0.0021 5.9932e-09 0 6.0482e-09 0 6.0512e-09 0.0021 6.0542e-09 0 6.1092e-09 0 6.1122e-09 0.0021 6.1152e-09 0 6.1702e-09 0 6.1732e-09 0.0021 6.1762e-09 0 6.2312e-09 0 6.2342e-09 0.0021 6.2372e-09 0 6.2922e-09 0 6.2952e-09 0.0021 6.2982e-09 0 6.3532e-09 0 6.3562e-09 0.0021 6.3592e-09 0 6.4142e-09 0 6.4172e-09 0.0021 6.4202e-09 0 6.4752e-09 0 6.4782e-09 0.0021 6.4812e-09 0 6.5362e-09 0 6.5392e-09 0.0021 6.5422e-09 0 6.5972e-09 0 6.6002e-09 0.0021 6.6032e-09 0 6.6582e-09 0 6.6612e-09 0.0021 6.6642e-09 0 6.7192e-09 0 6.7222e-09 0.0021 6.7252e-09 0 6.7802e-09 0 6.7832e-09 0.0021 6.7862e-09 0 6.8412e-09 0 6.8442e-09 0.0021 6.8472e-09 0 6.9022e-09 0 6.9052e-09 0.0021 6.9082e-09 0 6.9632e-09 0 6.9662e-09 0.0021 6.9692e-09 0 7.0242e-09 0 7.0272e-09 0.0021 7.0302e-09 0 7.0852e-09 0 7.0882e-09 0.0021 7.0912e-09 0 7.1462e-09 0 7.1492e-09 0.0021 7.1522e-09 0 7.2072e-09 0 7.2102e-09 0.0021 7.2132e-09 0 7.2682e-09 0 7.2712e-09 0.0021 7.2742e-09 0 7.3292e-09 0 7.3322e-09 0.0021 7.3352e-09 0 7.3902e-09 0 7.3932e-09 0.0021 7.3962e-09 0 7.4512e-09 0 7.4542e-09 0.0021 7.4572e-09 0 7.5122e-09 0 7.5152e-09 0.0021 7.5182e-09 0 7.5732e-09 0 7.5762e-09 0.0021 7.5792e-09 0 7.6342e-09 0 7.6372e-09 0.0021 7.6402e-09 0 7.6952e-09 0 7.6982e-09 0.0021 7.7012e-09 0 7.7562e-09 0 7.7592e-09 0.0021 7.7622e-09 0 7.8172e-09 0 7.8202e-09 0.0021 7.8232e-09 0 7.8782e-09 0 7.8812e-09 0.0021 7.8842e-09 0 7.9392e-09 0 7.9422e-09 0.0021 7.9452e-09 0 8.0002e-09 0 8.0032e-09 0.0021 8.0062e-09 0 8.0612e-09 0 8.0642e-09 0.0021 8.0672e-09 0 8.1222e-09 0 8.1252e-09 0.0021 8.1282e-09 0 8.1832e-09 0 8.1862e-09 0.0021 8.1892e-09 0 8.2442e-09 0 8.2472e-09 0.0021 8.2502e-09 0 8.3052e-09 0 8.3082e-09 0.0021 8.3112e-09 0 8.3662e-09 0 8.3692e-09 0.0021 8.3722e-09 0 8.4272e-09 0 8.4302e-09 0.0021 8.4332e-09 0 8.4882e-09 0 8.4912e-09 0.0021 8.4942e-09 0 8.5492e-09 0 8.5522e-09 0.0021 8.5552e-09 0 8.6102e-09 0 8.6132e-09 0.0021 8.6162e-09 0 8.6712e-09 0 8.6742e-09 0.0021 8.6772e-09 0 8.7322e-09 0 8.7352e-09 0.0021 8.7382e-09 0 8.7932e-09 0 8.7962e-09 0.0021 8.7992e-09 0 8.8542e-09 0 8.8572e-09 0.0021 8.8602e-09 0 8.9152e-09 0 8.9182e-09 0.0021 8.9212e-09 0 8.9762e-09 0 8.9792e-09 0.0021 8.9822e-09 0 9.0372e-09 0 9.0402e-09 0.0021 9.0432e-09 0 9.0982e-09 0 9.1012e-09 0.0021 9.1042e-09 0 9.1592e-09 0 9.1622e-09 0.0021 9.1652e-09 0 9.2202e-09 0 9.2232e-09 0.0021 9.2262e-09 0 9.2812e-09 0 9.2842e-09 0.0021 9.2872e-09 0 9.3422e-09 0 9.3452e-09 0.0021 9.3482e-09 0 9.4032e-09 0 9.4062e-09 0.0021 9.4092e-09 0 9.4642e-09 0 9.4672e-09 0.0021 9.4702e-09 0 9.5252e-09 0 9.5282e-09 0.0021 9.5312e-09 0 9.5862e-09 0 9.5892e-09 0.0021 9.5922e-09 0 9.6472e-09 0 9.6502e-09 0.0021 9.6532e-09 0 9.7082e-09 0 9.7112e-09 0.0021 9.7142e-09 0 9.7692e-09 0 9.7722e-09 0.0021 9.7752e-09 0 9.8302e-09 0 9.8332e-09 0.0021 9.8362e-09 0 9.8912e-09 0 9.8942e-09 0.0021 9.8972e-09 0 9.9522e-09 0 9.9552e-09 0.0021 9.9582e-09 0 1.00132e-08 0 1.00162e-08 0.0021 1.00192e-08 0 1.00742e-08 0 1.00772e-08 0.0021 1.00802e-08 0 1.01352e-08 0 1.01382e-08 0.0021 1.01412e-08 0 1.01962e-08 0 1.01992e-08 0.0021 1.02022e-08 0 1.02572e-08 0 1.02602e-08 0.0021 1.02632e-08 0 1.03182e-08 0 1.03212e-08 0.0021 1.03242e-08 0 1.03792e-08 0 1.03822e-08 0.0021 1.03852e-08 0 1.04402e-08 0 1.04432e-08 0.0021 1.04462e-08 0 1.05012e-08 0 1.05042e-08 0.0021 1.05072e-08 0 1.05622e-08 0 1.05652e-08 0.0021 1.05682e-08 0 1.06232e-08 0 1.06262e-08 0.0021 1.06292e-08 0 1.06842e-08 0 1.06872e-08 0.0021 1.06902e-08 0 1.07452e-08 0 1.07482e-08 0.0021 1.07512e-08 0 1.08062e-08 0 1.08092e-08 0.0021 1.08122e-08 0 1.08672e-08 0 1.08702e-08 0.0021 1.08732e-08 0 1.09282e-08 0 1.09312e-08 0.0021 1.09342e-08 0 1.09892e-08 0 1.09922e-08 0.0021 1.09952e-08 0 1.10502e-08 0 1.10532e-08 0.0021 1.10562e-08 0 1.11112e-08 0 1.11142e-08 0.0021 1.11172e-08 0 1.11722e-08 0 1.11752e-08 0.0021 1.11782e-08 0 1.12332e-08 0 1.12362e-08 0.0021 1.12392e-08 0 1.12942e-08 0 1.12972e-08 0.0021 1.13002e-08 0 1.13552e-08 0 1.13582e-08 0.0021 1.13612e-08 0 1.14162e-08 0 1.14192e-08 0.0021 1.14222e-08 0 1.14772e-08 0 1.14802e-08 0.0021 1.14832e-08 0 1.15382e-08 0 1.15412e-08 0.0021 1.15442e-08 0 1.15992e-08 0 1.16022e-08 0.0021 1.16052e-08 0 1.16602e-08 0 1.16632e-08 0.0021 1.16662e-08 0 1.17212e-08 0 1.17242e-08 0.0021 1.17272e-08 0 1.17822e-08 0 1.17852e-08 0.0021 1.17882e-08 0 1.18432e-08 0 1.18462e-08 0.0021 1.18492e-08 0 1.19042e-08 0 1.19072e-08 0.0021 1.19102e-08 0 1.19652e-08 0 1.19682e-08 0.0021 1.19712e-08 0 1.20262e-08 0 1.20292e-08 0.0021 1.20322e-08 0 1.20872e-08 0 1.20902e-08 0.0021 1.20932e-08 0 1.21482e-08 0 1.21512e-08 0.0021 1.21542e-08 0 1.22092e-08 0 1.22122e-08 0.0021 1.22152e-08 0 1.22702e-08 0 1.22732e-08 0.0021 1.22762e-08 0 1.23312e-08 0 1.23342e-08 0.0021 1.23372e-08 0 1.23922e-08 0 1.23952e-08 0.0021 1.23982e-08 0 1.24532e-08 0 1.24562e-08 0.0021 1.24592e-08 0 1.25142e-08 0 1.25172e-08 0.0021 1.25202e-08 0 1.25752e-08 0 1.25782e-08 0.0021 1.25812e-08 0 1.26362e-08 0 1.26392e-08 0.0021 1.26422e-08 0 1.26972e-08 0 1.27002e-08 0.0021 1.27032e-08 0 1.27582e-08 0 1.27612e-08 0.0021 1.27642e-08 0 1.28192e-08 0 1.28222e-08 0.0021 1.28252e-08 0 1.28802e-08 0 1.28832e-08 0.0021 1.28862e-08 0 1.29412e-08 0 1.29442e-08 0.0021 1.29472e-08 0 1.30022e-08 0 1.30052e-08 0.0021 1.30082e-08 0 1.30632e-08 0 1.30662e-08 0.0021 1.30692e-08 0 1.31242e-08 0 1.31272e-08 0.0021 1.31302e-08 0 1.31852e-08 0 1.31882e-08 0.0021 1.31912e-08 0 1.32462e-08 0 1.32492e-08 0.0021 1.32522e-08 0 1.33072e-08 0 1.33102e-08 0.0021 1.33132e-08 0 1.33682e-08 0 1.33712e-08 0.0021 1.33742e-08 0 1.34292e-08 0 1.34322e-08 0.0021 1.34352e-08 0 1.34902e-08 0 1.34932e-08 0.0021 1.34962e-08 0 1.35512e-08 0 1.35542e-08 0.0021 1.35572e-08 0 1.36122e-08 0 1.36152e-08 0.0021 1.36182e-08 0 1.36732e-08 0 1.36762e-08 0.0021 1.36792e-08 0 1.37342e-08 0 1.37372e-08 0.0021 1.37402e-08 0 1.37952e-08 0 1.37982e-08 0.0021 1.38012e-08 0 1.38562e-08 0 1.38592e-08 0.0021 1.38622e-08 0 1.39172e-08 0 1.39202e-08 0.0021 1.39232e-08 0 1.39782e-08 0 1.39812e-08 0.0021 1.39842e-08 0 1.40392e-08 0 1.40422e-08 0.0021 1.40452e-08 0 1.41002e-08 0 1.41032e-08 0.0021 1.41062e-08 0 1.41612e-08 0 1.41642e-08 0.0021 1.41672e-08 0 1.42222e-08 0 1.42252e-08 0.0021 1.42282e-08 0 1.42832e-08 0 1.42862e-08 0.0021 1.42892e-08 0 1.43442e-08 0 1.43472e-08 0.0021 1.43502e-08 0 1.44052e-08 0 1.44082e-08 0.0021 1.44112e-08 0 1.44662e-08 0 1.44692e-08 0.0021 1.44722e-08 0 1.45272e-08 0 1.45302e-08 0.0021 1.45332e-08 0 1.45882e-08 0 1.45912e-08 0.0021 1.45942e-08 0 1.46492e-08 0 1.46522e-08 0.0021 1.46552e-08 0 1.47102e-08 0 1.47132e-08 0.0021 1.47162e-08 0 1.47712e-08 0 1.47742e-08 0.0021 1.47772e-08 0 1.48322e-08 0 1.48352e-08 0.0021 1.48382e-08 0 1.48932e-08 0 1.48962e-08 0.0021 1.48992e-08 0 1.49542e-08 0 1.49572e-08 0.0021 1.49602e-08 0 1.50152e-08 0 1.50182e-08 0.0021 1.50212e-08 0 1.50762e-08 0 1.50792e-08 0.0021 1.50822e-08 0 1.51372e-08 0 1.51402e-08 0.0021 1.51432e-08 0 1.51982e-08 0 1.52012e-08 0.0021 1.52042e-08 0 1.52592e-08 0 1.52622e-08 0.0021 1.52652e-08 0 1.53202e-08 0 1.53232e-08 0.0021 1.53262e-08 0 1.53812e-08 0 1.53842e-08 0.0021 1.53872e-08 0 1.54422e-08 0 1.54452e-08 0.0021 1.54482e-08 0 1.55032e-08 0 1.55062e-08 0.0021 1.55092e-08 0 1.55642e-08 0 1.55672e-08 0.0021 1.55702e-08 0 1.56252e-08 0 1.56282e-08 0.0021 1.56312e-08 0 1.56862e-08 0 1.56892e-08 0.0021 1.56922e-08 0 1.57472e-08 0 1.57502e-08 0.0021 1.57532e-08 0 1.58082e-08 0 1.58112e-08 0.0021 1.58142e-08 0 1.58692e-08 0 1.58722e-08 0.0021 1.58752e-08 0 1.59302e-08 0 1.59332e-08 0.0021 1.59362e-08 0 1.59912e-08 0 1.59942e-08 0.0021 1.59972e-08 0 1.60522e-08 0 1.60552e-08 0.0021 1.60582e-08 0 1.61132e-08 0 1.61162e-08 0.0021 1.61192e-08 0 1.61742e-08 0 1.61772e-08 0.0021 1.61802e-08 0 1.62352e-08 0 1.62382e-08 0.0021 1.62412e-08 0 1.62962e-08 0 1.62992e-08 0.0021 1.63022e-08 0 1.63572e-08 0 1.63602e-08 0.0021 1.63632e-08 0 1.64182e-08 0 1.64212e-08 0.0021 1.64242e-08 0 1.64792e-08 0 1.64822e-08 0.0021 1.64852e-08 0 1.65402e-08 0 1.65432e-08 0.0021 1.65462e-08 0 1.66012e-08 0 1.66042e-08 0.0021 1.66072e-08 0 1.66622e-08 0 1.66652e-08 0.0021 1.66682e-08 0 1.67232e-08 0 1.67262e-08 0.0021 1.67292e-08 0 1.67842e-08 0 1.67872e-08 0.0021 1.67902e-08 0 1.68452e-08 0 1.68482e-08 0.0021 1.68512e-08 0 1.69062e-08 0 1.69092e-08 0.0021 1.69122e-08 0 1.69672e-08 0 1.69702e-08 0.0021 1.69732e-08 0 1.70282e-08 0 1.70312e-08 0.0021 1.70342e-08 0 1.70892e-08 0 1.70922e-08 0.0021 1.70952e-08 0 1.71502e-08 0 1.71532e-08 0.0021 1.71562e-08 0 1.72112e-08 0 1.72142e-08 0.0021 1.72172e-08 0 1.72722e-08 0 1.72752e-08 0.0021 1.72782e-08 0 1.73332e-08 0 1.73362e-08 0.0021 1.73392e-08 0 1.73942e-08 0 1.73972e-08 0.0021 1.74002e-08 0 1.74552e-08 0 1.74582e-08 0.0021 1.74612e-08 0 1.75162e-08 0 1.75192e-08 0.0021 1.75222e-08 0 1.75772e-08 0 1.75802e-08 0.0021 1.75832e-08 0 1.76382e-08 0 1.76412e-08 0.0021 1.76442e-08 0 1.76992e-08 0 1.77022e-08 0.0021 1.77052e-08 0 1.77602e-08 0 1.77632e-08 0.0021 1.77662e-08 0 1.78212e-08 0 1.78242e-08 0.0021 1.78272e-08 0 1.78822e-08 0 1.78852e-08 0.0021 1.78882e-08 0 1.79432e-08 0 1.79462e-08 0.0021 1.79492e-08 0 1.80042e-08 0 1.80072e-08 0.0021 1.80102e-08 0 1.80652e-08 0 1.80682e-08 0.0021 1.80712e-08 0 1.81262e-08 0 1.81292e-08 0.0021 1.81322e-08 0 1.81872e-08 0 1.81902e-08 0.0021 1.81932e-08 0 1.82482e-08 0 1.82512e-08 0.0021 1.82542e-08 0 1.83092e-08 0 1.83122e-08 0.0021 1.83152e-08 0 1.83702e-08 0 1.83732e-08 0.0021 1.83762e-08 0 1.84312e-08 0 1.84342e-08 0.0021 1.84372e-08 0 1.84922e-08 0 1.84952e-08 0.0021 1.84982e-08 0 1.85532e-08 0 1.85562e-08 0.0021 1.85592e-08 0 1.86142e-08 0 1.86172e-08 0.0021 1.86202e-08 0 1.86752e-08 0 1.86782e-08 0.0021 1.86812e-08 0 1.87362e-08 0 1.87392e-08 0.0021 1.87422e-08 0 1.87972e-08 0 1.88002e-08 0.0021 1.88032e-08 0 1.88582e-08 0 1.88612e-08 0.0021 1.88642e-08 0 1.89192e-08 0 1.89222e-08 0.0021 1.89252e-08 0 1.89802e-08 0 1.89832e-08 0.0021 1.89862e-08 0 1.90412e-08 0 1.90442e-08 0.0021 1.90472e-08 0 1.91022e-08 0 1.91052e-08 0.0021 1.91082e-08 0 1.91632e-08 0 1.91662e-08 0.0021 1.91692e-08 0 1.92242e-08 0 1.92272e-08 0.0021 1.92302e-08 0 1.92852e-08 0 1.92882e-08 0.0021 1.92912e-08 0 1.93462e-08 0 1.93492e-08 0.0021 1.93522e-08 0 1.94072e-08 0 1.94102e-08 0.0021 1.94132e-08 0 1.94682e-08 0 1.94712e-08 0.0021 1.94742e-08 0 1.95292e-08 0 1.95322e-08 0.0021 1.95352e-08 0 1.95902e-08 0 1.95932e-08 0.0021 1.95962e-08 0 1.96512e-08 0 1.96542e-08 0.0021 1.96572e-08 0 1.97122e-08 0 1.97152e-08 0.0021 1.97182e-08 0 1.97732e-08 0 1.97762e-08 0.0021 1.97792e-08 0 1.98342e-08 0 1.98372e-08 0.0021 1.98402e-08 0 1.98952e-08 0 1.98982e-08 0.0021 1.99012e-08 0 1.99562e-08 0 1.99592e-08 0.0021 1.99622e-08 0 2.00172e-08 0 2.00202e-08 0.0021 2.00232e-08 0 2.00782e-08 0 2.00812e-08 0.0021 2.00842e-08 0 2.01392e-08 0 2.01422e-08 0.0021 2.01452e-08 0 2.02002e-08 0 2.02032e-08 0.0021 2.02062e-08 0 2.02612e-08 0 2.02642e-08 0.0021 2.02672e-08 0 2.03222e-08 0 2.03252e-08 0.0021 2.03282e-08 0 2.03832e-08 0 2.03862e-08 0.0021 2.03892e-08 0 2.04442e-08 0 2.04472e-08 0.0021 2.04502e-08 0 2.05052e-08 0 2.05082e-08 0.0021 2.05112e-08 0 2.05662e-08 0 2.05692e-08 0.0021 2.05722e-08 0 2.06272e-08 0 2.06302e-08 0.0021 2.06332e-08 0 2.06882e-08 0 2.06912e-08 0.0021 2.06942e-08 0 2.07492e-08 0 2.07522e-08 0.0021 2.07552e-08 0 2.08102e-08 0 2.08132e-08 0.0021 2.08162e-08 0 2.08712e-08 0 2.08742e-08 0.0021 2.08772e-08 0 2.09322e-08 0 2.09352e-08 0.0021 2.09382e-08 0 2.09932e-08 0 2.09962e-08 0.0021 2.09992e-08 0 2.10542e-08 0 2.10572e-08 0.0021 2.10602e-08 0 2.11152e-08 0 2.11182e-08 0.0021 2.11212e-08 0 2.11762e-08 0 2.11792e-08 0.0021 2.11822e-08 0 2.12372e-08 0 2.12402e-08 0.0021 2.12432e-08 0 2.12982e-08 0 2.13012e-08 0.0021 2.13042e-08 0 2.13592e-08 0 2.13622e-08 0.0021 2.13652e-08 0 2.14202e-08 0 2.14232e-08 0.0021 2.14262e-08 0 2.14812e-08 0 2.14842e-08 0.0021 2.14872e-08 0 2.15422e-08 0 2.15452e-08 0.0021 2.15482e-08 0 2.16032e-08 0 2.16062e-08 0.0021 2.16092e-08 0 2.16642e-08 0 2.16672e-08 0.0021 2.16702e-08 0 2.17252e-08 0 2.17282e-08 0.0021 2.17312e-08 0 2.17862e-08 0 2.17892e-08 0.0021 2.17922e-08 0 2.18472e-08 0 2.18502e-08 0.0021 2.18532e-08 0 2.19082e-08 0 2.19112e-08 0.0021 2.19142e-08 0 2.19692e-08 0 2.19722e-08 0.0021 2.19752e-08 0 2.20302e-08 0 2.20332e-08 0.0021 2.20362e-08 0 2.20912e-08 0 2.20942e-08 0.0021 2.20972e-08 0 2.21522e-08 0 2.21552e-08 0.0021 2.21582e-08 0 2.22132e-08 0 2.22162e-08 0.0021 2.22192e-08 0 2.22742e-08 0 2.22772e-08 0.0021 2.22802e-08 0 2.23352e-08 0 2.23382e-08 0.0021 2.23412e-08 0 2.23962e-08 0 2.23992e-08 0.0021 2.24022e-08 0 2.24572e-08 0 2.24602e-08 0.0021 2.24632e-08 0 2.25182e-08 0 2.25212e-08 0.0021 2.25242e-08 0 2.25792e-08 0 2.25822e-08 0.0021 2.25852e-08 0 2.26402e-08 0 2.26432e-08 0.0021 2.26462e-08 0 2.27012e-08 0 2.27042e-08 0.0021 2.27072e-08 0 2.27622e-08 0 2.27652e-08 0.0021 2.27682e-08 0 2.28232e-08 0 2.28262e-08 0.0021 2.28292e-08 0 2.28842e-08 0 2.28872e-08 0.0021 2.28902e-08 0 2.29452e-08 0 2.29482e-08 0.0021 2.29512e-08 0 2.30062e-08 0 2.30092e-08 0.0021 2.30122e-08 0 2.30672e-08 0 2.30702e-08 0.0021 2.30732e-08 0 2.31282e-08 0 2.31312e-08 0.0021 2.31342e-08 0 2.31892e-08 0 2.31922e-08 0.0021 2.31952e-08 0 2.32502e-08 0 2.32532e-08 0.0021 2.32562e-08 0 2.33112e-08 0 2.33142e-08 0.0021 2.33172e-08 0 2.33722e-08 0 2.33752e-08 0.0021 2.33782e-08 0 2.34332e-08 0 2.34362e-08 0.0021 2.34392e-08 0 2.34942e-08 0 2.34972e-08 0.0021 2.35002e-08 0 2.35552e-08 0 2.35582e-08 0.0021 2.35612e-08 0 2.36162e-08 0 2.36192e-08 0.0021 2.36222e-08 0 2.36772e-08 0 2.36802e-08 0.0021 2.36832e-08 0 2.37382e-08 0 2.37412e-08 0.0021 2.37442e-08 0 2.37992e-08 0 2.38022e-08 0.0021 2.38052e-08 0 2.38602e-08 0 2.38632e-08 0.0021 2.38662e-08 0 2.39212e-08 0 2.39242e-08 0.0021 2.39272e-08 0 2.39822e-08 0 2.39852e-08 0.0021 2.39882e-08 0 2.40432e-08 0 2.40462e-08 0.0021 2.40492e-08 0 2.41042e-08 0 2.41072e-08 0.0021 2.41102e-08 0 2.41652e-08 0 2.41682e-08 0.0021 2.41712e-08 0 2.42262e-08 0 2.42292e-08 0.0021 2.42322e-08 0 2.42872e-08 0 2.42902e-08 0.0021 2.42932e-08 0)
IT01|T 0 T01  PWL(0 0 9.2e-12 0 1.22e-11 0.0021 1.52e-11 0 7.02e-11 0 7.32e-11 0.0021 7.62e-11 0 1.312e-10 0 1.342e-10 0.0021 1.372e-10 0 1.922e-10 0 1.952e-10 0.0021 1.982e-10 0 2.532e-10 0 2.562e-10 0.0021 2.592e-10 0 3.142e-10 0 3.172e-10 0.0021 3.202e-10 0 3.752e-10 0 3.782e-10 0.0021 3.812e-10 0 4.362e-10 0 4.392e-10 0.0021 4.422e-10 0 4.972e-10 0 5.002e-10 0.0021 5.032e-10 0 5.582e-10 0 5.612e-10 0.0021 5.642e-10 0 6.192e-10 0 6.222e-10 0.0021 6.252e-10 0 6.802e-10 0 6.832e-10 0.0021 6.862e-10 0 7.412e-10 0 7.442e-10 0.0021 7.472e-10 0 8.022e-10 0 8.052e-10 0.0021 8.082e-10 0 8.632e-10 0 8.662e-10 0.0021 8.692e-10 0 9.242e-10 0 9.272e-10 0.0021 9.302e-10 0 9.852e-10 0 9.882e-10 0.0021 9.912e-10 0 1.0462e-09 0 1.0492e-09 0.0021 1.0522e-09 0 1.1072e-09 0 1.1102e-09 0.0021 1.1132e-09 0 1.1682e-09 0 1.1712e-09 0.0021 1.1742e-09 0 1.2292e-09 0 1.2322e-09 0.0021 1.2352e-09 0 1.2902e-09 0 1.2932e-09 0.0021 1.2962e-09 0 1.3512e-09 0 1.3542e-09 0.0021 1.3572e-09 0 1.4122e-09 0 1.4152e-09 0.0021 1.4182e-09 0 1.4732e-09 0 1.4762e-09 0.0021 1.4792e-09 0 1.5342e-09 0 1.5372e-09 0.0021 1.5402e-09 0 1.5952e-09 0 1.5982e-09 0.0021 1.6012e-09 0 1.6562e-09 0 1.6592e-09 0.0021 1.6622e-09 0 1.7172e-09 0 1.7202e-09 0.0021 1.7232e-09 0 1.7782e-09 0 1.7812e-09 0.0021 1.7842e-09 0 1.8392e-09 0 1.8422e-09 0.0021 1.8452e-09 0 1.9002e-09 0 1.9032e-09 0.0021 1.9062e-09 0 1.9612e-09 0 1.9642e-09 0.0021 1.9672e-09 0 2.0222e-09 0 2.0252e-09 0.0021 2.0282e-09 0 2.0832e-09 0 2.0862e-09 0.0021 2.0892e-09 0 2.1442e-09 0 2.1472e-09 0.0021 2.1502e-09 0 2.2052e-09 0 2.2082e-09 0.0021 2.2112e-09 0 2.2662e-09 0 2.2692e-09 0.0021 2.2722e-09 0 2.3272e-09 0 2.3302e-09 0.0021 2.3332e-09 0 2.3882e-09 0 2.3912e-09 0.0021 2.3942e-09 0 2.4492e-09 0 2.4522e-09 0.0021 2.4552e-09 0 2.5102e-09 0 2.5132e-09 0.0021 2.5162e-09 0 2.5712e-09 0 2.5742e-09 0.0021 2.5772e-09 0 2.6322e-09 0 2.6352e-09 0.0021 2.6382e-09 0 2.6932e-09 0 2.6962e-09 0.0021 2.6992e-09 0 2.7542e-09 0 2.7572e-09 0.0021 2.7602e-09 0 2.8152e-09 0 2.8182e-09 0.0021 2.8212e-09 0 2.8762e-09 0 2.8792e-09 0.0021 2.8822e-09 0 2.9372e-09 0 2.9402e-09 0.0021 2.9432e-09 0 2.9982e-09 0 3.0012e-09 0.0021 3.0042e-09 0 3.0592e-09 0 3.0622e-09 0.0021 3.0652e-09 0 3.1202e-09 0 3.1232e-09 0.0021 3.1262e-09 0 3.1812e-09 0 3.1842e-09 0.0021 3.1872e-09 0 3.2422e-09 0 3.2452e-09 0.0021 3.2482e-09 0 3.3032e-09 0 3.3062e-09 0.0021 3.3092e-09 0 3.3642e-09 0 3.3672e-09 0.0021 3.3702e-09 0 3.4252e-09 0 3.4282e-09 0.0021 3.4312e-09 0 3.4862e-09 0 3.4892e-09 0.0021 3.4922e-09 0 3.5472e-09 0 3.5502e-09 0.0021 3.5532e-09 0 3.6082e-09 0 3.6112e-09 0.0021 3.6142e-09 0 3.6692e-09 0 3.6722e-09 0.0021 3.6752e-09 0 3.7302e-09 0 3.7332e-09 0.0021 3.7362e-09 0 3.7912e-09 0 3.7942e-09 0.0021 3.7972e-09 0 3.8522e-09 0 3.8552e-09 0.0021 3.8582e-09 0 3.9132e-09 0 3.9162e-09 0.0021 3.9192e-09 0 3.9742e-09 0 3.9772e-09 0.0021 3.9802e-09 0 4.0352e-09 0 4.0382e-09 0.0021 4.0412e-09 0 4.0962e-09 0 4.0992e-09 0.0021 4.1022e-09 0 4.1572e-09 0 4.1602e-09 0.0021 4.1632e-09 0 4.2182e-09 0 4.2212e-09 0.0021 4.2242e-09 0 4.2792e-09 0 4.2822e-09 0.0021 4.2852e-09 0 4.3402e-09 0 4.3432e-09 0.0021 4.3462e-09 0 4.4012e-09 0 4.4042e-09 0.0021 4.4072e-09 0 4.4622e-09 0 4.4652e-09 0.0021 4.4682e-09 0 4.5232e-09 0 4.5262e-09 0.0021 4.5292e-09 0 4.5842e-09 0 4.5872e-09 0.0021 4.5902e-09 0 4.6452e-09 0 4.6482e-09 0.0021 4.6512e-09 0 4.7062e-09 0 4.7092e-09 0.0021 4.7122e-09 0 4.7672e-09 0 4.7702e-09 0.0021 4.7732e-09 0 4.8282e-09 0 4.8312e-09 0.0021 4.8342e-09 0 4.8892e-09 0 4.8922e-09 0.0021 4.8952e-09 0 4.9502e-09 0 4.9532e-09 0.0021 4.9562e-09 0 5.0112e-09 0 5.0142e-09 0.0021 5.0172e-09 0 5.0722e-09 0 5.0752e-09 0.0021 5.0782e-09 0 5.1332e-09 0 5.1362e-09 0.0021 5.1392e-09 0 5.1942e-09 0 5.1972e-09 0.0021 5.2002e-09 0 5.2552e-09 0 5.2582e-09 0.0021 5.2612e-09 0 5.3162e-09 0 5.3192e-09 0.0021 5.3222e-09 0 5.3772e-09 0 5.3802e-09 0.0021 5.3832e-09 0 5.4382e-09 0 5.4412e-09 0.0021 5.4442e-09 0 5.4992e-09 0 5.5022e-09 0.0021 5.5052e-09 0 5.5602e-09 0 5.5632e-09 0.0021 5.5662e-09 0 5.6212e-09 0 5.6242e-09 0.0021 5.6272e-09 0 5.6822e-09 0 5.6852e-09 0.0021 5.6882e-09 0 5.7432e-09 0 5.7462e-09 0.0021 5.7492e-09 0 5.8042e-09 0 5.8072e-09 0.0021 5.8102e-09 0 5.8652e-09 0 5.8682e-09 0.0021 5.8712e-09 0 5.9262e-09 0 5.9292e-09 0.0021 5.9322e-09 0 5.9872e-09 0 5.9902e-09 0.0021 5.9932e-09 0 6.0482e-09 0 6.0512e-09 0.0021 6.0542e-09 0 6.1092e-09 0 6.1122e-09 0.0021 6.1152e-09 0 6.1702e-09 0 6.1732e-09 0.0021 6.1762e-09 0 6.2312e-09 0 6.2342e-09 0.0021 6.2372e-09 0 6.2922e-09 0 6.2952e-09 0.0021 6.2982e-09 0 6.3532e-09 0 6.3562e-09 0.0021 6.3592e-09 0 6.4142e-09 0 6.4172e-09 0.0021 6.4202e-09 0 6.4752e-09 0 6.4782e-09 0.0021 6.4812e-09 0 6.5362e-09 0 6.5392e-09 0.0021 6.5422e-09 0 6.5972e-09 0 6.6002e-09 0.0021 6.6032e-09 0 6.6582e-09 0 6.6612e-09 0.0021 6.6642e-09 0 6.7192e-09 0 6.7222e-09 0.0021 6.7252e-09 0 6.7802e-09 0 6.7832e-09 0.0021 6.7862e-09 0 6.8412e-09 0 6.8442e-09 0.0021 6.8472e-09 0 6.9022e-09 0 6.9052e-09 0.0021 6.9082e-09 0 6.9632e-09 0 6.9662e-09 0.0021 6.9692e-09 0 7.0242e-09 0 7.0272e-09 0.0021 7.0302e-09 0 7.0852e-09 0 7.0882e-09 0.0021 7.0912e-09 0 7.1462e-09 0 7.1492e-09 0.0021 7.1522e-09 0 7.2072e-09 0 7.2102e-09 0.0021 7.2132e-09 0 7.2682e-09 0 7.2712e-09 0.0021 7.2742e-09 0 7.3292e-09 0 7.3322e-09 0.0021 7.3352e-09 0 7.3902e-09 0 7.3932e-09 0.0021 7.3962e-09 0 7.4512e-09 0 7.4542e-09 0.0021 7.4572e-09 0 7.5122e-09 0 7.5152e-09 0.0021 7.5182e-09 0 7.5732e-09 0 7.5762e-09 0.0021 7.5792e-09 0 7.6342e-09 0 7.6372e-09 0.0021 7.6402e-09 0 7.6952e-09 0 7.6982e-09 0.0021 7.7012e-09 0 7.7562e-09 0 7.7592e-09 0.0021 7.7622e-09 0 7.8172e-09 0 7.8202e-09 0.0021 7.8232e-09 0 7.8782e-09 0 7.8812e-09 0.0021 7.8842e-09 0 7.9392e-09 0 7.9422e-09 0.0021 7.9452e-09 0 8.0002e-09 0 8.0032e-09 0.0021 8.0062e-09 0 8.0612e-09 0 8.0642e-09 0.0021 8.0672e-09 0 8.1222e-09 0 8.1252e-09 0.0021 8.1282e-09 0 8.1832e-09 0 8.1862e-09 0.0021 8.1892e-09 0 8.2442e-09 0 8.2472e-09 0.0021 8.2502e-09 0 8.3052e-09 0 8.3082e-09 0.0021 8.3112e-09 0 8.3662e-09 0 8.3692e-09 0.0021 8.3722e-09 0 8.4272e-09 0 8.4302e-09 0.0021 8.4332e-09 0 8.4882e-09 0 8.4912e-09 0.0021 8.4942e-09 0 8.5492e-09 0 8.5522e-09 0.0021 8.5552e-09 0 8.6102e-09 0 8.6132e-09 0.0021 8.6162e-09 0 8.6712e-09 0 8.6742e-09 0.0021 8.6772e-09 0 8.7322e-09 0 8.7352e-09 0.0021 8.7382e-09 0 8.7932e-09 0 8.7962e-09 0.0021 8.7992e-09 0 8.8542e-09 0 8.8572e-09 0.0021 8.8602e-09 0 8.9152e-09 0 8.9182e-09 0.0021 8.9212e-09 0 8.9762e-09 0 8.9792e-09 0.0021 8.9822e-09 0 9.0372e-09 0 9.0402e-09 0.0021 9.0432e-09 0 9.0982e-09 0 9.1012e-09 0.0021 9.1042e-09 0 9.1592e-09 0 9.1622e-09 0.0021 9.1652e-09 0 9.2202e-09 0 9.2232e-09 0.0021 9.2262e-09 0 9.2812e-09 0 9.2842e-09 0.0021 9.2872e-09 0 9.3422e-09 0 9.3452e-09 0.0021 9.3482e-09 0 9.4032e-09 0 9.4062e-09 0.0021 9.4092e-09 0 9.4642e-09 0 9.4672e-09 0.0021 9.4702e-09 0 9.5252e-09 0 9.5282e-09 0.0021 9.5312e-09 0 9.5862e-09 0 9.5892e-09 0.0021 9.5922e-09 0 9.6472e-09 0 9.6502e-09 0.0021 9.6532e-09 0 9.7082e-09 0 9.7112e-09 0.0021 9.7142e-09 0 9.7692e-09 0 9.7722e-09 0.0021 9.7752e-09 0 9.8302e-09 0 9.8332e-09 0.0021 9.8362e-09 0 9.8912e-09 0 9.8942e-09 0.0021 9.8972e-09 0 9.9522e-09 0 9.9552e-09 0.0021 9.9582e-09 0 1.00132e-08 0 1.00162e-08 0.0021 1.00192e-08 0 1.00742e-08 0 1.00772e-08 0.0021 1.00802e-08 0 1.01352e-08 0 1.01382e-08 0.0021 1.01412e-08 0 1.01962e-08 0 1.01992e-08 0.0021 1.02022e-08 0 1.02572e-08 0 1.02602e-08 0.0021 1.02632e-08 0 1.03182e-08 0 1.03212e-08 0.0021 1.03242e-08 0 1.03792e-08 0 1.03822e-08 0.0021 1.03852e-08 0 1.04402e-08 0 1.04432e-08 0.0021 1.04462e-08 0 1.05012e-08 0 1.05042e-08 0.0021 1.05072e-08 0 1.05622e-08 0 1.05652e-08 0.0021 1.05682e-08 0 1.06232e-08 0 1.06262e-08 0.0021 1.06292e-08 0 1.06842e-08 0 1.06872e-08 0.0021 1.06902e-08 0 1.07452e-08 0 1.07482e-08 0.0021 1.07512e-08 0 1.08062e-08 0 1.08092e-08 0.0021 1.08122e-08 0 1.08672e-08 0 1.08702e-08 0.0021 1.08732e-08 0 1.09282e-08 0 1.09312e-08 0.0021 1.09342e-08 0 1.09892e-08 0 1.09922e-08 0.0021 1.09952e-08 0 1.10502e-08 0 1.10532e-08 0.0021 1.10562e-08 0 1.11112e-08 0 1.11142e-08 0.0021 1.11172e-08 0 1.11722e-08 0 1.11752e-08 0.0021 1.11782e-08 0 1.12332e-08 0 1.12362e-08 0.0021 1.12392e-08 0 1.12942e-08 0 1.12972e-08 0.0021 1.13002e-08 0 1.13552e-08 0 1.13582e-08 0.0021 1.13612e-08 0 1.14162e-08 0 1.14192e-08 0.0021 1.14222e-08 0 1.14772e-08 0 1.14802e-08 0.0021 1.14832e-08 0 1.15382e-08 0 1.15412e-08 0.0021 1.15442e-08 0 1.15992e-08 0 1.16022e-08 0.0021 1.16052e-08 0 1.16602e-08 0 1.16632e-08 0.0021 1.16662e-08 0 1.17212e-08 0 1.17242e-08 0.0021 1.17272e-08 0 1.17822e-08 0 1.17852e-08 0.0021 1.17882e-08 0 1.18432e-08 0 1.18462e-08 0.0021 1.18492e-08 0 1.19042e-08 0 1.19072e-08 0.0021 1.19102e-08 0 1.19652e-08 0 1.19682e-08 0.0021 1.19712e-08 0 1.20262e-08 0 1.20292e-08 0.0021 1.20322e-08 0 1.20872e-08 0 1.20902e-08 0.0021 1.20932e-08 0 1.21482e-08 0 1.21512e-08 0.0021 1.21542e-08 0 1.22092e-08 0 1.22122e-08 0.0021 1.22152e-08 0 1.22702e-08 0 1.22732e-08 0.0021 1.22762e-08 0 1.23312e-08 0 1.23342e-08 0.0021 1.23372e-08 0 1.23922e-08 0 1.23952e-08 0.0021 1.23982e-08 0 1.24532e-08 0 1.24562e-08 0.0021 1.24592e-08 0 1.25142e-08 0 1.25172e-08 0.0021 1.25202e-08 0 1.25752e-08 0 1.25782e-08 0.0021 1.25812e-08 0 1.26362e-08 0 1.26392e-08 0.0021 1.26422e-08 0 1.26972e-08 0 1.27002e-08 0.0021 1.27032e-08 0 1.27582e-08 0 1.27612e-08 0.0021 1.27642e-08 0 1.28192e-08 0 1.28222e-08 0.0021 1.28252e-08 0 1.28802e-08 0 1.28832e-08 0.0021 1.28862e-08 0 1.29412e-08 0 1.29442e-08 0.0021 1.29472e-08 0 1.30022e-08 0 1.30052e-08 0.0021 1.30082e-08 0 1.30632e-08 0 1.30662e-08 0.0021 1.30692e-08 0 1.31242e-08 0 1.31272e-08 0.0021 1.31302e-08 0 1.31852e-08 0 1.31882e-08 0.0021 1.31912e-08 0 1.32462e-08 0 1.32492e-08 0.0021 1.32522e-08 0 1.33072e-08 0 1.33102e-08 0.0021 1.33132e-08 0 1.33682e-08 0 1.33712e-08 0.0021 1.33742e-08 0 1.34292e-08 0 1.34322e-08 0.0021 1.34352e-08 0 1.34902e-08 0 1.34932e-08 0.0021 1.34962e-08 0 1.35512e-08 0 1.35542e-08 0.0021 1.35572e-08 0 1.36122e-08 0 1.36152e-08 0.0021 1.36182e-08 0 1.36732e-08 0 1.36762e-08 0.0021 1.36792e-08 0 1.37342e-08 0 1.37372e-08 0.0021 1.37402e-08 0 1.37952e-08 0 1.37982e-08 0.0021 1.38012e-08 0 1.38562e-08 0 1.38592e-08 0.0021 1.38622e-08 0 1.39172e-08 0 1.39202e-08 0.0021 1.39232e-08 0 1.39782e-08 0 1.39812e-08 0.0021 1.39842e-08 0 1.40392e-08 0 1.40422e-08 0.0021 1.40452e-08 0 1.41002e-08 0 1.41032e-08 0.0021 1.41062e-08 0 1.41612e-08 0 1.41642e-08 0.0021 1.41672e-08 0 1.42222e-08 0 1.42252e-08 0.0021 1.42282e-08 0 1.42832e-08 0 1.42862e-08 0.0021 1.42892e-08 0 1.43442e-08 0 1.43472e-08 0.0021 1.43502e-08 0 1.44052e-08 0 1.44082e-08 0.0021 1.44112e-08 0 1.44662e-08 0 1.44692e-08 0.0021 1.44722e-08 0 1.45272e-08 0 1.45302e-08 0.0021 1.45332e-08 0 1.45882e-08 0 1.45912e-08 0.0021 1.45942e-08 0 1.46492e-08 0 1.46522e-08 0.0021 1.46552e-08 0 1.47102e-08 0 1.47132e-08 0.0021 1.47162e-08 0 1.47712e-08 0 1.47742e-08 0.0021 1.47772e-08 0 1.48322e-08 0 1.48352e-08 0.0021 1.48382e-08 0 1.48932e-08 0 1.48962e-08 0.0021 1.48992e-08 0 1.49542e-08 0 1.49572e-08 0.0021 1.49602e-08 0 1.50152e-08 0 1.50182e-08 0.0021 1.50212e-08 0 1.50762e-08 0 1.50792e-08 0.0021 1.50822e-08 0 1.51372e-08 0 1.51402e-08 0.0021 1.51432e-08 0 1.51982e-08 0 1.52012e-08 0.0021 1.52042e-08 0 1.52592e-08 0 1.52622e-08 0.0021 1.52652e-08 0 1.53202e-08 0 1.53232e-08 0.0021 1.53262e-08 0 1.53812e-08 0 1.53842e-08 0.0021 1.53872e-08 0 1.54422e-08 0 1.54452e-08 0.0021 1.54482e-08 0 1.55032e-08 0 1.55062e-08 0.0021 1.55092e-08 0 1.55642e-08 0 1.55672e-08 0.0021 1.55702e-08 0 1.56252e-08 0 1.56282e-08 0.0021 1.56312e-08 0 1.56862e-08 0 1.56892e-08 0.0021 1.56922e-08 0 1.57472e-08 0 1.57502e-08 0.0021 1.57532e-08 0 1.58082e-08 0 1.58112e-08 0.0021 1.58142e-08 0 1.58692e-08 0 1.58722e-08 0.0021 1.58752e-08 0 1.59302e-08 0 1.59332e-08 0.0021 1.59362e-08 0 1.59912e-08 0 1.59942e-08 0.0021 1.59972e-08 0 1.60522e-08 0 1.60552e-08 0.0021 1.60582e-08 0 1.61132e-08 0 1.61162e-08 0.0021 1.61192e-08 0 1.61742e-08 0 1.61772e-08 0.0021 1.61802e-08 0 1.62352e-08 0 1.62382e-08 0.0021 1.62412e-08 0 1.62962e-08 0 1.62992e-08 0.0021 1.63022e-08 0 1.63572e-08 0 1.63602e-08 0.0021 1.63632e-08 0 1.64182e-08 0 1.64212e-08 0.0021 1.64242e-08 0 1.64792e-08 0 1.64822e-08 0.0021 1.64852e-08 0 1.65402e-08 0 1.65432e-08 0.0021 1.65462e-08 0 1.66012e-08 0 1.66042e-08 0.0021 1.66072e-08 0 1.66622e-08 0 1.66652e-08 0.0021 1.66682e-08 0 1.67232e-08 0 1.67262e-08 0.0021 1.67292e-08 0 1.67842e-08 0 1.67872e-08 0.0021 1.67902e-08 0 1.68452e-08 0 1.68482e-08 0.0021 1.68512e-08 0 1.69062e-08 0 1.69092e-08 0.0021 1.69122e-08 0 1.69672e-08 0 1.69702e-08 0.0021 1.69732e-08 0 1.70282e-08 0 1.70312e-08 0.0021 1.70342e-08 0 1.70892e-08 0 1.70922e-08 0.0021 1.70952e-08 0 1.71502e-08 0 1.71532e-08 0.0021 1.71562e-08 0 1.72112e-08 0 1.72142e-08 0.0021 1.72172e-08 0 1.72722e-08 0 1.72752e-08 0.0021 1.72782e-08 0 1.73332e-08 0 1.73362e-08 0.0021 1.73392e-08 0 1.73942e-08 0 1.73972e-08 0.0021 1.74002e-08 0 1.74552e-08 0 1.74582e-08 0.0021 1.74612e-08 0 1.75162e-08 0 1.75192e-08 0.0021 1.75222e-08 0 1.75772e-08 0 1.75802e-08 0.0021 1.75832e-08 0 1.76382e-08 0 1.76412e-08 0.0021 1.76442e-08 0 1.76992e-08 0 1.77022e-08 0.0021 1.77052e-08 0 1.77602e-08 0 1.77632e-08 0.0021 1.77662e-08 0 1.78212e-08 0 1.78242e-08 0.0021 1.78272e-08 0 1.78822e-08 0 1.78852e-08 0.0021 1.78882e-08 0 1.79432e-08 0 1.79462e-08 0.0021 1.79492e-08 0 1.80042e-08 0 1.80072e-08 0.0021 1.80102e-08 0 1.80652e-08 0 1.80682e-08 0.0021 1.80712e-08 0 1.81262e-08 0 1.81292e-08 0.0021 1.81322e-08 0 1.81872e-08 0 1.81902e-08 0.0021 1.81932e-08 0 1.82482e-08 0 1.82512e-08 0.0021 1.82542e-08 0 1.83092e-08 0 1.83122e-08 0.0021 1.83152e-08 0 1.83702e-08 0 1.83732e-08 0.0021 1.83762e-08 0 1.84312e-08 0 1.84342e-08 0.0021 1.84372e-08 0 1.84922e-08 0 1.84952e-08 0.0021 1.84982e-08 0 1.85532e-08 0 1.85562e-08 0.0021 1.85592e-08 0 1.86142e-08 0 1.86172e-08 0.0021 1.86202e-08 0 1.86752e-08 0 1.86782e-08 0.0021 1.86812e-08 0 1.87362e-08 0 1.87392e-08 0.0021 1.87422e-08 0 1.87972e-08 0 1.88002e-08 0.0021 1.88032e-08 0 1.88582e-08 0 1.88612e-08 0.0021 1.88642e-08 0 1.89192e-08 0 1.89222e-08 0.0021 1.89252e-08 0 1.89802e-08 0 1.89832e-08 0.0021 1.89862e-08 0 1.90412e-08 0 1.90442e-08 0.0021 1.90472e-08 0 1.91022e-08 0 1.91052e-08 0.0021 1.91082e-08 0 1.91632e-08 0 1.91662e-08 0.0021 1.91692e-08 0 1.92242e-08 0 1.92272e-08 0.0021 1.92302e-08 0 1.92852e-08 0 1.92882e-08 0.0021 1.92912e-08 0 1.93462e-08 0 1.93492e-08 0.0021 1.93522e-08 0 1.94072e-08 0 1.94102e-08 0.0021 1.94132e-08 0 1.94682e-08 0 1.94712e-08 0.0021 1.94742e-08 0 1.95292e-08 0 1.95322e-08 0.0021 1.95352e-08 0 1.95902e-08 0 1.95932e-08 0.0021 1.95962e-08 0 1.96512e-08 0 1.96542e-08 0.0021 1.96572e-08 0 1.97122e-08 0 1.97152e-08 0.0021 1.97182e-08 0 1.97732e-08 0 1.97762e-08 0.0021 1.97792e-08 0 1.98342e-08 0 1.98372e-08 0.0021 1.98402e-08 0 1.98952e-08 0 1.98982e-08 0.0021 1.99012e-08 0 1.99562e-08 0 1.99592e-08 0.0021 1.99622e-08 0 2.00172e-08 0 2.00202e-08 0.0021 2.00232e-08 0 2.00782e-08 0 2.00812e-08 0.0021 2.00842e-08 0 2.01392e-08 0 2.01422e-08 0.0021 2.01452e-08 0 2.02002e-08 0 2.02032e-08 0.0021 2.02062e-08 0 2.02612e-08 0 2.02642e-08 0.0021 2.02672e-08 0 2.03222e-08 0 2.03252e-08 0.0021 2.03282e-08 0 2.03832e-08 0 2.03862e-08 0.0021 2.03892e-08 0 2.04442e-08 0 2.04472e-08 0.0021 2.04502e-08 0 2.05052e-08 0 2.05082e-08 0.0021 2.05112e-08 0 2.05662e-08 0 2.05692e-08 0.0021 2.05722e-08 0 2.06272e-08 0 2.06302e-08 0.0021 2.06332e-08 0 2.06882e-08 0 2.06912e-08 0.0021 2.06942e-08 0 2.07492e-08 0 2.07522e-08 0.0021 2.07552e-08 0 2.08102e-08 0 2.08132e-08 0.0021 2.08162e-08 0 2.08712e-08 0 2.08742e-08 0.0021 2.08772e-08 0 2.09322e-08 0 2.09352e-08 0.0021 2.09382e-08 0 2.09932e-08 0 2.09962e-08 0.0021 2.09992e-08 0 2.10542e-08 0 2.10572e-08 0.0021 2.10602e-08 0 2.11152e-08 0 2.11182e-08 0.0021 2.11212e-08 0 2.11762e-08 0 2.11792e-08 0.0021 2.11822e-08 0 2.12372e-08 0 2.12402e-08 0.0021 2.12432e-08 0 2.12982e-08 0 2.13012e-08 0.0021 2.13042e-08 0 2.13592e-08 0 2.13622e-08 0.0021 2.13652e-08 0 2.14202e-08 0 2.14232e-08 0.0021 2.14262e-08 0 2.14812e-08 0 2.14842e-08 0.0021 2.14872e-08 0 2.15422e-08 0 2.15452e-08 0.0021 2.15482e-08 0 2.16032e-08 0 2.16062e-08 0.0021 2.16092e-08 0 2.16642e-08 0 2.16672e-08 0.0021 2.16702e-08 0 2.17252e-08 0 2.17282e-08 0.0021 2.17312e-08 0 2.17862e-08 0 2.17892e-08 0.0021 2.17922e-08 0 2.18472e-08 0 2.18502e-08 0.0021 2.18532e-08 0 2.19082e-08 0 2.19112e-08 0.0021 2.19142e-08 0 2.19692e-08 0 2.19722e-08 0.0021 2.19752e-08 0 2.20302e-08 0 2.20332e-08 0.0021 2.20362e-08 0 2.20912e-08 0 2.20942e-08 0.0021 2.20972e-08 0 2.21522e-08 0 2.21552e-08 0.0021 2.21582e-08 0 2.22132e-08 0 2.22162e-08 0.0021 2.22192e-08 0 2.22742e-08 0 2.22772e-08 0.0021 2.22802e-08 0 2.23352e-08 0 2.23382e-08 0.0021 2.23412e-08 0 2.23962e-08 0 2.23992e-08 0.0021 2.24022e-08 0 2.24572e-08 0 2.24602e-08 0.0021 2.24632e-08 0 2.25182e-08 0 2.25212e-08 0.0021 2.25242e-08 0 2.25792e-08 0 2.25822e-08 0.0021 2.25852e-08 0 2.26402e-08 0 2.26432e-08 0.0021 2.26462e-08 0 2.27012e-08 0 2.27042e-08 0.0021 2.27072e-08 0 2.27622e-08 0 2.27652e-08 0.0021 2.27682e-08 0 2.28232e-08 0 2.28262e-08 0.0021 2.28292e-08 0 2.28842e-08 0 2.28872e-08 0.0021 2.28902e-08 0 2.29452e-08 0 2.29482e-08 0.0021 2.29512e-08 0 2.30062e-08 0 2.30092e-08 0.0021 2.30122e-08 0 2.30672e-08 0 2.30702e-08 0.0021 2.30732e-08 0 2.31282e-08 0 2.31312e-08 0.0021 2.31342e-08 0 2.31892e-08 0 2.31922e-08 0.0021 2.31952e-08 0 2.32502e-08 0 2.32532e-08 0.0021 2.32562e-08 0 2.33112e-08 0 2.33142e-08 0.0021 2.33172e-08 0 2.33722e-08 0 2.33752e-08 0.0021 2.33782e-08 0 2.34332e-08 0 2.34362e-08 0.0021 2.34392e-08 0 2.34942e-08 0 2.34972e-08 0.0021 2.35002e-08 0 2.35552e-08 0 2.35582e-08 0.0021 2.35612e-08 0 2.36162e-08 0 2.36192e-08 0.0021 2.36222e-08 0 2.36772e-08 0 2.36802e-08 0.0021 2.36832e-08 0 2.37382e-08 0 2.37412e-08 0.0021 2.37442e-08 0 2.37992e-08 0 2.38022e-08 0.0021 2.38052e-08 0 2.38602e-08 0 2.38632e-08 0.0021 2.38662e-08 0 2.39212e-08 0 2.39242e-08 0.0021 2.39272e-08 0 2.39822e-08 0 2.39852e-08 0.0021 2.39882e-08 0 2.40432e-08 0 2.40462e-08 0.0021 2.40492e-08 0 2.41042e-08 0 2.41072e-08 0.0021 2.41102e-08 0 2.41652e-08 0 2.41682e-08 0.0021 2.41712e-08 0 2.42262e-08 0 2.42292e-08 0.0021 2.42322e-08 0 2.42872e-08 0 2.42902e-08 0.0021 2.42932e-08 0)
IT02|T 0 T02  PWL(0 0 9.2e-12 0 1.22e-11 0.0021 1.52e-11 0 7.02e-11 0 7.32e-11 0.0021 7.62e-11 0 1.312e-10 0 1.342e-10 0.0021 1.372e-10 0 1.922e-10 0 1.952e-10 0.0021 1.982e-10 0 2.532e-10 0 2.562e-10 0.0021 2.592e-10 0 3.142e-10 0 3.172e-10 0.0021 3.202e-10 0 3.752e-10 0 3.782e-10 0.0021 3.812e-10 0 4.362e-10 0 4.392e-10 0.0021 4.422e-10 0 4.972e-10 0 5.002e-10 0.0021 5.032e-10 0 5.582e-10 0 5.612e-10 0.0021 5.642e-10 0 6.192e-10 0 6.222e-10 0.0021 6.252e-10 0 6.802e-10 0 6.832e-10 0.0021 6.862e-10 0 7.412e-10 0 7.442e-10 0.0021 7.472e-10 0 8.022e-10 0 8.052e-10 0.0021 8.082e-10 0 8.632e-10 0 8.662e-10 0.0021 8.692e-10 0 9.242e-10 0 9.272e-10 0.0021 9.302e-10 0 9.852e-10 0 9.882e-10 0.0021 9.912e-10 0 1.0462e-09 0 1.0492e-09 0.0021 1.0522e-09 0 1.1072e-09 0 1.1102e-09 0.0021 1.1132e-09 0 1.1682e-09 0 1.1712e-09 0.0021 1.1742e-09 0 1.2292e-09 0 1.2322e-09 0.0021 1.2352e-09 0 1.2902e-09 0 1.2932e-09 0.0021 1.2962e-09 0 1.3512e-09 0 1.3542e-09 0.0021 1.3572e-09 0 1.4122e-09 0 1.4152e-09 0.0021 1.4182e-09 0 1.4732e-09 0 1.4762e-09 0.0021 1.4792e-09 0 1.5342e-09 0 1.5372e-09 0.0021 1.5402e-09 0 1.5952e-09 0 1.5982e-09 0.0021 1.6012e-09 0 1.6562e-09 0 1.6592e-09 0.0021 1.6622e-09 0 1.7172e-09 0 1.7202e-09 0.0021 1.7232e-09 0 1.7782e-09 0 1.7812e-09 0.0021 1.7842e-09 0 1.8392e-09 0 1.8422e-09 0.0021 1.8452e-09 0 1.9002e-09 0 1.9032e-09 0.0021 1.9062e-09 0 1.9612e-09 0 1.9642e-09 0.0021 1.9672e-09 0 2.0222e-09 0 2.0252e-09 0.0021 2.0282e-09 0 2.0832e-09 0 2.0862e-09 0.0021 2.0892e-09 0 2.1442e-09 0 2.1472e-09 0.0021 2.1502e-09 0 2.2052e-09 0 2.2082e-09 0.0021 2.2112e-09 0 2.2662e-09 0 2.2692e-09 0.0021 2.2722e-09 0 2.3272e-09 0 2.3302e-09 0.0021 2.3332e-09 0 2.3882e-09 0 2.3912e-09 0.0021 2.3942e-09 0 2.4492e-09 0 2.4522e-09 0.0021 2.4552e-09 0 2.5102e-09 0 2.5132e-09 0.0021 2.5162e-09 0 2.5712e-09 0 2.5742e-09 0.0021 2.5772e-09 0 2.6322e-09 0 2.6352e-09 0.0021 2.6382e-09 0 2.6932e-09 0 2.6962e-09 0.0021 2.6992e-09 0 2.7542e-09 0 2.7572e-09 0.0021 2.7602e-09 0 2.8152e-09 0 2.8182e-09 0.0021 2.8212e-09 0 2.8762e-09 0 2.8792e-09 0.0021 2.8822e-09 0 2.9372e-09 0 2.9402e-09 0.0021 2.9432e-09 0 2.9982e-09 0 3.0012e-09 0.0021 3.0042e-09 0 3.0592e-09 0 3.0622e-09 0.0021 3.0652e-09 0 3.1202e-09 0 3.1232e-09 0.0021 3.1262e-09 0 3.1812e-09 0 3.1842e-09 0.0021 3.1872e-09 0 3.2422e-09 0 3.2452e-09 0.0021 3.2482e-09 0 3.3032e-09 0 3.3062e-09 0.0021 3.3092e-09 0 3.3642e-09 0 3.3672e-09 0.0021 3.3702e-09 0 3.4252e-09 0 3.4282e-09 0.0021 3.4312e-09 0 3.4862e-09 0 3.4892e-09 0.0021 3.4922e-09 0 3.5472e-09 0 3.5502e-09 0.0021 3.5532e-09 0 3.6082e-09 0 3.6112e-09 0.0021 3.6142e-09 0 3.6692e-09 0 3.6722e-09 0.0021 3.6752e-09 0 3.7302e-09 0 3.7332e-09 0.0021 3.7362e-09 0 3.7912e-09 0 3.7942e-09 0.0021 3.7972e-09 0 3.8522e-09 0 3.8552e-09 0.0021 3.8582e-09 0 3.9132e-09 0 3.9162e-09 0.0021 3.9192e-09 0 3.9742e-09 0 3.9772e-09 0.0021 3.9802e-09 0 4.0352e-09 0 4.0382e-09 0.0021 4.0412e-09 0 4.0962e-09 0 4.0992e-09 0.0021 4.1022e-09 0 4.1572e-09 0 4.1602e-09 0.0021 4.1632e-09 0 4.2182e-09 0 4.2212e-09 0.0021 4.2242e-09 0 4.2792e-09 0 4.2822e-09 0.0021 4.2852e-09 0 4.3402e-09 0 4.3432e-09 0.0021 4.3462e-09 0 4.4012e-09 0 4.4042e-09 0.0021 4.4072e-09 0 4.4622e-09 0 4.4652e-09 0.0021 4.4682e-09 0 4.5232e-09 0 4.5262e-09 0.0021 4.5292e-09 0 4.5842e-09 0 4.5872e-09 0.0021 4.5902e-09 0 4.6452e-09 0 4.6482e-09 0.0021 4.6512e-09 0 4.7062e-09 0 4.7092e-09 0.0021 4.7122e-09 0 4.7672e-09 0 4.7702e-09 0.0021 4.7732e-09 0 4.8282e-09 0 4.8312e-09 0.0021 4.8342e-09 0 4.8892e-09 0 4.8922e-09 0.0021 4.8952e-09 0 4.9502e-09 0 4.9532e-09 0.0021 4.9562e-09 0 5.0112e-09 0 5.0142e-09 0.0021 5.0172e-09 0 5.0722e-09 0 5.0752e-09 0.0021 5.0782e-09 0 5.1332e-09 0 5.1362e-09 0.0021 5.1392e-09 0 5.1942e-09 0 5.1972e-09 0.0021 5.2002e-09 0 5.2552e-09 0 5.2582e-09 0.0021 5.2612e-09 0 5.3162e-09 0 5.3192e-09 0.0021 5.3222e-09 0 5.3772e-09 0 5.3802e-09 0.0021 5.3832e-09 0 5.4382e-09 0 5.4412e-09 0.0021 5.4442e-09 0 5.4992e-09 0 5.5022e-09 0.0021 5.5052e-09 0 5.5602e-09 0 5.5632e-09 0.0021 5.5662e-09 0 5.6212e-09 0 5.6242e-09 0.0021 5.6272e-09 0 5.6822e-09 0 5.6852e-09 0.0021 5.6882e-09 0 5.7432e-09 0 5.7462e-09 0.0021 5.7492e-09 0 5.8042e-09 0 5.8072e-09 0.0021 5.8102e-09 0 5.8652e-09 0 5.8682e-09 0.0021 5.8712e-09 0 5.9262e-09 0 5.9292e-09 0.0021 5.9322e-09 0 5.9872e-09 0 5.9902e-09 0.0021 5.9932e-09 0 6.0482e-09 0 6.0512e-09 0.0021 6.0542e-09 0 6.1092e-09 0 6.1122e-09 0.0021 6.1152e-09 0 6.1702e-09 0 6.1732e-09 0.0021 6.1762e-09 0 6.2312e-09 0 6.2342e-09 0.0021 6.2372e-09 0 6.2922e-09 0 6.2952e-09 0.0021 6.2982e-09 0 6.3532e-09 0 6.3562e-09 0.0021 6.3592e-09 0 6.4142e-09 0 6.4172e-09 0.0021 6.4202e-09 0 6.4752e-09 0 6.4782e-09 0.0021 6.4812e-09 0 6.5362e-09 0 6.5392e-09 0.0021 6.5422e-09 0 6.5972e-09 0 6.6002e-09 0.0021 6.6032e-09 0 6.6582e-09 0 6.6612e-09 0.0021 6.6642e-09 0 6.7192e-09 0 6.7222e-09 0.0021 6.7252e-09 0 6.7802e-09 0 6.7832e-09 0.0021 6.7862e-09 0 6.8412e-09 0 6.8442e-09 0.0021 6.8472e-09 0 6.9022e-09 0 6.9052e-09 0.0021 6.9082e-09 0 6.9632e-09 0 6.9662e-09 0.0021 6.9692e-09 0 7.0242e-09 0 7.0272e-09 0.0021 7.0302e-09 0 7.0852e-09 0 7.0882e-09 0.0021 7.0912e-09 0 7.1462e-09 0 7.1492e-09 0.0021 7.1522e-09 0 7.2072e-09 0 7.2102e-09 0.0021 7.2132e-09 0 7.2682e-09 0 7.2712e-09 0.0021 7.2742e-09 0 7.3292e-09 0 7.3322e-09 0.0021 7.3352e-09 0 7.3902e-09 0 7.3932e-09 0.0021 7.3962e-09 0 7.4512e-09 0 7.4542e-09 0.0021 7.4572e-09 0 7.5122e-09 0 7.5152e-09 0.0021 7.5182e-09 0 7.5732e-09 0 7.5762e-09 0.0021 7.5792e-09 0 7.6342e-09 0 7.6372e-09 0.0021 7.6402e-09 0 7.6952e-09 0 7.6982e-09 0.0021 7.7012e-09 0 7.7562e-09 0 7.7592e-09 0.0021 7.7622e-09 0 7.8172e-09 0 7.8202e-09 0.0021 7.8232e-09 0 7.8782e-09 0 7.8812e-09 0.0021 7.8842e-09 0 7.9392e-09 0 7.9422e-09 0.0021 7.9452e-09 0 8.0002e-09 0 8.0032e-09 0.0021 8.0062e-09 0 8.0612e-09 0 8.0642e-09 0.0021 8.0672e-09 0 8.1222e-09 0 8.1252e-09 0.0021 8.1282e-09 0 8.1832e-09 0 8.1862e-09 0.0021 8.1892e-09 0 8.2442e-09 0 8.2472e-09 0.0021 8.2502e-09 0 8.3052e-09 0 8.3082e-09 0.0021 8.3112e-09 0 8.3662e-09 0 8.3692e-09 0.0021 8.3722e-09 0 8.4272e-09 0 8.4302e-09 0.0021 8.4332e-09 0 8.4882e-09 0 8.4912e-09 0.0021 8.4942e-09 0 8.5492e-09 0 8.5522e-09 0.0021 8.5552e-09 0 8.6102e-09 0 8.6132e-09 0.0021 8.6162e-09 0 8.6712e-09 0 8.6742e-09 0.0021 8.6772e-09 0 8.7322e-09 0 8.7352e-09 0.0021 8.7382e-09 0 8.7932e-09 0 8.7962e-09 0.0021 8.7992e-09 0 8.8542e-09 0 8.8572e-09 0.0021 8.8602e-09 0 8.9152e-09 0 8.9182e-09 0.0021 8.9212e-09 0 8.9762e-09 0 8.9792e-09 0.0021 8.9822e-09 0 9.0372e-09 0 9.0402e-09 0.0021 9.0432e-09 0 9.0982e-09 0 9.1012e-09 0.0021 9.1042e-09 0 9.1592e-09 0 9.1622e-09 0.0021 9.1652e-09 0 9.2202e-09 0 9.2232e-09 0.0021 9.2262e-09 0 9.2812e-09 0 9.2842e-09 0.0021 9.2872e-09 0 9.3422e-09 0 9.3452e-09 0.0021 9.3482e-09 0 9.4032e-09 0 9.4062e-09 0.0021 9.4092e-09 0 9.4642e-09 0 9.4672e-09 0.0021 9.4702e-09 0 9.5252e-09 0 9.5282e-09 0.0021 9.5312e-09 0 9.5862e-09 0 9.5892e-09 0.0021 9.5922e-09 0 9.6472e-09 0 9.6502e-09 0.0021 9.6532e-09 0 9.7082e-09 0 9.7112e-09 0.0021 9.7142e-09 0 9.7692e-09 0 9.7722e-09 0.0021 9.7752e-09 0 9.8302e-09 0 9.8332e-09 0.0021 9.8362e-09 0 9.8912e-09 0 9.8942e-09 0.0021 9.8972e-09 0 9.9522e-09 0 9.9552e-09 0.0021 9.9582e-09 0 1.00132e-08 0 1.00162e-08 0.0021 1.00192e-08 0 1.00742e-08 0 1.00772e-08 0.0021 1.00802e-08 0 1.01352e-08 0 1.01382e-08 0.0021 1.01412e-08 0 1.01962e-08 0 1.01992e-08 0.0021 1.02022e-08 0 1.02572e-08 0 1.02602e-08 0.0021 1.02632e-08 0 1.03182e-08 0 1.03212e-08 0.0021 1.03242e-08 0 1.03792e-08 0 1.03822e-08 0.0021 1.03852e-08 0 1.04402e-08 0 1.04432e-08 0.0021 1.04462e-08 0 1.05012e-08 0 1.05042e-08 0.0021 1.05072e-08 0 1.05622e-08 0 1.05652e-08 0.0021 1.05682e-08 0 1.06232e-08 0 1.06262e-08 0.0021 1.06292e-08 0 1.06842e-08 0 1.06872e-08 0.0021 1.06902e-08 0 1.07452e-08 0 1.07482e-08 0.0021 1.07512e-08 0 1.08062e-08 0 1.08092e-08 0.0021 1.08122e-08 0 1.08672e-08 0 1.08702e-08 0.0021 1.08732e-08 0 1.09282e-08 0 1.09312e-08 0.0021 1.09342e-08 0 1.09892e-08 0 1.09922e-08 0.0021 1.09952e-08 0 1.10502e-08 0 1.10532e-08 0.0021 1.10562e-08 0 1.11112e-08 0 1.11142e-08 0.0021 1.11172e-08 0 1.11722e-08 0 1.11752e-08 0.0021 1.11782e-08 0 1.12332e-08 0 1.12362e-08 0.0021 1.12392e-08 0 1.12942e-08 0 1.12972e-08 0.0021 1.13002e-08 0 1.13552e-08 0 1.13582e-08 0.0021 1.13612e-08 0 1.14162e-08 0 1.14192e-08 0.0021 1.14222e-08 0 1.14772e-08 0 1.14802e-08 0.0021 1.14832e-08 0 1.15382e-08 0 1.15412e-08 0.0021 1.15442e-08 0 1.15992e-08 0 1.16022e-08 0.0021 1.16052e-08 0 1.16602e-08 0 1.16632e-08 0.0021 1.16662e-08 0 1.17212e-08 0 1.17242e-08 0.0021 1.17272e-08 0 1.17822e-08 0 1.17852e-08 0.0021 1.17882e-08 0 1.18432e-08 0 1.18462e-08 0.0021 1.18492e-08 0 1.19042e-08 0 1.19072e-08 0.0021 1.19102e-08 0 1.19652e-08 0 1.19682e-08 0.0021 1.19712e-08 0 1.20262e-08 0 1.20292e-08 0.0021 1.20322e-08 0 1.20872e-08 0 1.20902e-08 0.0021 1.20932e-08 0 1.21482e-08 0 1.21512e-08 0.0021 1.21542e-08 0 1.22092e-08 0 1.22122e-08 0.0021 1.22152e-08 0 1.22702e-08 0 1.22732e-08 0.0021 1.22762e-08 0 1.23312e-08 0 1.23342e-08 0.0021 1.23372e-08 0 1.23922e-08 0 1.23952e-08 0.0021 1.23982e-08 0 1.24532e-08 0 1.24562e-08 0.0021 1.24592e-08 0 1.25142e-08 0 1.25172e-08 0.0021 1.25202e-08 0 1.25752e-08 0 1.25782e-08 0.0021 1.25812e-08 0 1.26362e-08 0 1.26392e-08 0.0021 1.26422e-08 0 1.26972e-08 0 1.27002e-08 0.0021 1.27032e-08 0 1.27582e-08 0 1.27612e-08 0.0021 1.27642e-08 0 1.28192e-08 0 1.28222e-08 0.0021 1.28252e-08 0 1.28802e-08 0 1.28832e-08 0.0021 1.28862e-08 0 1.29412e-08 0 1.29442e-08 0.0021 1.29472e-08 0 1.30022e-08 0 1.30052e-08 0.0021 1.30082e-08 0 1.30632e-08 0 1.30662e-08 0.0021 1.30692e-08 0 1.31242e-08 0 1.31272e-08 0.0021 1.31302e-08 0 1.31852e-08 0 1.31882e-08 0.0021 1.31912e-08 0 1.32462e-08 0 1.32492e-08 0.0021 1.32522e-08 0 1.33072e-08 0 1.33102e-08 0.0021 1.33132e-08 0 1.33682e-08 0 1.33712e-08 0.0021 1.33742e-08 0 1.34292e-08 0 1.34322e-08 0.0021 1.34352e-08 0 1.34902e-08 0 1.34932e-08 0.0021 1.34962e-08 0 1.35512e-08 0 1.35542e-08 0.0021 1.35572e-08 0 1.36122e-08 0 1.36152e-08 0.0021 1.36182e-08 0 1.36732e-08 0 1.36762e-08 0.0021 1.36792e-08 0 1.37342e-08 0 1.37372e-08 0.0021 1.37402e-08 0 1.37952e-08 0 1.37982e-08 0.0021 1.38012e-08 0 1.38562e-08 0 1.38592e-08 0.0021 1.38622e-08 0 1.39172e-08 0 1.39202e-08 0.0021 1.39232e-08 0 1.39782e-08 0 1.39812e-08 0.0021 1.39842e-08 0 1.40392e-08 0 1.40422e-08 0.0021 1.40452e-08 0 1.41002e-08 0 1.41032e-08 0.0021 1.41062e-08 0 1.41612e-08 0 1.41642e-08 0.0021 1.41672e-08 0 1.42222e-08 0 1.42252e-08 0.0021 1.42282e-08 0 1.42832e-08 0 1.42862e-08 0.0021 1.42892e-08 0 1.43442e-08 0 1.43472e-08 0.0021 1.43502e-08 0 1.44052e-08 0 1.44082e-08 0.0021 1.44112e-08 0 1.44662e-08 0 1.44692e-08 0.0021 1.44722e-08 0 1.45272e-08 0 1.45302e-08 0.0021 1.45332e-08 0 1.45882e-08 0 1.45912e-08 0.0021 1.45942e-08 0 1.46492e-08 0 1.46522e-08 0.0021 1.46552e-08 0 1.47102e-08 0 1.47132e-08 0.0021 1.47162e-08 0 1.47712e-08 0 1.47742e-08 0.0021 1.47772e-08 0 1.48322e-08 0 1.48352e-08 0.0021 1.48382e-08 0 1.48932e-08 0 1.48962e-08 0.0021 1.48992e-08 0 1.49542e-08 0 1.49572e-08 0.0021 1.49602e-08 0 1.50152e-08 0 1.50182e-08 0.0021 1.50212e-08 0 1.50762e-08 0 1.50792e-08 0.0021 1.50822e-08 0 1.51372e-08 0 1.51402e-08 0.0021 1.51432e-08 0 1.51982e-08 0 1.52012e-08 0.0021 1.52042e-08 0 1.52592e-08 0 1.52622e-08 0.0021 1.52652e-08 0 1.53202e-08 0 1.53232e-08 0.0021 1.53262e-08 0 1.53812e-08 0 1.53842e-08 0.0021 1.53872e-08 0 1.54422e-08 0 1.54452e-08 0.0021 1.54482e-08 0 1.55032e-08 0 1.55062e-08 0.0021 1.55092e-08 0 1.55642e-08 0 1.55672e-08 0.0021 1.55702e-08 0 1.56252e-08 0 1.56282e-08 0.0021 1.56312e-08 0 1.56862e-08 0 1.56892e-08 0.0021 1.56922e-08 0 1.57472e-08 0 1.57502e-08 0.0021 1.57532e-08 0 1.58082e-08 0 1.58112e-08 0.0021 1.58142e-08 0 1.58692e-08 0 1.58722e-08 0.0021 1.58752e-08 0 1.59302e-08 0 1.59332e-08 0.0021 1.59362e-08 0 1.59912e-08 0 1.59942e-08 0.0021 1.59972e-08 0 1.60522e-08 0 1.60552e-08 0.0021 1.60582e-08 0 1.61132e-08 0 1.61162e-08 0.0021 1.61192e-08 0 1.61742e-08 0 1.61772e-08 0.0021 1.61802e-08 0 1.62352e-08 0 1.62382e-08 0.0021 1.62412e-08 0 1.62962e-08 0 1.62992e-08 0.0021 1.63022e-08 0 1.63572e-08 0 1.63602e-08 0.0021 1.63632e-08 0 1.64182e-08 0 1.64212e-08 0.0021 1.64242e-08 0 1.64792e-08 0 1.64822e-08 0.0021 1.64852e-08 0 1.65402e-08 0 1.65432e-08 0.0021 1.65462e-08 0 1.66012e-08 0 1.66042e-08 0.0021 1.66072e-08 0 1.66622e-08 0 1.66652e-08 0.0021 1.66682e-08 0 1.67232e-08 0 1.67262e-08 0.0021 1.67292e-08 0 1.67842e-08 0 1.67872e-08 0.0021 1.67902e-08 0 1.68452e-08 0 1.68482e-08 0.0021 1.68512e-08 0 1.69062e-08 0 1.69092e-08 0.0021 1.69122e-08 0 1.69672e-08 0 1.69702e-08 0.0021 1.69732e-08 0 1.70282e-08 0 1.70312e-08 0.0021 1.70342e-08 0 1.70892e-08 0 1.70922e-08 0.0021 1.70952e-08 0 1.71502e-08 0 1.71532e-08 0.0021 1.71562e-08 0 1.72112e-08 0 1.72142e-08 0.0021 1.72172e-08 0 1.72722e-08 0 1.72752e-08 0.0021 1.72782e-08 0 1.73332e-08 0 1.73362e-08 0.0021 1.73392e-08 0 1.73942e-08 0 1.73972e-08 0.0021 1.74002e-08 0 1.74552e-08 0 1.74582e-08 0.0021 1.74612e-08 0 1.75162e-08 0 1.75192e-08 0.0021 1.75222e-08 0 1.75772e-08 0 1.75802e-08 0.0021 1.75832e-08 0 1.76382e-08 0 1.76412e-08 0.0021 1.76442e-08 0 1.76992e-08 0 1.77022e-08 0.0021 1.77052e-08 0 1.77602e-08 0 1.77632e-08 0.0021 1.77662e-08 0 1.78212e-08 0 1.78242e-08 0.0021 1.78272e-08 0 1.78822e-08 0 1.78852e-08 0.0021 1.78882e-08 0 1.79432e-08 0 1.79462e-08 0.0021 1.79492e-08 0 1.80042e-08 0 1.80072e-08 0.0021 1.80102e-08 0 1.80652e-08 0 1.80682e-08 0.0021 1.80712e-08 0 1.81262e-08 0 1.81292e-08 0.0021 1.81322e-08 0 1.81872e-08 0 1.81902e-08 0.0021 1.81932e-08 0 1.82482e-08 0 1.82512e-08 0.0021 1.82542e-08 0 1.83092e-08 0 1.83122e-08 0.0021 1.83152e-08 0 1.83702e-08 0 1.83732e-08 0.0021 1.83762e-08 0 1.84312e-08 0 1.84342e-08 0.0021 1.84372e-08 0 1.84922e-08 0 1.84952e-08 0.0021 1.84982e-08 0 1.85532e-08 0 1.85562e-08 0.0021 1.85592e-08 0 1.86142e-08 0 1.86172e-08 0.0021 1.86202e-08 0 1.86752e-08 0 1.86782e-08 0.0021 1.86812e-08 0 1.87362e-08 0 1.87392e-08 0.0021 1.87422e-08 0 1.87972e-08 0 1.88002e-08 0.0021 1.88032e-08 0 1.88582e-08 0 1.88612e-08 0.0021 1.88642e-08 0 1.89192e-08 0 1.89222e-08 0.0021 1.89252e-08 0 1.89802e-08 0 1.89832e-08 0.0021 1.89862e-08 0 1.90412e-08 0 1.90442e-08 0.0021 1.90472e-08 0 1.91022e-08 0 1.91052e-08 0.0021 1.91082e-08 0 1.91632e-08 0 1.91662e-08 0.0021 1.91692e-08 0 1.92242e-08 0 1.92272e-08 0.0021 1.92302e-08 0 1.92852e-08 0 1.92882e-08 0.0021 1.92912e-08 0 1.93462e-08 0 1.93492e-08 0.0021 1.93522e-08 0 1.94072e-08 0 1.94102e-08 0.0021 1.94132e-08 0 1.94682e-08 0 1.94712e-08 0.0021 1.94742e-08 0 1.95292e-08 0 1.95322e-08 0.0021 1.95352e-08 0 1.95902e-08 0 1.95932e-08 0.0021 1.95962e-08 0 1.96512e-08 0 1.96542e-08 0.0021 1.96572e-08 0 1.97122e-08 0 1.97152e-08 0.0021 1.97182e-08 0 1.97732e-08 0 1.97762e-08 0.0021 1.97792e-08 0 1.98342e-08 0 1.98372e-08 0.0021 1.98402e-08 0 1.98952e-08 0 1.98982e-08 0.0021 1.99012e-08 0 1.99562e-08 0 1.99592e-08 0.0021 1.99622e-08 0 2.00172e-08 0 2.00202e-08 0.0021 2.00232e-08 0 2.00782e-08 0 2.00812e-08 0.0021 2.00842e-08 0 2.01392e-08 0 2.01422e-08 0.0021 2.01452e-08 0 2.02002e-08 0 2.02032e-08 0.0021 2.02062e-08 0 2.02612e-08 0 2.02642e-08 0.0021 2.02672e-08 0 2.03222e-08 0 2.03252e-08 0.0021 2.03282e-08 0 2.03832e-08 0 2.03862e-08 0.0021 2.03892e-08 0 2.04442e-08 0 2.04472e-08 0.0021 2.04502e-08 0 2.05052e-08 0 2.05082e-08 0.0021 2.05112e-08 0 2.05662e-08 0 2.05692e-08 0.0021 2.05722e-08 0 2.06272e-08 0 2.06302e-08 0.0021 2.06332e-08 0 2.06882e-08 0 2.06912e-08 0.0021 2.06942e-08 0 2.07492e-08 0 2.07522e-08 0.0021 2.07552e-08 0 2.08102e-08 0 2.08132e-08 0.0021 2.08162e-08 0 2.08712e-08 0 2.08742e-08 0.0021 2.08772e-08 0 2.09322e-08 0 2.09352e-08 0.0021 2.09382e-08 0 2.09932e-08 0 2.09962e-08 0.0021 2.09992e-08 0 2.10542e-08 0 2.10572e-08 0.0021 2.10602e-08 0 2.11152e-08 0 2.11182e-08 0.0021 2.11212e-08 0 2.11762e-08 0 2.11792e-08 0.0021 2.11822e-08 0 2.12372e-08 0 2.12402e-08 0.0021 2.12432e-08 0 2.12982e-08 0 2.13012e-08 0.0021 2.13042e-08 0 2.13592e-08 0 2.13622e-08 0.0021 2.13652e-08 0 2.14202e-08 0 2.14232e-08 0.0021 2.14262e-08 0 2.14812e-08 0 2.14842e-08 0.0021 2.14872e-08 0 2.15422e-08 0 2.15452e-08 0.0021 2.15482e-08 0 2.16032e-08 0 2.16062e-08 0.0021 2.16092e-08 0 2.16642e-08 0 2.16672e-08 0.0021 2.16702e-08 0 2.17252e-08 0 2.17282e-08 0.0021 2.17312e-08 0 2.17862e-08 0 2.17892e-08 0.0021 2.17922e-08 0 2.18472e-08 0 2.18502e-08 0.0021 2.18532e-08 0 2.19082e-08 0 2.19112e-08 0.0021 2.19142e-08 0 2.19692e-08 0 2.19722e-08 0.0021 2.19752e-08 0 2.20302e-08 0 2.20332e-08 0.0021 2.20362e-08 0 2.20912e-08 0 2.20942e-08 0.0021 2.20972e-08 0 2.21522e-08 0 2.21552e-08 0.0021 2.21582e-08 0 2.22132e-08 0 2.22162e-08 0.0021 2.22192e-08 0 2.22742e-08 0 2.22772e-08 0.0021 2.22802e-08 0 2.23352e-08 0 2.23382e-08 0.0021 2.23412e-08 0 2.23962e-08 0 2.23992e-08 0.0021 2.24022e-08 0 2.24572e-08 0 2.24602e-08 0.0021 2.24632e-08 0 2.25182e-08 0 2.25212e-08 0.0021 2.25242e-08 0 2.25792e-08 0 2.25822e-08 0.0021 2.25852e-08 0 2.26402e-08 0 2.26432e-08 0.0021 2.26462e-08 0 2.27012e-08 0 2.27042e-08 0.0021 2.27072e-08 0 2.27622e-08 0 2.27652e-08 0.0021 2.27682e-08 0 2.28232e-08 0 2.28262e-08 0.0021 2.28292e-08 0 2.28842e-08 0 2.28872e-08 0.0021 2.28902e-08 0 2.29452e-08 0 2.29482e-08 0.0021 2.29512e-08 0 2.30062e-08 0 2.30092e-08 0.0021 2.30122e-08 0 2.30672e-08 0 2.30702e-08 0.0021 2.30732e-08 0 2.31282e-08 0 2.31312e-08 0.0021 2.31342e-08 0 2.31892e-08 0 2.31922e-08 0.0021 2.31952e-08 0 2.32502e-08 0 2.32532e-08 0.0021 2.32562e-08 0 2.33112e-08 0 2.33142e-08 0.0021 2.33172e-08 0 2.33722e-08 0 2.33752e-08 0.0021 2.33782e-08 0 2.34332e-08 0 2.34362e-08 0.0021 2.34392e-08 0 2.34942e-08 0 2.34972e-08 0.0021 2.35002e-08 0 2.35552e-08 0 2.35582e-08 0.0021 2.35612e-08 0 2.36162e-08 0 2.36192e-08 0.0021 2.36222e-08 0 2.36772e-08 0 2.36802e-08 0.0021 2.36832e-08 0 2.37382e-08 0 2.37412e-08 0.0021 2.37442e-08 0 2.37992e-08 0 2.38022e-08 0.0021 2.38052e-08 0 2.38602e-08 0 2.38632e-08 0.0021 2.38662e-08 0 2.39212e-08 0 2.39242e-08 0.0021 2.39272e-08 0 2.39822e-08 0 2.39852e-08 0.0021 2.39882e-08 0 2.40432e-08 0 2.40462e-08 0.0021 2.40492e-08 0 2.41042e-08 0 2.41072e-08 0.0021 2.41102e-08 0 2.41652e-08 0 2.41682e-08 0.0021 2.41712e-08 0 2.42262e-08 0 2.42292e-08 0.0021 2.42322e-08 0 2.42872e-08 0 2.42902e-08 0.0021 2.42932e-08 0)
IT03|T 0 T03  PWL(0 0 9.2e-12 0 1.22e-11 0.0021 1.52e-11 0 7.02e-11 0 7.32e-11 0.0021 7.62e-11 0 1.312e-10 0 1.342e-10 0.0021 1.372e-10 0 1.922e-10 0 1.952e-10 0.0021 1.982e-10 0 2.532e-10 0 2.562e-10 0.0021 2.592e-10 0 3.142e-10 0 3.172e-10 0.0021 3.202e-10 0 3.752e-10 0 3.782e-10 0.0021 3.812e-10 0 4.362e-10 0 4.392e-10 0.0021 4.422e-10 0 4.972e-10 0 5.002e-10 0.0021 5.032e-10 0 5.582e-10 0 5.612e-10 0.0021 5.642e-10 0 6.192e-10 0 6.222e-10 0.0021 6.252e-10 0 6.802e-10 0 6.832e-10 0.0021 6.862e-10 0 7.412e-10 0 7.442e-10 0.0021 7.472e-10 0 8.022e-10 0 8.052e-10 0.0021 8.082e-10 0 8.632e-10 0 8.662e-10 0.0021 8.692e-10 0 9.242e-10 0 9.272e-10 0.0021 9.302e-10 0 9.852e-10 0 9.882e-10 0.0021 9.912e-10 0 1.0462e-09 0 1.0492e-09 0.0021 1.0522e-09 0 1.1072e-09 0 1.1102e-09 0.0021 1.1132e-09 0 1.1682e-09 0 1.1712e-09 0.0021 1.1742e-09 0 1.2292e-09 0 1.2322e-09 0.0021 1.2352e-09 0 1.2902e-09 0 1.2932e-09 0.0021 1.2962e-09 0 1.3512e-09 0 1.3542e-09 0.0021 1.3572e-09 0 1.4122e-09 0 1.4152e-09 0.0021 1.4182e-09 0 1.4732e-09 0 1.4762e-09 0.0021 1.4792e-09 0 1.5342e-09 0 1.5372e-09 0.0021 1.5402e-09 0 1.5952e-09 0 1.5982e-09 0.0021 1.6012e-09 0 1.6562e-09 0 1.6592e-09 0.0021 1.6622e-09 0 1.7172e-09 0 1.7202e-09 0.0021 1.7232e-09 0 1.7782e-09 0 1.7812e-09 0.0021 1.7842e-09 0 1.8392e-09 0 1.8422e-09 0.0021 1.8452e-09 0 1.9002e-09 0 1.9032e-09 0.0021 1.9062e-09 0 1.9612e-09 0 1.9642e-09 0.0021 1.9672e-09 0 2.0222e-09 0 2.0252e-09 0.0021 2.0282e-09 0 2.0832e-09 0 2.0862e-09 0.0021 2.0892e-09 0 2.1442e-09 0 2.1472e-09 0.0021 2.1502e-09 0 2.2052e-09 0 2.2082e-09 0.0021 2.2112e-09 0 2.2662e-09 0 2.2692e-09 0.0021 2.2722e-09 0 2.3272e-09 0 2.3302e-09 0.0021 2.3332e-09 0 2.3882e-09 0 2.3912e-09 0.0021 2.3942e-09 0 2.4492e-09 0 2.4522e-09 0.0021 2.4552e-09 0 2.5102e-09 0 2.5132e-09 0.0021 2.5162e-09 0 2.5712e-09 0 2.5742e-09 0.0021 2.5772e-09 0 2.6322e-09 0 2.6352e-09 0.0021 2.6382e-09 0 2.6932e-09 0 2.6962e-09 0.0021 2.6992e-09 0 2.7542e-09 0 2.7572e-09 0.0021 2.7602e-09 0 2.8152e-09 0 2.8182e-09 0.0021 2.8212e-09 0 2.8762e-09 0 2.8792e-09 0.0021 2.8822e-09 0 2.9372e-09 0 2.9402e-09 0.0021 2.9432e-09 0 2.9982e-09 0 3.0012e-09 0.0021 3.0042e-09 0 3.0592e-09 0 3.0622e-09 0.0021 3.0652e-09 0 3.1202e-09 0 3.1232e-09 0.0021 3.1262e-09 0 3.1812e-09 0 3.1842e-09 0.0021 3.1872e-09 0 3.2422e-09 0 3.2452e-09 0.0021 3.2482e-09 0 3.3032e-09 0 3.3062e-09 0.0021 3.3092e-09 0 3.3642e-09 0 3.3672e-09 0.0021 3.3702e-09 0 3.4252e-09 0 3.4282e-09 0.0021 3.4312e-09 0 3.4862e-09 0 3.4892e-09 0.0021 3.4922e-09 0 3.5472e-09 0 3.5502e-09 0.0021 3.5532e-09 0 3.6082e-09 0 3.6112e-09 0.0021 3.6142e-09 0 3.6692e-09 0 3.6722e-09 0.0021 3.6752e-09 0 3.7302e-09 0 3.7332e-09 0.0021 3.7362e-09 0 3.7912e-09 0 3.7942e-09 0.0021 3.7972e-09 0 3.8522e-09 0 3.8552e-09 0.0021 3.8582e-09 0 3.9132e-09 0 3.9162e-09 0.0021 3.9192e-09 0 3.9742e-09 0 3.9772e-09 0.0021 3.9802e-09 0 4.0352e-09 0 4.0382e-09 0.0021 4.0412e-09 0 4.0962e-09 0 4.0992e-09 0.0021 4.1022e-09 0 4.1572e-09 0 4.1602e-09 0.0021 4.1632e-09 0 4.2182e-09 0 4.2212e-09 0.0021 4.2242e-09 0 4.2792e-09 0 4.2822e-09 0.0021 4.2852e-09 0 4.3402e-09 0 4.3432e-09 0.0021 4.3462e-09 0 4.4012e-09 0 4.4042e-09 0.0021 4.4072e-09 0 4.4622e-09 0 4.4652e-09 0.0021 4.4682e-09 0 4.5232e-09 0 4.5262e-09 0.0021 4.5292e-09 0 4.5842e-09 0 4.5872e-09 0.0021 4.5902e-09 0 4.6452e-09 0 4.6482e-09 0.0021 4.6512e-09 0 4.7062e-09 0 4.7092e-09 0.0021 4.7122e-09 0 4.7672e-09 0 4.7702e-09 0.0021 4.7732e-09 0 4.8282e-09 0 4.8312e-09 0.0021 4.8342e-09 0 4.8892e-09 0 4.8922e-09 0.0021 4.8952e-09 0 4.9502e-09 0 4.9532e-09 0.0021 4.9562e-09 0 5.0112e-09 0 5.0142e-09 0.0021 5.0172e-09 0 5.0722e-09 0 5.0752e-09 0.0021 5.0782e-09 0 5.1332e-09 0 5.1362e-09 0.0021 5.1392e-09 0 5.1942e-09 0 5.1972e-09 0.0021 5.2002e-09 0 5.2552e-09 0 5.2582e-09 0.0021 5.2612e-09 0 5.3162e-09 0 5.3192e-09 0.0021 5.3222e-09 0 5.3772e-09 0 5.3802e-09 0.0021 5.3832e-09 0 5.4382e-09 0 5.4412e-09 0.0021 5.4442e-09 0 5.4992e-09 0 5.5022e-09 0.0021 5.5052e-09 0 5.5602e-09 0 5.5632e-09 0.0021 5.5662e-09 0 5.6212e-09 0 5.6242e-09 0.0021 5.6272e-09 0 5.6822e-09 0 5.6852e-09 0.0021 5.6882e-09 0 5.7432e-09 0 5.7462e-09 0.0021 5.7492e-09 0 5.8042e-09 0 5.8072e-09 0.0021 5.8102e-09 0 5.8652e-09 0 5.8682e-09 0.0021 5.8712e-09 0 5.9262e-09 0 5.9292e-09 0.0021 5.9322e-09 0 5.9872e-09 0 5.9902e-09 0.0021 5.9932e-09 0 6.0482e-09 0 6.0512e-09 0.0021 6.0542e-09 0 6.1092e-09 0 6.1122e-09 0.0021 6.1152e-09 0 6.1702e-09 0 6.1732e-09 0.0021 6.1762e-09 0 6.2312e-09 0 6.2342e-09 0.0021 6.2372e-09 0 6.2922e-09 0 6.2952e-09 0.0021 6.2982e-09 0 6.3532e-09 0 6.3562e-09 0.0021 6.3592e-09 0 6.4142e-09 0 6.4172e-09 0.0021 6.4202e-09 0 6.4752e-09 0 6.4782e-09 0.0021 6.4812e-09 0 6.5362e-09 0 6.5392e-09 0.0021 6.5422e-09 0 6.5972e-09 0 6.6002e-09 0.0021 6.6032e-09 0 6.6582e-09 0 6.6612e-09 0.0021 6.6642e-09 0 6.7192e-09 0 6.7222e-09 0.0021 6.7252e-09 0 6.7802e-09 0 6.7832e-09 0.0021 6.7862e-09 0 6.8412e-09 0 6.8442e-09 0.0021 6.8472e-09 0 6.9022e-09 0 6.9052e-09 0.0021 6.9082e-09 0 6.9632e-09 0 6.9662e-09 0.0021 6.9692e-09 0 7.0242e-09 0 7.0272e-09 0.0021 7.0302e-09 0 7.0852e-09 0 7.0882e-09 0.0021 7.0912e-09 0 7.1462e-09 0 7.1492e-09 0.0021 7.1522e-09 0 7.2072e-09 0 7.2102e-09 0.0021 7.2132e-09 0 7.2682e-09 0 7.2712e-09 0.0021 7.2742e-09 0 7.3292e-09 0 7.3322e-09 0.0021 7.3352e-09 0 7.3902e-09 0 7.3932e-09 0.0021 7.3962e-09 0 7.4512e-09 0 7.4542e-09 0.0021 7.4572e-09 0 7.5122e-09 0 7.5152e-09 0.0021 7.5182e-09 0 7.5732e-09 0 7.5762e-09 0.0021 7.5792e-09 0 7.6342e-09 0 7.6372e-09 0.0021 7.6402e-09 0 7.6952e-09 0 7.6982e-09 0.0021 7.7012e-09 0 7.7562e-09 0 7.7592e-09 0.0021 7.7622e-09 0 7.8172e-09 0 7.8202e-09 0.0021 7.8232e-09 0 7.8782e-09 0 7.8812e-09 0.0021 7.8842e-09 0 7.9392e-09 0 7.9422e-09 0.0021 7.9452e-09 0 8.0002e-09 0 8.0032e-09 0.0021 8.0062e-09 0 8.0612e-09 0 8.0642e-09 0.0021 8.0672e-09 0 8.1222e-09 0 8.1252e-09 0.0021 8.1282e-09 0 8.1832e-09 0 8.1862e-09 0.0021 8.1892e-09 0 8.2442e-09 0 8.2472e-09 0.0021 8.2502e-09 0 8.3052e-09 0 8.3082e-09 0.0021 8.3112e-09 0 8.3662e-09 0 8.3692e-09 0.0021 8.3722e-09 0 8.4272e-09 0 8.4302e-09 0.0021 8.4332e-09 0 8.4882e-09 0 8.4912e-09 0.0021 8.4942e-09 0 8.5492e-09 0 8.5522e-09 0.0021 8.5552e-09 0 8.6102e-09 0 8.6132e-09 0.0021 8.6162e-09 0 8.6712e-09 0 8.6742e-09 0.0021 8.6772e-09 0 8.7322e-09 0 8.7352e-09 0.0021 8.7382e-09 0 8.7932e-09 0 8.7962e-09 0.0021 8.7992e-09 0 8.8542e-09 0 8.8572e-09 0.0021 8.8602e-09 0 8.9152e-09 0 8.9182e-09 0.0021 8.9212e-09 0 8.9762e-09 0 8.9792e-09 0.0021 8.9822e-09 0 9.0372e-09 0 9.0402e-09 0.0021 9.0432e-09 0 9.0982e-09 0 9.1012e-09 0.0021 9.1042e-09 0 9.1592e-09 0 9.1622e-09 0.0021 9.1652e-09 0 9.2202e-09 0 9.2232e-09 0.0021 9.2262e-09 0 9.2812e-09 0 9.2842e-09 0.0021 9.2872e-09 0 9.3422e-09 0 9.3452e-09 0.0021 9.3482e-09 0 9.4032e-09 0 9.4062e-09 0.0021 9.4092e-09 0 9.4642e-09 0 9.4672e-09 0.0021 9.4702e-09 0 9.5252e-09 0 9.5282e-09 0.0021 9.5312e-09 0 9.5862e-09 0 9.5892e-09 0.0021 9.5922e-09 0 9.6472e-09 0 9.6502e-09 0.0021 9.6532e-09 0 9.7082e-09 0 9.7112e-09 0.0021 9.7142e-09 0 9.7692e-09 0 9.7722e-09 0.0021 9.7752e-09 0 9.8302e-09 0 9.8332e-09 0.0021 9.8362e-09 0 9.8912e-09 0 9.8942e-09 0.0021 9.8972e-09 0 9.9522e-09 0 9.9552e-09 0.0021 9.9582e-09 0 1.00132e-08 0 1.00162e-08 0.0021 1.00192e-08 0 1.00742e-08 0 1.00772e-08 0.0021 1.00802e-08 0 1.01352e-08 0 1.01382e-08 0.0021 1.01412e-08 0 1.01962e-08 0 1.01992e-08 0.0021 1.02022e-08 0 1.02572e-08 0 1.02602e-08 0.0021 1.02632e-08 0 1.03182e-08 0 1.03212e-08 0.0021 1.03242e-08 0 1.03792e-08 0 1.03822e-08 0.0021 1.03852e-08 0 1.04402e-08 0 1.04432e-08 0.0021 1.04462e-08 0 1.05012e-08 0 1.05042e-08 0.0021 1.05072e-08 0 1.05622e-08 0 1.05652e-08 0.0021 1.05682e-08 0 1.06232e-08 0 1.06262e-08 0.0021 1.06292e-08 0 1.06842e-08 0 1.06872e-08 0.0021 1.06902e-08 0 1.07452e-08 0 1.07482e-08 0.0021 1.07512e-08 0 1.08062e-08 0 1.08092e-08 0.0021 1.08122e-08 0 1.08672e-08 0 1.08702e-08 0.0021 1.08732e-08 0 1.09282e-08 0 1.09312e-08 0.0021 1.09342e-08 0 1.09892e-08 0 1.09922e-08 0.0021 1.09952e-08 0 1.10502e-08 0 1.10532e-08 0.0021 1.10562e-08 0 1.11112e-08 0 1.11142e-08 0.0021 1.11172e-08 0 1.11722e-08 0 1.11752e-08 0.0021 1.11782e-08 0 1.12332e-08 0 1.12362e-08 0.0021 1.12392e-08 0 1.12942e-08 0 1.12972e-08 0.0021 1.13002e-08 0 1.13552e-08 0 1.13582e-08 0.0021 1.13612e-08 0 1.14162e-08 0 1.14192e-08 0.0021 1.14222e-08 0 1.14772e-08 0 1.14802e-08 0.0021 1.14832e-08 0 1.15382e-08 0 1.15412e-08 0.0021 1.15442e-08 0 1.15992e-08 0 1.16022e-08 0.0021 1.16052e-08 0 1.16602e-08 0 1.16632e-08 0.0021 1.16662e-08 0 1.17212e-08 0 1.17242e-08 0.0021 1.17272e-08 0 1.17822e-08 0 1.17852e-08 0.0021 1.17882e-08 0 1.18432e-08 0 1.18462e-08 0.0021 1.18492e-08 0 1.19042e-08 0 1.19072e-08 0.0021 1.19102e-08 0 1.19652e-08 0 1.19682e-08 0.0021 1.19712e-08 0 1.20262e-08 0 1.20292e-08 0.0021 1.20322e-08 0 1.20872e-08 0 1.20902e-08 0.0021 1.20932e-08 0 1.21482e-08 0 1.21512e-08 0.0021 1.21542e-08 0 1.22092e-08 0 1.22122e-08 0.0021 1.22152e-08 0 1.22702e-08 0 1.22732e-08 0.0021 1.22762e-08 0 1.23312e-08 0 1.23342e-08 0.0021 1.23372e-08 0 1.23922e-08 0 1.23952e-08 0.0021 1.23982e-08 0 1.24532e-08 0 1.24562e-08 0.0021 1.24592e-08 0 1.25142e-08 0 1.25172e-08 0.0021 1.25202e-08 0 1.25752e-08 0 1.25782e-08 0.0021 1.25812e-08 0 1.26362e-08 0 1.26392e-08 0.0021 1.26422e-08 0 1.26972e-08 0 1.27002e-08 0.0021 1.27032e-08 0 1.27582e-08 0 1.27612e-08 0.0021 1.27642e-08 0 1.28192e-08 0 1.28222e-08 0.0021 1.28252e-08 0 1.28802e-08 0 1.28832e-08 0.0021 1.28862e-08 0 1.29412e-08 0 1.29442e-08 0.0021 1.29472e-08 0 1.30022e-08 0 1.30052e-08 0.0021 1.30082e-08 0 1.30632e-08 0 1.30662e-08 0.0021 1.30692e-08 0 1.31242e-08 0 1.31272e-08 0.0021 1.31302e-08 0 1.31852e-08 0 1.31882e-08 0.0021 1.31912e-08 0 1.32462e-08 0 1.32492e-08 0.0021 1.32522e-08 0 1.33072e-08 0 1.33102e-08 0.0021 1.33132e-08 0 1.33682e-08 0 1.33712e-08 0.0021 1.33742e-08 0 1.34292e-08 0 1.34322e-08 0.0021 1.34352e-08 0 1.34902e-08 0 1.34932e-08 0.0021 1.34962e-08 0 1.35512e-08 0 1.35542e-08 0.0021 1.35572e-08 0 1.36122e-08 0 1.36152e-08 0.0021 1.36182e-08 0 1.36732e-08 0 1.36762e-08 0.0021 1.36792e-08 0 1.37342e-08 0 1.37372e-08 0.0021 1.37402e-08 0 1.37952e-08 0 1.37982e-08 0.0021 1.38012e-08 0 1.38562e-08 0 1.38592e-08 0.0021 1.38622e-08 0 1.39172e-08 0 1.39202e-08 0.0021 1.39232e-08 0 1.39782e-08 0 1.39812e-08 0.0021 1.39842e-08 0 1.40392e-08 0 1.40422e-08 0.0021 1.40452e-08 0 1.41002e-08 0 1.41032e-08 0.0021 1.41062e-08 0 1.41612e-08 0 1.41642e-08 0.0021 1.41672e-08 0 1.42222e-08 0 1.42252e-08 0.0021 1.42282e-08 0 1.42832e-08 0 1.42862e-08 0.0021 1.42892e-08 0 1.43442e-08 0 1.43472e-08 0.0021 1.43502e-08 0 1.44052e-08 0 1.44082e-08 0.0021 1.44112e-08 0 1.44662e-08 0 1.44692e-08 0.0021 1.44722e-08 0 1.45272e-08 0 1.45302e-08 0.0021 1.45332e-08 0 1.45882e-08 0 1.45912e-08 0.0021 1.45942e-08 0 1.46492e-08 0 1.46522e-08 0.0021 1.46552e-08 0 1.47102e-08 0 1.47132e-08 0.0021 1.47162e-08 0 1.47712e-08 0 1.47742e-08 0.0021 1.47772e-08 0 1.48322e-08 0 1.48352e-08 0.0021 1.48382e-08 0 1.48932e-08 0 1.48962e-08 0.0021 1.48992e-08 0 1.49542e-08 0 1.49572e-08 0.0021 1.49602e-08 0 1.50152e-08 0 1.50182e-08 0.0021 1.50212e-08 0 1.50762e-08 0 1.50792e-08 0.0021 1.50822e-08 0 1.51372e-08 0 1.51402e-08 0.0021 1.51432e-08 0 1.51982e-08 0 1.52012e-08 0.0021 1.52042e-08 0 1.52592e-08 0 1.52622e-08 0.0021 1.52652e-08 0 1.53202e-08 0 1.53232e-08 0.0021 1.53262e-08 0 1.53812e-08 0 1.53842e-08 0.0021 1.53872e-08 0 1.54422e-08 0 1.54452e-08 0.0021 1.54482e-08 0 1.55032e-08 0 1.55062e-08 0.0021 1.55092e-08 0 1.55642e-08 0 1.55672e-08 0.0021 1.55702e-08 0 1.56252e-08 0 1.56282e-08 0.0021 1.56312e-08 0 1.56862e-08 0 1.56892e-08 0.0021 1.56922e-08 0 1.57472e-08 0 1.57502e-08 0.0021 1.57532e-08 0 1.58082e-08 0 1.58112e-08 0.0021 1.58142e-08 0 1.58692e-08 0 1.58722e-08 0.0021 1.58752e-08 0 1.59302e-08 0 1.59332e-08 0.0021 1.59362e-08 0 1.59912e-08 0 1.59942e-08 0.0021 1.59972e-08 0 1.60522e-08 0 1.60552e-08 0.0021 1.60582e-08 0 1.61132e-08 0 1.61162e-08 0.0021 1.61192e-08 0 1.61742e-08 0 1.61772e-08 0.0021 1.61802e-08 0 1.62352e-08 0 1.62382e-08 0.0021 1.62412e-08 0 1.62962e-08 0 1.62992e-08 0.0021 1.63022e-08 0 1.63572e-08 0 1.63602e-08 0.0021 1.63632e-08 0 1.64182e-08 0 1.64212e-08 0.0021 1.64242e-08 0 1.64792e-08 0 1.64822e-08 0.0021 1.64852e-08 0 1.65402e-08 0 1.65432e-08 0.0021 1.65462e-08 0 1.66012e-08 0 1.66042e-08 0.0021 1.66072e-08 0 1.66622e-08 0 1.66652e-08 0.0021 1.66682e-08 0 1.67232e-08 0 1.67262e-08 0.0021 1.67292e-08 0 1.67842e-08 0 1.67872e-08 0.0021 1.67902e-08 0 1.68452e-08 0 1.68482e-08 0.0021 1.68512e-08 0 1.69062e-08 0 1.69092e-08 0.0021 1.69122e-08 0 1.69672e-08 0 1.69702e-08 0.0021 1.69732e-08 0 1.70282e-08 0 1.70312e-08 0.0021 1.70342e-08 0 1.70892e-08 0 1.70922e-08 0.0021 1.70952e-08 0 1.71502e-08 0 1.71532e-08 0.0021 1.71562e-08 0 1.72112e-08 0 1.72142e-08 0.0021 1.72172e-08 0 1.72722e-08 0 1.72752e-08 0.0021 1.72782e-08 0 1.73332e-08 0 1.73362e-08 0.0021 1.73392e-08 0 1.73942e-08 0 1.73972e-08 0.0021 1.74002e-08 0 1.74552e-08 0 1.74582e-08 0.0021 1.74612e-08 0 1.75162e-08 0 1.75192e-08 0.0021 1.75222e-08 0 1.75772e-08 0 1.75802e-08 0.0021 1.75832e-08 0 1.76382e-08 0 1.76412e-08 0.0021 1.76442e-08 0 1.76992e-08 0 1.77022e-08 0.0021 1.77052e-08 0 1.77602e-08 0 1.77632e-08 0.0021 1.77662e-08 0 1.78212e-08 0 1.78242e-08 0.0021 1.78272e-08 0 1.78822e-08 0 1.78852e-08 0.0021 1.78882e-08 0 1.79432e-08 0 1.79462e-08 0.0021 1.79492e-08 0 1.80042e-08 0 1.80072e-08 0.0021 1.80102e-08 0 1.80652e-08 0 1.80682e-08 0.0021 1.80712e-08 0 1.81262e-08 0 1.81292e-08 0.0021 1.81322e-08 0 1.81872e-08 0 1.81902e-08 0.0021 1.81932e-08 0 1.82482e-08 0 1.82512e-08 0.0021 1.82542e-08 0 1.83092e-08 0 1.83122e-08 0.0021 1.83152e-08 0 1.83702e-08 0 1.83732e-08 0.0021 1.83762e-08 0 1.84312e-08 0 1.84342e-08 0.0021 1.84372e-08 0 1.84922e-08 0 1.84952e-08 0.0021 1.84982e-08 0 1.85532e-08 0 1.85562e-08 0.0021 1.85592e-08 0 1.86142e-08 0 1.86172e-08 0.0021 1.86202e-08 0 1.86752e-08 0 1.86782e-08 0.0021 1.86812e-08 0 1.87362e-08 0 1.87392e-08 0.0021 1.87422e-08 0 1.87972e-08 0 1.88002e-08 0.0021 1.88032e-08 0 1.88582e-08 0 1.88612e-08 0.0021 1.88642e-08 0 1.89192e-08 0 1.89222e-08 0.0021 1.89252e-08 0 1.89802e-08 0 1.89832e-08 0.0021 1.89862e-08 0 1.90412e-08 0 1.90442e-08 0.0021 1.90472e-08 0 1.91022e-08 0 1.91052e-08 0.0021 1.91082e-08 0 1.91632e-08 0 1.91662e-08 0.0021 1.91692e-08 0 1.92242e-08 0 1.92272e-08 0.0021 1.92302e-08 0 1.92852e-08 0 1.92882e-08 0.0021 1.92912e-08 0 1.93462e-08 0 1.93492e-08 0.0021 1.93522e-08 0 1.94072e-08 0 1.94102e-08 0.0021 1.94132e-08 0 1.94682e-08 0 1.94712e-08 0.0021 1.94742e-08 0 1.95292e-08 0 1.95322e-08 0.0021 1.95352e-08 0 1.95902e-08 0 1.95932e-08 0.0021 1.95962e-08 0 1.96512e-08 0 1.96542e-08 0.0021 1.96572e-08 0 1.97122e-08 0 1.97152e-08 0.0021 1.97182e-08 0 1.97732e-08 0 1.97762e-08 0.0021 1.97792e-08 0 1.98342e-08 0 1.98372e-08 0.0021 1.98402e-08 0 1.98952e-08 0 1.98982e-08 0.0021 1.99012e-08 0 1.99562e-08 0 1.99592e-08 0.0021 1.99622e-08 0 2.00172e-08 0 2.00202e-08 0.0021 2.00232e-08 0 2.00782e-08 0 2.00812e-08 0.0021 2.00842e-08 0 2.01392e-08 0 2.01422e-08 0.0021 2.01452e-08 0 2.02002e-08 0 2.02032e-08 0.0021 2.02062e-08 0 2.02612e-08 0 2.02642e-08 0.0021 2.02672e-08 0 2.03222e-08 0 2.03252e-08 0.0021 2.03282e-08 0 2.03832e-08 0 2.03862e-08 0.0021 2.03892e-08 0 2.04442e-08 0 2.04472e-08 0.0021 2.04502e-08 0 2.05052e-08 0 2.05082e-08 0.0021 2.05112e-08 0 2.05662e-08 0 2.05692e-08 0.0021 2.05722e-08 0 2.06272e-08 0 2.06302e-08 0.0021 2.06332e-08 0 2.06882e-08 0 2.06912e-08 0.0021 2.06942e-08 0 2.07492e-08 0 2.07522e-08 0.0021 2.07552e-08 0 2.08102e-08 0 2.08132e-08 0.0021 2.08162e-08 0 2.08712e-08 0 2.08742e-08 0.0021 2.08772e-08 0 2.09322e-08 0 2.09352e-08 0.0021 2.09382e-08 0 2.09932e-08 0 2.09962e-08 0.0021 2.09992e-08 0 2.10542e-08 0 2.10572e-08 0.0021 2.10602e-08 0 2.11152e-08 0 2.11182e-08 0.0021 2.11212e-08 0 2.11762e-08 0 2.11792e-08 0.0021 2.11822e-08 0 2.12372e-08 0 2.12402e-08 0.0021 2.12432e-08 0 2.12982e-08 0 2.13012e-08 0.0021 2.13042e-08 0 2.13592e-08 0 2.13622e-08 0.0021 2.13652e-08 0 2.14202e-08 0 2.14232e-08 0.0021 2.14262e-08 0 2.14812e-08 0 2.14842e-08 0.0021 2.14872e-08 0 2.15422e-08 0 2.15452e-08 0.0021 2.15482e-08 0 2.16032e-08 0 2.16062e-08 0.0021 2.16092e-08 0 2.16642e-08 0 2.16672e-08 0.0021 2.16702e-08 0 2.17252e-08 0 2.17282e-08 0.0021 2.17312e-08 0 2.17862e-08 0 2.17892e-08 0.0021 2.17922e-08 0 2.18472e-08 0 2.18502e-08 0.0021 2.18532e-08 0 2.19082e-08 0 2.19112e-08 0.0021 2.19142e-08 0 2.19692e-08 0 2.19722e-08 0.0021 2.19752e-08 0 2.20302e-08 0 2.20332e-08 0.0021 2.20362e-08 0 2.20912e-08 0 2.20942e-08 0.0021 2.20972e-08 0 2.21522e-08 0 2.21552e-08 0.0021 2.21582e-08 0 2.22132e-08 0 2.22162e-08 0.0021 2.22192e-08 0 2.22742e-08 0 2.22772e-08 0.0021 2.22802e-08 0 2.23352e-08 0 2.23382e-08 0.0021 2.23412e-08 0 2.23962e-08 0 2.23992e-08 0.0021 2.24022e-08 0 2.24572e-08 0 2.24602e-08 0.0021 2.24632e-08 0 2.25182e-08 0 2.25212e-08 0.0021 2.25242e-08 0 2.25792e-08 0 2.25822e-08 0.0021 2.25852e-08 0 2.26402e-08 0 2.26432e-08 0.0021 2.26462e-08 0 2.27012e-08 0 2.27042e-08 0.0021 2.27072e-08 0 2.27622e-08 0 2.27652e-08 0.0021 2.27682e-08 0 2.28232e-08 0 2.28262e-08 0.0021 2.28292e-08 0 2.28842e-08 0 2.28872e-08 0.0021 2.28902e-08 0 2.29452e-08 0 2.29482e-08 0.0021 2.29512e-08 0 2.30062e-08 0 2.30092e-08 0.0021 2.30122e-08 0 2.30672e-08 0 2.30702e-08 0.0021 2.30732e-08 0 2.31282e-08 0 2.31312e-08 0.0021 2.31342e-08 0 2.31892e-08 0 2.31922e-08 0.0021 2.31952e-08 0 2.32502e-08 0 2.32532e-08 0.0021 2.32562e-08 0 2.33112e-08 0 2.33142e-08 0.0021 2.33172e-08 0 2.33722e-08 0 2.33752e-08 0.0021 2.33782e-08 0 2.34332e-08 0 2.34362e-08 0.0021 2.34392e-08 0 2.34942e-08 0 2.34972e-08 0.0021 2.35002e-08 0 2.35552e-08 0 2.35582e-08 0.0021 2.35612e-08 0 2.36162e-08 0 2.36192e-08 0.0021 2.36222e-08 0 2.36772e-08 0 2.36802e-08 0.0021 2.36832e-08 0 2.37382e-08 0 2.37412e-08 0.0021 2.37442e-08 0 2.37992e-08 0 2.38022e-08 0.0021 2.38052e-08 0 2.38602e-08 0 2.38632e-08 0.0021 2.38662e-08 0 2.39212e-08 0 2.39242e-08 0.0021 2.39272e-08 0 2.39822e-08 0 2.39852e-08 0.0021 2.39882e-08 0 2.40432e-08 0 2.40462e-08 0.0021 2.40492e-08 0 2.41042e-08 0 2.41072e-08 0.0021 2.41102e-08 0 2.41652e-08 0 2.41682e-08 0.0021 2.41712e-08 0 2.42262e-08 0 2.42292e-08 0.0021 2.42322e-08 0 2.42872e-08 0 2.42902e-08 0.0021 2.42932e-08 0)
LSPL_IG0_0|1 IG0_0_RX SPL_IG0_0|D1  2e-12
LSPL_IG0_0|2 SPL_IG0_0|D1 SPL_IG0_0|D2  4.135667696e-12
LSPL_IG0_0|3 SPL_IG0_0|D2 SPL_IG0_0|JCT  9.84682784761905e-13
LSPL_IG0_0|4 SPL_IG0_0|JCT SPL_IG0_0|QA1  9.84682784761905e-13
LSPL_IG0_0|5 SPL_IG0_0|QA1 IG0_0_TO0  2e-12
LSPL_IG0_0|6 SPL_IG0_0|JCT SPL_IG0_0|QB1  9.84682784761905e-13
LSPL_IG0_0|7 SPL_IG0_0|QB1 IG0_0_TO1  2e-12
LSPL_IP1_0|1 IP1_0_RX SPL_IP1_0|D1  2e-12
LSPL_IP1_0|2 SPL_IP1_0|D1 SPL_IP1_0|D2  4.135667696e-12
LSPL_IP1_0|3 SPL_IP1_0|D2 SPL_IP1_0|JCT  9.84682784761905e-13
LSPL_IP1_0|4 SPL_IP1_0|JCT SPL_IP1_0|QA1  9.84682784761905e-13
LSPL_IP1_0|5 SPL_IP1_0|QA1 IP1_0_TO1  2e-12
LSPL_IP1_0|6 SPL_IP1_0|JCT SPL_IP1_0|QB1  9.84682784761905e-13
LSPL_IP1_0|7 SPL_IP1_0|QB1 IP1_0_OUT  2e-12
LSPL_IG2_0|1 IG2_0_RX SPL_IG2_0|D1  2e-12
LSPL_IG2_0|2 SPL_IG2_0|D1 SPL_IG2_0|D2  4.135667696e-12
LSPL_IG2_0|3 SPL_IG2_0|D2 SPL_IG2_0|JCT  9.84682784761905e-13
LSPL_IG2_0|4 SPL_IG2_0|JCT SPL_IG2_0|QA1  9.84682784761905e-13
LSPL_IG2_0|5 SPL_IG2_0|QA1 IG2_0_TO2  2e-12
LSPL_IG2_0|6 SPL_IG2_0|JCT SPL_IG2_0|QB1  9.84682784761905e-13
LSPL_IG2_0|7 SPL_IG2_0|QB1 IG2_0_TO3  2e-12
LSPL_IP3_0|1 IP3_0_RX SPL_IP3_0|D1  2e-12
LSPL_IP3_0|2 SPL_IP3_0|D1 SPL_IP3_0|D2  4.135667696e-12
LSPL_IP3_0|3 SPL_IP3_0|D2 SPL_IP3_0|JCT  9.84682784761905e-13
LSPL_IP3_0|4 SPL_IP3_0|JCT SPL_IP3_0|QA1  9.84682784761905e-13
LSPL_IP3_0|5 SPL_IP3_0|QA1 IP3_0_TO1  2e-12
LSPL_IP3_0|6 SPL_IP3_0|JCT SPL_IP3_0|QB1  9.84682784761905e-13
LSPL_IP3_0|7 SPL_IP3_0|QB1 IP3_0_OUT  2e-12
IT04|T 0 T04  PWL(0 0 6.15e-12 0 9.15e-12 0.0014 1.215e-11 0 6.715e-11 0 7.015e-11 0.0014 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0014 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0014 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0014 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0014 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0014 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0014 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0014 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0014 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0014 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0014 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0014 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0014 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0014 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0014 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0014 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0014 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0014 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0014 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0014 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0014 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0014 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0014 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0014 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0014 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0014 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0014 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0014 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0014 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0014 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0014 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0014 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0014 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0014 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0014 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0014 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0014 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0014 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0014 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0014 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0014 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0014 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0014 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0014 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0014 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0014 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0014 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0014 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0014 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0014 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0014 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0014 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0014 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0014 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0014 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0014 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0014 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0014 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0014 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0014 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0014 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0014 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0014 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0014 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0014 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0014 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0014 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0014 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0014 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0014 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0014 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0014 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0014 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0014 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0014 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0014 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0014 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0014 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0014 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0014 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0014 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0014 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0014 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0014 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0014 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0014 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0014 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0014 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0014 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0014 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0014 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0014 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0014 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0014 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0014 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0014 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0014 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0014 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0014 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0014 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0014 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0014 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0014 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0014 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0014 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0014 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0014 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0014 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0014 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0014 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0014 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0014 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0014 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0014 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0014 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0014 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0014 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0014 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0014 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0014 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0014 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0014 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0014 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0014 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0014 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0014 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0014 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0014 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0014 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0014 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0014 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0014 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0014 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0014 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0014 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0014 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0014 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0014 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0014 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0014 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0014 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0014 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0014 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0014 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0014 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0014 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0014 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0014 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0014 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0014 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0014 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0014 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0014 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0014 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0014 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0014 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0014 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0014 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0014 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0014 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0014 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0014 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0014 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0014 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0014 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0014 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0014 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0014 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0014 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0014 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0014 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0014 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0014 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0014 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0014 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0014 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0014 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0014 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0014 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0014 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0014 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0014 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0014 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0014 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0014 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0014 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0014 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0014 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0014 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0014 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0014 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0014 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0014 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0014 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0014 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0014 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0014 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0014 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0014 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0014 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0014 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0014 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0014 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0014 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0014 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0014 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0014 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0014 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0014 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0014 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0014 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0014 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0014 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0014 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0014 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0014 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0014 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0014 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0014 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0014 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0014 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0014 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0014 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0014 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0014 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0014 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0014 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0014 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0014 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0014 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0014 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0014 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0014 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0014 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0014 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0014 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0014 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0014 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0014 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0014 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0014 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0014 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0014 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0014 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0014 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0014 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0014 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0014 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0014 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0014 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0014 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0014 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0014 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0014 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0014 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0014 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0014 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0014 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0014 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0014 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0014 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0014 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0014 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0014 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0014 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0014 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0014 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0014 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0014 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0014 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0014 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0014 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0014 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0014 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0014 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0014 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0014 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0014 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0014 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0014 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0014 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0014 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0014 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0014 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0014 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0014 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0014 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0014 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0014 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0014 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0014 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0014 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0014 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0014 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0014 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0014 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0014 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0014 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0014 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0014 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0014 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0014 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0014 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0014 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0014 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0014 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0014 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0014 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0014 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0014 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0014 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0014 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0014 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0014 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0014 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0014 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0014 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0014 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0014 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0014 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0014 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0014 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0014 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0014 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0014 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0014 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0014 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0014 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0014 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0014 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0014 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0014 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0014 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0014 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0014 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0014 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0014 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0014 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0014 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0014 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0014 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0014 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0014 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0014 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0014 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0014 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0014 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0014 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0014 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0014 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0014 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0014 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0014 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0014 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0014 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0014 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0014 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0014 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0014 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0014 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0014 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0014 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0014 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0014 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0014 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0014 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0014 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0014 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0014 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0014 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0014 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0014 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0014 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0014 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0014 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0014 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0014 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0014 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0014 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0014 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0014 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0014 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0014 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0014 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0014 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0014 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0014 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0014 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0014 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0014 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0014 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0014 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0014 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0014 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0014 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0014 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0014 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0014 2.42901e-08 0)
IT05|T 0 T05  PWL(0 0 6.15e-12 0 9.15e-12 0.0014 1.215e-11 0 6.715e-11 0 7.015e-11 0.0014 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0014 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0014 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0014 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0014 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0014 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0014 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0014 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0014 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0014 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0014 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0014 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0014 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0014 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0014 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0014 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0014 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0014 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0014 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0014 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0014 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0014 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0014 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0014 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0014 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0014 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0014 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0014 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0014 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0014 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0014 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0014 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0014 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0014 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0014 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0014 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0014 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0014 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0014 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0014 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0014 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0014 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0014 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0014 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0014 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0014 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0014 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0014 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0014 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0014 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0014 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0014 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0014 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0014 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0014 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0014 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0014 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0014 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0014 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0014 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0014 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0014 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0014 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0014 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0014 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0014 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0014 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0014 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0014 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0014 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0014 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0014 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0014 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0014 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0014 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0014 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0014 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0014 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0014 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0014 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0014 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0014 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0014 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0014 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0014 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0014 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0014 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0014 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0014 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0014 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0014 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0014 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0014 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0014 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0014 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0014 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0014 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0014 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0014 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0014 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0014 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0014 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0014 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0014 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0014 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0014 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0014 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0014 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0014 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0014 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0014 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0014 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0014 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0014 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0014 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0014 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0014 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0014 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0014 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0014 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0014 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0014 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0014 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0014 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0014 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0014 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0014 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0014 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0014 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0014 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0014 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0014 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0014 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0014 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0014 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0014 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0014 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0014 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0014 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0014 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0014 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0014 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0014 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0014 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0014 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0014 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0014 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0014 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0014 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0014 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0014 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0014 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0014 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0014 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0014 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0014 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0014 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0014 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0014 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0014 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0014 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0014 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0014 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0014 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0014 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0014 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0014 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0014 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0014 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0014 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0014 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0014 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0014 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0014 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0014 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0014 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0014 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0014 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0014 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0014 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0014 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0014 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0014 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0014 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0014 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0014 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0014 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0014 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0014 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0014 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0014 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0014 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0014 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0014 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0014 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0014 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0014 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0014 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0014 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0014 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0014 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0014 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0014 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0014 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0014 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0014 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0014 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0014 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0014 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0014 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0014 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0014 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0014 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0014 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0014 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0014 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0014 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0014 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0014 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0014 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0014 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0014 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0014 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0014 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0014 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0014 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0014 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0014 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0014 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0014 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0014 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0014 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0014 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0014 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0014 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0014 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0014 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0014 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0014 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0014 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0014 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0014 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0014 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0014 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0014 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0014 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0014 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0014 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0014 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0014 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0014 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0014 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0014 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0014 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0014 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0014 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0014 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0014 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0014 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0014 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0014 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0014 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0014 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0014 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0014 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0014 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0014 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0014 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0014 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0014 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0014 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0014 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0014 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0014 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0014 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0014 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0014 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0014 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0014 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0014 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0014 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0014 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0014 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0014 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0014 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0014 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0014 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0014 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0014 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0014 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0014 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0014 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0014 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0014 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0014 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0014 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0014 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0014 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0014 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0014 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0014 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0014 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0014 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0014 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0014 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0014 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0014 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0014 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0014 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0014 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0014 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0014 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0014 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0014 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0014 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0014 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0014 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0014 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0014 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0014 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0014 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0014 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0014 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0014 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0014 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0014 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0014 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0014 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0014 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0014 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0014 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0014 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0014 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0014 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0014 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0014 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0014 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0014 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0014 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0014 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0014 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0014 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0014 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0014 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0014 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0014 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0014 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0014 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0014 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0014 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0014 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0014 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0014 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0014 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0014 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0014 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0014 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0014 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0014 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0014 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0014 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0014 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0014 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0014 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0014 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0014 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0014 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0014 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0014 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0014 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0014 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0014 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0014 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0014 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0014 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0014 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0014 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0014 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0014 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0014 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0014 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0014 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0014 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0014 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0014 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0014 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0014 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0014 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0014 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0014 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0014 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0014 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0014 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0014 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0014 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0014 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0014 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0014 2.42901e-08 0)
IT06|T 0 T06  PWL(0 0 6.15e-12 0 9.15e-12 0.0014 1.215e-11 0 6.715e-11 0 7.015e-11 0.0014 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0014 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0014 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0014 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0014 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0014 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0014 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0014 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0014 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0014 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0014 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0014 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0014 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0014 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0014 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0014 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0014 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0014 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0014 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0014 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0014 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0014 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0014 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0014 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0014 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0014 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0014 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0014 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0014 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0014 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0014 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0014 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0014 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0014 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0014 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0014 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0014 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0014 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0014 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0014 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0014 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0014 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0014 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0014 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0014 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0014 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0014 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0014 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0014 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0014 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0014 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0014 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0014 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0014 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0014 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0014 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0014 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0014 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0014 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0014 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0014 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0014 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0014 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0014 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0014 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0014 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0014 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0014 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0014 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0014 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0014 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0014 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0014 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0014 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0014 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0014 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0014 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0014 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0014 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0014 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0014 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0014 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0014 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0014 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0014 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0014 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0014 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0014 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0014 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0014 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0014 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0014 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0014 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0014 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0014 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0014 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0014 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0014 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0014 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0014 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0014 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0014 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0014 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0014 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0014 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0014 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0014 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0014 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0014 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0014 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0014 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0014 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0014 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0014 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0014 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0014 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0014 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0014 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0014 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0014 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0014 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0014 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0014 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0014 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0014 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0014 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0014 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0014 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0014 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0014 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0014 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0014 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0014 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0014 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0014 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0014 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0014 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0014 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0014 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0014 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0014 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0014 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0014 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0014 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0014 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0014 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0014 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0014 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0014 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0014 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0014 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0014 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0014 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0014 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0014 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0014 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0014 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0014 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0014 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0014 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0014 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0014 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0014 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0014 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0014 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0014 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0014 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0014 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0014 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0014 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0014 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0014 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0014 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0014 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0014 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0014 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0014 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0014 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0014 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0014 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0014 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0014 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0014 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0014 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0014 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0014 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0014 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0014 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0014 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0014 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0014 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0014 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0014 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0014 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0014 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0014 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0014 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0014 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0014 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0014 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0014 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0014 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0014 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0014 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0014 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0014 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0014 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0014 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0014 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0014 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0014 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0014 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0014 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0014 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0014 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0014 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0014 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0014 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0014 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0014 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0014 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0014 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0014 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0014 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0014 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0014 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0014 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0014 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0014 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0014 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0014 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0014 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0014 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0014 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0014 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0014 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0014 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0014 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0014 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0014 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0014 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0014 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0014 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0014 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0014 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0014 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0014 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0014 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0014 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0014 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0014 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0014 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0014 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0014 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0014 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0014 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0014 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0014 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0014 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0014 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0014 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0014 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0014 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0014 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0014 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0014 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0014 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0014 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0014 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0014 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0014 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0014 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0014 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0014 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0014 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0014 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0014 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0014 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0014 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0014 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0014 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0014 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0014 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0014 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0014 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0014 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0014 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0014 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0014 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0014 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0014 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0014 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0014 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0014 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0014 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0014 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0014 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0014 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0014 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0014 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0014 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0014 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0014 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0014 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0014 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0014 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0014 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0014 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0014 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0014 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0014 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0014 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0014 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0014 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0014 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0014 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0014 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0014 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0014 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0014 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0014 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0014 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0014 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0014 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0014 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0014 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0014 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0014 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0014 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0014 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0014 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0014 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0014 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0014 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0014 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0014 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0014 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0014 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0014 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0014 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0014 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0014 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0014 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0014 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0014 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0014 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0014 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0014 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0014 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0014 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0014 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0014 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0014 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0014 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0014 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0014 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0014 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0014 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0014 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0014 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0014 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0014 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0014 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0014 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0014 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0014 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0014 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0014 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0014 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0014 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0014 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0014 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0014 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0014 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0014 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0014 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0014 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0014 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0014 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0014 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0014 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0014 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0014 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0014 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0014 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0014 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0014 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0014 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0014 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0014 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0014 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0014 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0014 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0014 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0014 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0014 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0014 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0014 2.42901e-08 0)
IT07|T 0 T07  PWL(0 0 6.15e-12 0 9.15e-12 0.0028 1.215e-11 0 6.715e-11 0 7.015e-11 0.0028 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0028 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0028 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0028 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0028 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0028 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0028 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0028 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0028 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0028 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0028 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0028 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0028 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0028 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0028 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0028 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0028 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0028 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0028 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0028 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0028 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0028 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0028 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0028 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0028 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0028 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0028 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0028 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0028 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0028 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0028 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0028 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0028 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0028 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0028 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0028 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0028 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0028 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0028 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0028 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0028 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0028 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0028 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0028 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0028 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0028 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0028 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0028 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0028 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0028 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0028 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0028 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0028 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0028 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0028 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0028 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0028 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0028 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0028 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0028 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0028 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0028 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0028 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0028 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0028 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0028 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0028 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0028 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0028 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0028 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0028 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0028 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0028 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0028 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0028 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0028 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0028 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0028 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0028 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0028 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0028 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0028 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0028 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0028 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0028 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0028 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0028 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0028 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0028 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0028 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0028 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0028 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0028 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0028 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0028 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0028 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0028 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0028 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0028 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0028 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0028 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0028 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0028 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0028 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0028 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0028 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0028 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0028 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0028 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0028 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0028 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0028 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0028 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0028 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0028 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0028 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0028 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0028 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0028 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0028 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0028 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0028 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0028 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0028 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0028 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0028 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0028 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0028 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0028 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0028 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0028 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0028 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0028 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0028 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0028 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0028 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0028 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0028 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0028 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0028 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0028 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0028 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0028 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0028 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0028 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0028 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0028 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0028 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0028 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0028 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0028 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0028 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0028 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0028 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0028 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0028 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0028 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0028 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0028 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0028 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0028 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0028 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0028 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0028 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0028 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0028 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0028 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0028 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0028 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0028 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0028 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0028 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0028 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0028 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0028 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0028 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0028 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0028 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0028 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0028 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0028 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0028 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0028 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0028 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0028 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0028 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0028 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0028 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0028 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0028 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0028 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0028 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0028 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0028 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0028 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0028 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0028 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0028 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0028 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0028 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0028 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0028 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0028 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0028 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0028 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0028 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0028 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0028 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0028 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0028 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0028 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0028 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0028 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0028 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0028 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0028 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0028 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0028 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0028 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0028 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0028 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0028 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0028 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0028 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0028 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0028 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0028 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0028 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0028 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0028 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0028 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0028 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0028 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0028 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0028 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0028 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0028 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0028 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0028 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0028 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0028 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0028 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0028 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0028 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0028 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0028 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0028 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0028 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0028 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0028 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0028 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0028 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0028 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0028 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0028 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0028 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0028 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0028 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0028 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0028 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0028 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0028 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0028 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0028 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0028 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0028 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0028 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0028 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0028 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0028 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0028 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0028 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0028 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0028 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0028 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0028 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0028 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0028 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0028 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0028 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0028 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0028 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0028 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0028 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0028 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0028 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0028 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0028 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0028 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0028 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0028 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0028 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0028 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0028 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0028 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0028 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0028 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0028 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0028 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0028 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0028 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0028 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0028 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0028 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0028 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0028 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0028 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0028 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0028 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0028 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0028 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0028 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0028 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0028 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0028 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0028 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0028 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0028 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0028 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0028 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0028 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0028 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0028 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0028 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0028 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0028 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0028 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0028 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0028 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0028 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0028 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0028 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0028 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0028 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0028 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0028 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0028 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0028 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0028 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0028 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0028 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0028 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0028 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0028 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0028 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0028 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0028 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0028 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0028 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0028 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0028 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0028 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0028 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0028 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0028 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0028 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0028 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0028 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0028 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0028 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0028 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0028 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0028 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0028 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0028 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0028 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0028 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0028 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0028 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0028 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0028 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0028 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0028 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0028 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0028 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0028 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0028 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0028 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0028 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0028 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0028 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0028 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0028 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0028 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0028 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0028 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0028 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0028 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0028 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0028 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0028 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0028 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0028 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0028 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0028 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0028 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0028 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0028 2.42901e-08 0)
ID01|T 0 D01  PWL(0 0 6.15e-12 0 9.15e-12 0.0007 1.215e-11 0 6.715e-11 0 7.015e-11 0.0007 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0007 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0007 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0007 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0007 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0007 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0007 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0007 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0007 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0007 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0007 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0007 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0007 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0007 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0007 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0007 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0007 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0007 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0007 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0007 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0007 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0007 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0007 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0007 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0007 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0007 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0007 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0007 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0007 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0007 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0007 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0007 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0007 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0007 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0007 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0007 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0007 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0007 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0007 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0007 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0007 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0007 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0007 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0007 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0007 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0007 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0007 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0007 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0007 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0007 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0007 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0007 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0007 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0007 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0007 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0007 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0007 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0007 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0007 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0007 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0007 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0007 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0007 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0007 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0007 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0007 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0007 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0007 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0007 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0007 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0007 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0007 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0007 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0007 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0007 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0007 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0007 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0007 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0007 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0007 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0007 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0007 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0007 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0007 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0007 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0007 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0007 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0007 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0007 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0007 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0007 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0007 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0007 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0007 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0007 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0007 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0007 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0007 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0007 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0007 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0007 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0007 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0007 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0007 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0007 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0007 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0007 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0007 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0007 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0007 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0007 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0007 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0007 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0007 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0007 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0007 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0007 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0007 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0007 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0007 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0007 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0007 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0007 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0007 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0007 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0007 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0007 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0007 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0007 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0007 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0007 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0007 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0007 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0007 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0007 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0007 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0007 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0007 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0007 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0007 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0007 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0007 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0007 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0007 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0007 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0007 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0007 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0007 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0007 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0007 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0007 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0007 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0007 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0007 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0007 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0007 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0007 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0007 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0007 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0007 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0007 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0007 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0007 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0007 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0007 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0007 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0007 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0007 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0007 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0007 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0007 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0007 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0007 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0007 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0007 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0007 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0007 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0007 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0007 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0007 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0007 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0007 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0007 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0007 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0007 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0007 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0007 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0007 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0007 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0007 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0007 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0007 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0007 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0007 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0007 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0007 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0007 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0007 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0007 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0007 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0007 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0007 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0007 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0007 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0007 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0007 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0007 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0007 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0007 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0007 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0007 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0007 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0007 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0007 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0007 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0007 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0007 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0007 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0007 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0007 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0007 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0007 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0007 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0007 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0007 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0007 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0007 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0007 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0007 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0007 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0007 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0007 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0007 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0007 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0007 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0007 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0007 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0007 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0007 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0007 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0007 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0007 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0007 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0007 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0007 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0007 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0007 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0007 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0007 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0007 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0007 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0007 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0007 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0007 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0007 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0007 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0007 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0007 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0007 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0007 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0007 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0007 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0007 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0007 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0007 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0007 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0007 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0007 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0007 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0007 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0007 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0007 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0007 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0007 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0007 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0007 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0007 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0007 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0007 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0007 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0007 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0007 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0007 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0007 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0007 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0007 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0007 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0007 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0007 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0007 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0007 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0007 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0007 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0007 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0007 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0007 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0007 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0007 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0007 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0007 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0007 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0007 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0007 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0007 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0007 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0007 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0007 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0007 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0007 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0007 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0007 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0007 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0007 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0007 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0007 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0007 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0007 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0007 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0007 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0007 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0007 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0007 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0007 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0007 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0007 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0007 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0007 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0007 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0007 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0007 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0007 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0007 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0007 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0007 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0007 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0007 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0007 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0007 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0007 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0007 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0007 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0007 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0007 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0007 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0007 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0007 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0007 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0007 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0007 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0007 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0007 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0007 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0007 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0007 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0007 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0007 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0007 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0007 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0007 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0007 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0007 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0007 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0007 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0007 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0007 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0007 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0007 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0007 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0007 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0007 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0007 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0007 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0007 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0007 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0007 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0007 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0007 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0007 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0007 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0007 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0007 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0007 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0007 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0007 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0007 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0007 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0007 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0007 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0007 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0007 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0007 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0007 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0007 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0007 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0007 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0007 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0007 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0007 2.42901e-08 0)
L_DFF_IP1_01|1 IP1_0_OUT _DFF_IP1_01|A1  2.067833848e-12
L_DFF_IP1_01|2 _DFF_IP1_01|A1 _DFF_IP1_01|A2  4.135667696e-12
L_DFF_IP1_01|3 _DFF_IP1_01|A3 _DFF_IP1_01|A4  8.271335392e-12
L_DFF_IP1_01|T D01 _DFF_IP1_01|T1  2.067833848e-12
L_DFF_IP1_01|4 _DFF_IP1_01|T1 _DFF_IP1_01|T2  4.135667696e-12
L_DFF_IP1_01|5 _DFF_IP1_01|A4 _DFF_IP1_01|Q1  4.135667696e-12
L_DFF_IP1_01|6 _DFF_IP1_01|Q1 IP1_1_OUT  2.067833848e-12
ID02|T 0 D02  PWL(0 0 6.15e-12 0 9.15e-12 0.0007 1.215e-11 0 6.715e-11 0 7.015e-11 0.0007 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0007 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0007 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0007 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0007 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0007 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0007 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0007 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0007 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0007 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0007 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0007 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0007 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0007 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0007 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0007 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0007 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0007 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0007 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0007 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0007 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0007 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0007 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0007 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0007 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0007 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0007 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0007 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0007 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0007 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0007 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0007 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0007 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0007 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0007 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0007 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0007 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0007 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0007 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0007 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0007 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0007 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0007 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0007 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0007 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0007 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0007 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0007 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0007 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0007 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0007 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0007 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0007 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0007 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0007 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0007 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0007 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0007 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0007 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0007 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0007 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0007 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0007 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0007 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0007 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0007 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0007 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0007 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0007 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0007 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0007 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0007 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0007 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0007 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0007 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0007 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0007 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0007 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0007 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0007 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0007 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0007 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0007 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0007 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0007 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0007 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0007 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0007 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0007 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0007 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0007 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0007 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0007 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0007 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0007 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0007 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0007 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0007 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0007 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0007 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0007 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0007 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0007 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0007 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0007 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0007 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0007 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0007 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0007 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0007 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0007 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0007 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0007 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0007 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0007 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0007 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0007 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0007 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0007 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0007 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0007 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0007 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0007 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0007 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0007 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0007 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0007 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0007 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0007 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0007 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0007 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0007 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0007 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0007 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0007 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0007 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0007 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0007 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0007 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0007 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0007 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0007 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0007 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0007 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0007 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0007 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0007 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0007 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0007 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0007 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0007 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0007 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0007 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0007 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0007 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0007 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0007 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0007 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0007 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0007 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0007 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0007 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0007 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0007 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0007 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0007 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0007 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0007 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0007 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0007 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0007 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0007 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0007 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0007 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0007 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0007 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0007 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0007 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0007 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0007 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0007 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0007 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0007 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0007 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0007 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0007 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0007 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0007 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0007 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0007 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0007 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0007 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0007 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0007 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0007 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0007 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0007 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0007 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0007 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0007 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0007 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0007 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0007 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0007 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0007 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0007 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0007 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0007 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0007 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0007 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0007 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0007 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0007 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0007 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0007 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0007 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0007 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0007 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0007 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0007 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0007 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0007 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0007 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0007 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0007 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0007 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0007 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0007 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0007 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0007 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0007 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0007 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0007 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0007 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0007 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0007 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0007 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0007 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0007 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0007 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0007 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0007 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0007 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0007 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0007 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0007 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0007 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0007 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0007 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0007 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0007 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0007 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0007 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0007 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0007 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0007 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0007 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0007 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0007 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0007 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0007 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0007 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0007 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0007 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0007 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0007 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0007 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0007 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0007 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0007 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0007 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0007 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0007 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0007 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0007 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0007 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0007 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0007 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0007 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0007 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0007 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0007 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0007 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0007 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0007 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0007 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0007 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0007 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0007 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0007 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0007 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0007 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0007 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0007 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0007 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0007 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0007 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0007 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0007 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0007 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0007 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0007 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0007 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0007 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0007 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0007 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0007 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0007 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0007 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0007 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0007 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0007 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0007 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0007 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0007 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0007 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0007 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0007 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0007 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0007 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0007 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0007 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0007 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0007 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0007 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0007 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0007 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0007 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0007 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0007 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0007 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0007 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0007 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0007 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0007 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0007 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0007 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0007 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0007 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0007 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0007 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0007 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0007 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0007 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0007 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0007 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0007 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0007 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0007 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0007 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0007 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0007 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0007 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0007 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0007 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0007 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0007 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0007 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0007 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0007 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0007 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0007 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0007 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0007 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0007 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0007 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0007 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0007 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0007 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0007 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0007 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0007 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0007 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0007 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0007 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0007 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0007 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0007 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0007 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0007 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0007 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0007 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0007 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0007 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0007 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0007 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0007 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0007 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0007 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0007 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0007 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0007 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0007 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0007 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0007 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0007 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0007 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0007 2.42901e-08 0)
L_DFF_IP2_01|1 IP2_0_OUT _DFF_IP2_01|A1  2.067833848e-12
L_DFF_IP2_01|2 _DFF_IP2_01|A1 _DFF_IP2_01|A2  4.135667696e-12
L_DFF_IP2_01|3 _DFF_IP2_01|A3 _DFF_IP2_01|A4  8.271335392e-12
L_DFF_IP2_01|T D02 _DFF_IP2_01|T1  2.067833848e-12
L_DFF_IP2_01|4 _DFF_IP2_01|T1 _DFF_IP2_01|T2  4.135667696e-12
L_DFF_IP2_01|5 _DFF_IP2_01|A4 _DFF_IP2_01|Q1  4.135667696e-12
L_DFF_IP2_01|6 _DFF_IP2_01|Q1 IP2_1_OUT  2.067833848e-12
ID03|T 0 D03  PWL(0 0 6.15e-12 0 9.15e-12 0.0007 1.215e-11 0 6.715e-11 0 7.015e-11 0.0007 7.315e-11 0 1.2815e-10 0 1.3115e-10 0.0007 1.3415e-10 0 1.8915e-10 0 1.9215e-10 0.0007 1.9515e-10 0 2.5015e-10 0 2.5315e-10 0.0007 2.5615e-10 0 3.1115e-10 0 3.1415e-10 0.0007 3.1715e-10 0 3.7215e-10 0 3.7515e-10 0.0007 3.7815e-10 0 4.3315e-10 0 4.3615e-10 0.0007 4.3915e-10 0 4.9415e-10 0 4.9715e-10 0.0007 5.0015e-10 0 5.5515e-10 0 5.5815e-10 0.0007 5.6115e-10 0 6.1615e-10 0 6.1915e-10 0.0007 6.2215e-10 0 6.7715e-10 0 6.8015e-10 0.0007 6.8315e-10 0 7.3815e-10 0 7.4115e-10 0.0007 7.4415e-10 0 7.9915e-10 0 8.0215e-10 0.0007 8.0515e-10 0 8.6015e-10 0 8.6315e-10 0.0007 8.6615e-10 0 9.2115e-10 0 9.2415e-10 0.0007 9.2715e-10 0 9.8215e-10 0 9.8515e-10 0.0007 9.8815e-10 0 1.04315e-09 0 1.04615e-09 0.0007 1.04915e-09 0 1.10415e-09 0 1.10715e-09 0.0007 1.11015e-09 0 1.16515e-09 0 1.16815e-09 0.0007 1.17115e-09 0 1.22615e-09 0 1.22915e-09 0.0007 1.23215e-09 0 1.28715e-09 0 1.29015e-09 0.0007 1.29315e-09 0 1.34815e-09 0 1.35115e-09 0.0007 1.35415e-09 0 1.40915e-09 0 1.41215e-09 0.0007 1.41515e-09 0 1.47015e-09 0 1.47315e-09 0.0007 1.47615e-09 0 1.53115e-09 0 1.53415e-09 0.0007 1.53715e-09 0 1.59215e-09 0 1.59515e-09 0.0007 1.59815e-09 0 1.65315e-09 0 1.65615e-09 0.0007 1.65915e-09 0 1.71415e-09 0 1.71715e-09 0.0007 1.72015e-09 0 1.77515e-09 0 1.77815e-09 0.0007 1.78115e-09 0 1.83615e-09 0 1.83915e-09 0.0007 1.84215e-09 0 1.89715e-09 0 1.90015e-09 0.0007 1.90315e-09 0 1.95815e-09 0 1.96115e-09 0.0007 1.96415e-09 0 2.01915e-09 0 2.02215e-09 0.0007 2.02515e-09 0 2.08015e-09 0 2.08315e-09 0.0007 2.08615e-09 0 2.14115e-09 0 2.14415e-09 0.0007 2.14715e-09 0 2.20215e-09 0 2.20515e-09 0.0007 2.20815e-09 0 2.26315e-09 0 2.26615e-09 0.0007 2.26915e-09 0 2.32415e-09 0 2.32715e-09 0.0007 2.33015e-09 0 2.38515e-09 0 2.38815e-09 0.0007 2.39115e-09 0 2.44615e-09 0 2.44915e-09 0.0007 2.45215e-09 0 2.50715e-09 0 2.51015e-09 0.0007 2.51315e-09 0 2.56815e-09 0 2.57115e-09 0.0007 2.57415e-09 0 2.62915e-09 0 2.63215e-09 0.0007 2.63515e-09 0 2.69015e-09 0 2.69315e-09 0.0007 2.69615e-09 0 2.75115e-09 0 2.75415e-09 0.0007 2.75715e-09 0 2.81215e-09 0 2.81515e-09 0.0007 2.81815e-09 0 2.87315e-09 0 2.87615e-09 0.0007 2.87915e-09 0 2.93415e-09 0 2.93715e-09 0.0007 2.94015e-09 0 2.99515e-09 0 2.99815e-09 0.0007 3.00115e-09 0 3.05615e-09 0 3.05915e-09 0.0007 3.06215e-09 0 3.11715e-09 0 3.12015e-09 0.0007 3.12315e-09 0 3.17815e-09 0 3.18115e-09 0.0007 3.18415e-09 0 3.23915e-09 0 3.24215e-09 0.0007 3.24515e-09 0 3.30015e-09 0 3.30315e-09 0.0007 3.30615e-09 0 3.36115e-09 0 3.36415e-09 0.0007 3.36715e-09 0 3.42215e-09 0 3.42515e-09 0.0007 3.42815e-09 0 3.48315e-09 0 3.48615e-09 0.0007 3.48915e-09 0 3.54415e-09 0 3.54715e-09 0.0007 3.55015e-09 0 3.60515e-09 0 3.60815e-09 0.0007 3.61115e-09 0 3.66615e-09 0 3.66915e-09 0.0007 3.67215e-09 0 3.72715e-09 0 3.73015e-09 0.0007 3.73315e-09 0 3.78815e-09 0 3.79115e-09 0.0007 3.79415e-09 0 3.84915e-09 0 3.85215e-09 0.0007 3.85515e-09 0 3.91015e-09 0 3.91315e-09 0.0007 3.91615e-09 0 3.97115e-09 0 3.97415e-09 0.0007 3.97715e-09 0 4.03215e-09 0 4.03515e-09 0.0007 4.03815e-09 0 4.09315e-09 0 4.09615e-09 0.0007 4.09915e-09 0 4.15415e-09 0 4.15715e-09 0.0007 4.16015e-09 0 4.21515e-09 0 4.21815e-09 0.0007 4.22115e-09 0 4.27615e-09 0 4.27915e-09 0.0007 4.28215e-09 0 4.33715e-09 0 4.34015e-09 0.0007 4.34315e-09 0 4.39815e-09 0 4.40115e-09 0.0007 4.40415e-09 0 4.45915e-09 0 4.46215e-09 0.0007 4.46515e-09 0 4.52015e-09 0 4.52315e-09 0.0007 4.52615e-09 0 4.58115e-09 0 4.58415e-09 0.0007 4.58715e-09 0 4.64215e-09 0 4.64515e-09 0.0007 4.64815e-09 0 4.70315e-09 0 4.70615e-09 0.0007 4.70915e-09 0 4.76415e-09 0 4.76715e-09 0.0007 4.77015e-09 0 4.82515e-09 0 4.82815e-09 0.0007 4.83115e-09 0 4.88615e-09 0 4.88915e-09 0.0007 4.89215e-09 0 4.94715e-09 0 4.95015e-09 0.0007 4.95315e-09 0 5.00815e-09 0 5.01115e-09 0.0007 5.01415e-09 0 5.06915e-09 0 5.07215e-09 0.0007 5.07515e-09 0 5.13015e-09 0 5.13315e-09 0.0007 5.13615e-09 0 5.19115e-09 0 5.19415e-09 0.0007 5.19715e-09 0 5.25215e-09 0 5.25515e-09 0.0007 5.25815e-09 0 5.31315e-09 0 5.31615e-09 0.0007 5.31915e-09 0 5.37415e-09 0 5.37715e-09 0.0007 5.38015e-09 0 5.43515e-09 0 5.43815e-09 0.0007 5.44115e-09 0 5.49615e-09 0 5.49915e-09 0.0007 5.50215e-09 0 5.55715e-09 0 5.56015e-09 0.0007 5.56315e-09 0 5.61815e-09 0 5.62115e-09 0.0007 5.62415e-09 0 5.67915e-09 0 5.68215e-09 0.0007 5.68515e-09 0 5.74015e-09 0 5.74315e-09 0.0007 5.74615e-09 0 5.80115e-09 0 5.80415e-09 0.0007 5.80715e-09 0 5.86215e-09 0 5.86515e-09 0.0007 5.86815e-09 0 5.92315e-09 0 5.92615e-09 0.0007 5.92915e-09 0 5.98415e-09 0 5.98715e-09 0.0007 5.99015e-09 0 6.04515e-09 0 6.04815e-09 0.0007 6.05115e-09 0 6.10615e-09 0 6.10915e-09 0.0007 6.11215e-09 0 6.16715e-09 0 6.17015e-09 0.0007 6.17315e-09 0 6.22815e-09 0 6.23115e-09 0.0007 6.23415e-09 0 6.28915e-09 0 6.29215e-09 0.0007 6.29515e-09 0 6.35015e-09 0 6.35315e-09 0.0007 6.35615e-09 0 6.41115e-09 0 6.41415e-09 0.0007 6.41715e-09 0 6.47215e-09 0 6.47515e-09 0.0007 6.47815e-09 0 6.53315e-09 0 6.53615e-09 0.0007 6.53915e-09 0 6.59415e-09 0 6.59715e-09 0.0007 6.60015e-09 0 6.65515e-09 0 6.65815e-09 0.0007 6.66115e-09 0 6.71615e-09 0 6.71915e-09 0.0007 6.72215e-09 0 6.77715e-09 0 6.78015e-09 0.0007 6.78315e-09 0 6.83815e-09 0 6.84115e-09 0.0007 6.84415e-09 0 6.89915e-09 0 6.90215e-09 0.0007 6.90515e-09 0 6.96015e-09 0 6.96315e-09 0.0007 6.96615e-09 0 7.02115e-09 0 7.02415e-09 0.0007 7.02715e-09 0 7.08215e-09 0 7.08515e-09 0.0007 7.08815e-09 0 7.14315e-09 0 7.14615e-09 0.0007 7.14915e-09 0 7.20415e-09 0 7.20715e-09 0.0007 7.21015e-09 0 7.26515e-09 0 7.26815e-09 0.0007 7.27115e-09 0 7.32615e-09 0 7.32915e-09 0.0007 7.33215e-09 0 7.38715e-09 0 7.39015e-09 0.0007 7.39315e-09 0 7.44815e-09 0 7.45115e-09 0.0007 7.45415e-09 0 7.50915e-09 0 7.51215e-09 0.0007 7.51515e-09 0 7.57015e-09 0 7.57315e-09 0.0007 7.57615e-09 0 7.63115e-09 0 7.63415e-09 0.0007 7.63715e-09 0 7.69215e-09 0 7.69515e-09 0.0007 7.69815e-09 0 7.75315e-09 0 7.75615e-09 0.0007 7.75915e-09 0 7.81415e-09 0 7.81715e-09 0.0007 7.82015e-09 0 7.87515e-09 0 7.87815e-09 0.0007 7.88115e-09 0 7.93615e-09 0 7.93915e-09 0.0007 7.94215e-09 0 7.99715e-09 0 8.00015e-09 0.0007 8.00315e-09 0 8.05815e-09 0 8.06115e-09 0.0007 8.06415e-09 0 8.11915e-09 0 8.12215e-09 0.0007 8.12515e-09 0 8.18015e-09 0 8.18315e-09 0.0007 8.18615e-09 0 8.24115e-09 0 8.24415e-09 0.0007 8.24715e-09 0 8.30215e-09 0 8.30515e-09 0.0007 8.30815e-09 0 8.36315e-09 0 8.36615e-09 0.0007 8.36915e-09 0 8.42415e-09 0 8.42715e-09 0.0007 8.43015e-09 0 8.48515e-09 0 8.48815e-09 0.0007 8.49115e-09 0 8.54615e-09 0 8.54915e-09 0.0007 8.55215e-09 0 8.60715e-09 0 8.61015e-09 0.0007 8.61315e-09 0 8.66815e-09 0 8.67115e-09 0.0007 8.67415e-09 0 8.72915e-09 0 8.73215e-09 0.0007 8.73515e-09 0 8.79015e-09 0 8.79315e-09 0.0007 8.79615e-09 0 8.85115e-09 0 8.85415e-09 0.0007 8.85715e-09 0 8.91215e-09 0 8.91515e-09 0.0007 8.91815e-09 0 8.97315e-09 0 8.97615e-09 0.0007 8.97915e-09 0 9.03415e-09 0 9.03715e-09 0.0007 9.04015e-09 0 9.09515e-09 0 9.09815e-09 0.0007 9.10115e-09 0 9.15615e-09 0 9.15915e-09 0.0007 9.16215e-09 0 9.21715e-09 0 9.22015e-09 0.0007 9.22315e-09 0 9.27815e-09 0 9.28115e-09 0.0007 9.28415e-09 0 9.33915e-09 0 9.34215e-09 0.0007 9.34515e-09 0 9.40015e-09 0 9.40315e-09 0.0007 9.40615e-09 0 9.46115e-09 0 9.46415e-09 0.0007 9.46715e-09 0 9.52215e-09 0 9.52515e-09 0.0007 9.52815e-09 0 9.58315e-09 0 9.58615e-09 0.0007 9.58915e-09 0 9.64415e-09 0 9.64715e-09 0.0007 9.65015e-09 0 9.70515e-09 0 9.70815e-09 0.0007 9.71115e-09 0 9.76615e-09 0 9.76915e-09 0.0007 9.77215e-09 0 9.82715e-09 0 9.83015e-09 0.0007 9.83315e-09 0 9.88815e-09 0 9.89115e-09 0.0007 9.89415e-09 0 9.94915e-09 0 9.95215e-09 0.0007 9.95515e-09 0 1.00101e-08 0 1.00131e-08 0.0007 1.00161e-08 0 1.00711e-08 0 1.00741e-08 0.0007 1.00771e-08 0 1.01321e-08 0 1.01351e-08 0.0007 1.01381e-08 0 1.01932e-08 0 1.01962e-08 0.0007 1.01992e-08 0 1.02542e-08 0 1.02572e-08 0.0007 1.02602e-08 0 1.03151e-08 0 1.03181e-08 0.0007 1.03212e-08 0 1.03761e-08 0 1.03791e-08 0.0007 1.03821e-08 0 1.04371e-08 0 1.04401e-08 0.0007 1.04431e-08 0 1.04981e-08 0 1.05011e-08 0.0007 1.05041e-08 0 1.05592e-08 0 1.05622e-08 0.0007 1.05652e-08 0 1.06201e-08 0 1.06232e-08 0.0007 1.06262e-08 0 1.06811e-08 0 1.06841e-08 0.0007 1.06871e-08 0 1.07421e-08 0 1.07451e-08 0.0007 1.07481e-08 0 1.08031e-08 0 1.08061e-08 0.0007 1.08091e-08 0 1.08642e-08 0 1.08672e-08 0.0007 1.08702e-08 0 1.09252e-08 0 1.09282e-08 0.0007 1.09312e-08 0 1.09861e-08 0 1.09891e-08 0.0007 1.09921e-08 0 1.10471e-08 0 1.10501e-08 0.0007 1.10531e-08 0 1.11081e-08 0 1.11111e-08 0.0007 1.11141e-08 0 1.11691e-08 0 1.11721e-08 0.0007 1.11751e-08 0 1.12302e-08 0 1.12332e-08 0.0007 1.12362e-08 0 1.12911e-08 0 1.12941e-08 0.0007 1.12972e-08 0 1.13521e-08 0 1.13551e-08 0.0007 1.13581e-08 0 1.14131e-08 0 1.14161e-08 0.0007 1.14191e-08 0 1.14741e-08 0 1.14771e-08 0.0007 1.14801e-08 0 1.15352e-08 0 1.15382e-08 0.0007 1.15412e-08 0 1.15961e-08 0 1.15992e-08 0.0007 1.16022e-08 0 1.16571e-08 0 1.16601e-08 0.0007 1.16631e-08 0 1.17181e-08 0 1.17211e-08 0.0007 1.17241e-08 0 1.17791e-08 0 1.17821e-08 0.0007 1.17851e-08 0 1.18402e-08 0 1.18432e-08 0.0007 1.18462e-08 0 1.19011e-08 0 1.19042e-08 0.0007 1.19072e-08 0 1.19621e-08 0 1.19651e-08 0.0007 1.19681e-08 0 1.20231e-08 0 1.20261e-08 0.0007 1.20291e-08 0 1.20841e-08 0 1.20871e-08 0.0007 1.20901e-08 0 1.21452e-08 0 1.21482e-08 0.0007 1.21512e-08 0 1.22062e-08 0 1.22092e-08 0.0007 1.22122e-08 0 1.22671e-08 0 1.22701e-08 0.0007 1.22731e-08 0 1.23281e-08 0 1.23311e-08 0.0007 1.23341e-08 0 1.23891e-08 0 1.23921e-08 0.0007 1.23951e-08 0 1.24501e-08 0 1.24531e-08 0.0007 1.24561e-08 0 1.25112e-08 0 1.25142e-08 0.0007 1.25172e-08 0 1.25721e-08 0 1.25751e-08 0.0007 1.25782e-08 0 1.26331e-08 0 1.26361e-08 0.0007 1.26391e-08 0 1.26941e-08 0 1.26971e-08 0.0007 1.27001e-08 0 1.27551e-08 0 1.27581e-08 0.0007 1.27611e-08 0 1.28162e-08 0 1.28192e-08 0.0007 1.28222e-08 0 1.28771e-08 0 1.28802e-08 0.0007 1.28832e-08 0 1.29381e-08 0 1.29411e-08 0.0007 1.29441e-08 0 1.29991e-08 0 1.30021e-08 0.0007 1.30051e-08 0 1.30601e-08 0 1.30631e-08 0.0007 1.30661e-08 0 1.31211e-08 0 1.31241e-08 0.0007 1.31271e-08 0 1.31822e-08 0 1.31852e-08 0.0007 1.31882e-08 0 1.32431e-08 0 1.32461e-08 0.0007 1.32491e-08 0 1.33041e-08 0 1.33071e-08 0.0007 1.33101e-08 0 1.33651e-08 0 1.33681e-08 0.0007 1.33711e-08 0 1.34261e-08 0 1.34291e-08 0.0007 1.34321e-08 0 1.34872e-08 0 1.34902e-08 0.0007 1.34932e-08 0 1.35481e-08 0 1.35511e-08 0.0007 1.35541e-08 0 1.36091e-08 0 1.36121e-08 0.0007 1.36151e-08 0 1.36701e-08 0 1.36731e-08 0.0007 1.36761e-08 0 1.37311e-08 0 1.37341e-08 0.0007 1.37371e-08 0 1.37922e-08 0 1.37952e-08 0.0007 1.37982e-08 0 1.38531e-08 0 1.38561e-08 0.0007 1.38592e-08 0 1.39141e-08 0 1.39171e-08 0.0007 1.39201e-08 0 1.39751e-08 0 1.39781e-08 0.0007 1.39811e-08 0 1.40361e-08 0 1.40391e-08 0.0007 1.40421e-08 0 1.40972e-08 0 1.41002e-08 0.0007 1.41032e-08 0 1.41581e-08 0 1.41612e-08 0.0007 1.41642e-08 0 1.42191e-08 0 1.42221e-08 0.0007 1.42251e-08 0 1.42801e-08 0 1.42831e-08 0.0007 1.42861e-08 0 1.43411e-08 0 1.43441e-08 0.0007 1.43471e-08 0 1.44021e-08 0 1.44051e-08 0.0007 1.44081e-08 0 1.44632e-08 0 1.44662e-08 0.0007 1.44692e-08 0 1.45241e-08 0 1.45271e-08 0.0007 1.45301e-08 0 1.45851e-08 0 1.45881e-08 0.0007 1.45911e-08 0 1.46461e-08 0 1.46491e-08 0.0007 1.46521e-08 0 1.47071e-08 0 1.47101e-08 0.0007 1.47131e-08 0 1.47682e-08 0 1.47712e-08 0.0007 1.47742e-08 0 1.48291e-08 0 1.48321e-08 0.0007 1.48351e-08 0 1.48901e-08 0 1.48931e-08 0.0007 1.48961e-08 0 1.49511e-08 0 1.49541e-08 0.0007 1.49571e-08 0 1.50121e-08 0 1.50151e-08 0.0007 1.50181e-08 0 1.50731e-08 0 1.50761e-08 0.0007 1.50791e-08 0 1.51341e-08 0 1.51371e-08 0.0007 1.51401e-08 0 1.51951e-08 0 1.51981e-08 0.0007 1.52011e-08 0 1.52561e-08 0 1.52591e-08 0.0007 1.52621e-08 0 1.53171e-08 0 1.53201e-08 0.0007 1.53231e-08 0 1.53781e-08 0 1.53811e-08 0.0007 1.53841e-08 0 1.54391e-08 0 1.54421e-08 0.0007 1.54451e-08 0 1.55001e-08 0 1.55031e-08 0.0007 1.55061e-08 0 1.55611e-08 0 1.55641e-08 0.0007 1.55671e-08 0 1.56221e-08 0 1.56251e-08 0.0007 1.56281e-08 0 1.56831e-08 0 1.56861e-08 0.0007 1.56891e-08 0 1.57441e-08 0 1.57471e-08 0.0007 1.57501e-08 0 1.58051e-08 0 1.58081e-08 0.0007 1.58111e-08 0 1.58661e-08 0 1.58691e-08 0.0007 1.58721e-08 0 1.59271e-08 0 1.59301e-08 0.0007 1.59331e-08 0 1.59881e-08 0 1.59911e-08 0.0007 1.59941e-08 0 1.60491e-08 0 1.60521e-08 0.0007 1.60551e-08 0 1.61101e-08 0 1.61131e-08 0.0007 1.61161e-08 0 1.61711e-08 0 1.61741e-08 0.0007 1.61771e-08 0 1.62321e-08 0 1.62351e-08 0.0007 1.62381e-08 0 1.62931e-08 0 1.62961e-08 0.0007 1.62991e-08 0 1.63541e-08 0 1.63571e-08 0.0007 1.63601e-08 0 1.64151e-08 0 1.64181e-08 0.0007 1.64211e-08 0 1.64761e-08 0 1.64791e-08 0.0007 1.64821e-08 0 1.65371e-08 0 1.65401e-08 0.0007 1.65431e-08 0 1.65981e-08 0 1.66011e-08 0.0007 1.66041e-08 0 1.66591e-08 0 1.66621e-08 0.0007 1.66651e-08 0 1.67201e-08 0 1.67231e-08 0.0007 1.67261e-08 0 1.67811e-08 0 1.67841e-08 0.0007 1.67871e-08 0 1.68421e-08 0 1.68451e-08 0.0007 1.68481e-08 0 1.69031e-08 0 1.69061e-08 0.0007 1.69091e-08 0 1.69641e-08 0 1.69671e-08 0.0007 1.69701e-08 0 1.70251e-08 0 1.70281e-08 0.0007 1.70311e-08 0 1.70861e-08 0 1.70891e-08 0.0007 1.70921e-08 0 1.71471e-08 0 1.71501e-08 0.0007 1.71531e-08 0 1.72081e-08 0 1.72111e-08 0.0007 1.72141e-08 0 1.72691e-08 0 1.72721e-08 0.0007 1.72751e-08 0 1.73301e-08 0 1.73331e-08 0.0007 1.73361e-08 0 1.73911e-08 0 1.73941e-08 0.0007 1.73971e-08 0 1.74521e-08 0 1.74551e-08 0.0007 1.74581e-08 0 1.75131e-08 0 1.75161e-08 0.0007 1.75191e-08 0 1.75741e-08 0 1.75771e-08 0.0007 1.75801e-08 0 1.76351e-08 0 1.76381e-08 0.0007 1.76411e-08 0 1.76961e-08 0 1.76991e-08 0.0007 1.77021e-08 0 1.77571e-08 0 1.77601e-08 0.0007 1.77631e-08 0 1.78181e-08 0 1.78211e-08 0.0007 1.78241e-08 0 1.78791e-08 0 1.78821e-08 0.0007 1.78851e-08 0 1.79401e-08 0 1.79431e-08 0.0007 1.79461e-08 0 1.80011e-08 0 1.80041e-08 0.0007 1.80071e-08 0 1.80621e-08 0 1.80651e-08 0.0007 1.80681e-08 0 1.81231e-08 0 1.81261e-08 0.0007 1.81291e-08 0 1.81841e-08 0 1.81871e-08 0.0007 1.81901e-08 0 1.82451e-08 0 1.82481e-08 0.0007 1.82511e-08 0 1.83061e-08 0 1.83091e-08 0.0007 1.83121e-08 0 1.83671e-08 0 1.83701e-08 0.0007 1.83731e-08 0 1.84281e-08 0 1.84311e-08 0.0007 1.84341e-08 0 1.84891e-08 0 1.84921e-08 0.0007 1.84951e-08 0 1.85501e-08 0 1.85531e-08 0.0007 1.85561e-08 0 1.86111e-08 0 1.86141e-08 0.0007 1.86171e-08 0 1.86721e-08 0 1.86751e-08 0.0007 1.86781e-08 0 1.87331e-08 0 1.87361e-08 0.0007 1.87391e-08 0 1.87941e-08 0 1.87971e-08 0.0007 1.88001e-08 0 1.88551e-08 0 1.88581e-08 0.0007 1.88611e-08 0 1.89161e-08 0 1.89191e-08 0.0007 1.89221e-08 0 1.89771e-08 0 1.89801e-08 0.0007 1.89831e-08 0 1.90381e-08 0 1.90411e-08 0.0007 1.90441e-08 0 1.90991e-08 0 1.91021e-08 0.0007 1.91051e-08 0 1.91601e-08 0 1.91631e-08 0.0007 1.91661e-08 0 1.92211e-08 0 1.92241e-08 0.0007 1.92271e-08 0 1.92821e-08 0 1.92851e-08 0.0007 1.92881e-08 0 1.93431e-08 0 1.93461e-08 0.0007 1.93491e-08 0 1.94041e-08 0 1.94071e-08 0.0007 1.94101e-08 0 1.94651e-08 0 1.94681e-08 0.0007 1.94711e-08 0 1.95261e-08 0 1.95291e-08 0.0007 1.95321e-08 0 1.95871e-08 0 1.95901e-08 0.0007 1.95931e-08 0 1.96481e-08 0 1.96511e-08 0.0007 1.96541e-08 0 1.97091e-08 0 1.97121e-08 0.0007 1.97151e-08 0 1.97701e-08 0 1.97731e-08 0.0007 1.97761e-08 0 1.98311e-08 0 1.98341e-08 0.0007 1.98371e-08 0 1.98921e-08 0 1.98951e-08 0.0007 1.98981e-08 0 1.99531e-08 0 1.99561e-08 0.0007 1.99591e-08 0 2.00141e-08 0 2.00171e-08 0.0007 2.00201e-08 0 2.00751e-08 0 2.00781e-08 0.0007 2.00811e-08 0 2.01361e-08 0 2.01391e-08 0.0007 2.01421e-08 0 2.01971e-08 0 2.02001e-08 0.0007 2.02031e-08 0 2.02581e-08 0 2.02611e-08 0.0007 2.02641e-08 0 2.03191e-08 0 2.03221e-08 0.0007 2.03251e-08 0 2.03801e-08 0 2.03831e-08 0.0007 2.03861e-08 0 2.04411e-08 0 2.04441e-08 0.0007 2.04471e-08 0 2.05021e-08 0 2.05051e-08 0.0007 2.05081e-08 0 2.05631e-08 0 2.05661e-08 0.0007 2.05691e-08 0 2.06241e-08 0 2.06271e-08 0.0007 2.06301e-08 0 2.06851e-08 0 2.06881e-08 0.0007 2.06911e-08 0 2.07461e-08 0 2.07491e-08 0.0007 2.07521e-08 0 2.08071e-08 0 2.08101e-08 0.0007 2.08131e-08 0 2.08681e-08 0 2.08711e-08 0.0007 2.08741e-08 0 2.09291e-08 0 2.09321e-08 0.0007 2.09351e-08 0 2.09901e-08 0 2.09931e-08 0.0007 2.09961e-08 0 2.10511e-08 0 2.10541e-08 0.0007 2.10571e-08 0 2.11121e-08 0 2.11151e-08 0.0007 2.11181e-08 0 2.11731e-08 0 2.11761e-08 0.0007 2.11791e-08 0 2.12341e-08 0 2.12371e-08 0.0007 2.12401e-08 0 2.12951e-08 0 2.12981e-08 0.0007 2.13011e-08 0 2.13561e-08 0 2.13591e-08 0.0007 2.13621e-08 0 2.14171e-08 0 2.14201e-08 0.0007 2.14231e-08 0 2.14781e-08 0 2.14811e-08 0.0007 2.14841e-08 0 2.15391e-08 0 2.15421e-08 0.0007 2.15451e-08 0 2.16001e-08 0 2.16031e-08 0.0007 2.16061e-08 0 2.16611e-08 0 2.16641e-08 0.0007 2.16671e-08 0 2.17221e-08 0 2.17251e-08 0.0007 2.17281e-08 0 2.17831e-08 0 2.17861e-08 0.0007 2.17891e-08 0 2.18441e-08 0 2.18471e-08 0.0007 2.18501e-08 0 2.19051e-08 0 2.19081e-08 0.0007 2.19111e-08 0 2.19661e-08 0 2.19691e-08 0.0007 2.19721e-08 0 2.20271e-08 0 2.20301e-08 0.0007 2.20331e-08 0 2.20881e-08 0 2.20911e-08 0.0007 2.20941e-08 0 2.21491e-08 0 2.21521e-08 0.0007 2.21551e-08 0 2.22101e-08 0 2.22131e-08 0.0007 2.22161e-08 0 2.22711e-08 0 2.22741e-08 0.0007 2.22771e-08 0 2.23321e-08 0 2.23351e-08 0.0007 2.23381e-08 0 2.23931e-08 0 2.23961e-08 0.0007 2.23991e-08 0 2.24541e-08 0 2.24571e-08 0.0007 2.24601e-08 0 2.25151e-08 0 2.25181e-08 0.0007 2.25211e-08 0 2.25761e-08 0 2.25791e-08 0.0007 2.25821e-08 0 2.26371e-08 0 2.26401e-08 0.0007 2.26431e-08 0 2.26981e-08 0 2.27011e-08 0.0007 2.27041e-08 0 2.27591e-08 0 2.27621e-08 0.0007 2.27651e-08 0 2.28201e-08 0 2.28231e-08 0.0007 2.28261e-08 0 2.28811e-08 0 2.28841e-08 0.0007 2.28871e-08 0 2.29421e-08 0 2.29451e-08 0.0007 2.29481e-08 0 2.30031e-08 0 2.30061e-08 0.0007 2.30091e-08 0 2.30641e-08 0 2.30671e-08 0.0007 2.30701e-08 0 2.31251e-08 0 2.31281e-08 0.0007 2.31311e-08 0 2.31861e-08 0 2.31891e-08 0.0007 2.31921e-08 0 2.32471e-08 0 2.32501e-08 0.0007 2.32531e-08 0 2.33081e-08 0 2.33111e-08 0.0007 2.33141e-08 0 2.33691e-08 0 2.33721e-08 0.0007 2.33751e-08 0 2.34301e-08 0 2.34331e-08 0.0007 2.34361e-08 0 2.34911e-08 0 2.34941e-08 0.0007 2.34971e-08 0 2.35521e-08 0 2.35551e-08 0.0007 2.35581e-08 0 2.36131e-08 0 2.36161e-08 0.0007 2.36191e-08 0 2.36741e-08 0 2.36771e-08 0.0007 2.36801e-08 0 2.37351e-08 0 2.37381e-08 0.0007 2.37411e-08 0 2.37961e-08 0 2.37991e-08 0.0007 2.38021e-08 0 2.38571e-08 0 2.38601e-08 0.0007 2.38631e-08 0 2.39181e-08 0 2.39211e-08 0.0007 2.39241e-08 0 2.39791e-08 0 2.39821e-08 0.0007 2.39851e-08 0 2.40401e-08 0 2.40431e-08 0.0007 2.40461e-08 0 2.41011e-08 0 2.41041e-08 0.0007 2.41071e-08 0 2.41621e-08 0 2.41651e-08 0.0007 2.41681e-08 0 2.42231e-08 0 2.42261e-08 0.0007 2.42291e-08 0 2.42841e-08 0 2.42871e-08 0.0007 2.42901e-08 0)
L_DFF_IP3_01|1 IP3_0_OUT _DFF_IP3_01|A1  2.067833848e-12
L_DFF_IP3_01|2 _DFF_IP3_01|A1 _DFF_IP3_01|A2  4.135667696e-12
L_DFF_IP3_01|3 _DFF_IP3_01|A3 _DFF_IP3_01|A4  8.271335392e-12
L_DFF_IP3_01|T D03 _DFF_IP3_01|T1  2.067833848e-12
L_DFF_IP3_01|4 _DFF_IP3_01|T1 _DFF_IP3_01|T2  4.135667696e-12
L_DFF_IP3_01|5 _DFF_IP3_01|A4 _DFF_IP3_01|Q1  4.135667696e-12
L_DFF_IP3_01|6 _DFF_IP3_01|Q1 IP3_1_OUT  2.067833848e-12
IT08|T 0 T08  PWL(0 0 3.1e-12 0 6.1e-12 0.0014 9.1e-12 0 6.41e-11 0 6.71e-11 0.0014 7.01e-11 0 1.251e-10 0 1.281e-10 0.0014 1.311e-10 0 1.861e-10 0 1.891e-10 0.0014 1.921e-10 0 2.471e-10 0 2.501e-10 0.0014 2.531e-10 0 3.081e-10 0 3.111e-10 0.0014 3.141e-10 0 3.691e-10 0 3.721e-10 0.0014 3.751e-10 0 4.301e-10 0 4.331e-10 0.0014 4.361e-10 0 4.911e-10 0 4.941e-10 0.0014 4.971e-10 0 5.521e-10 0 5.551e-10 0.0014 5.581e-10 0 6.131e-10 0 6.161e-10 0.0014 6.191e-10 0 6.741e-10 0 6.771e-10 0.0014 6.801e-10 0 7.351e-10 0 7.381e-10 0.0014 7.411e-10 0 7.961e-10 0 7.991e-10 0.0014 8.021e-10 0 8.571e-10 0 8.601e-10 0.0014 8.631e-10 0 9.181e-10 0 9.211e-10 0.0014 9.241e-10 0 9.791e-10 0 9.821e-10 0.0014 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0014 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0014 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0014 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0014 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0014 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0014 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0014 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0014 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0014 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0014 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0014 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0014 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0014 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0014 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0014 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0014 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0014 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0014 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0014 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0014 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0014 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0014 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0014 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0014 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0014 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0014 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0014 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0014 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0014 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0014 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0014 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0014 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0014 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0014 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0014 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0014 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0014 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0014 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0014 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0014 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0014 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0014 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0014 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0014 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0014 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0014 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0014 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0014 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0014 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0014 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0014 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0014 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0014 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0014 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0014 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0014 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0014 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0014 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0014 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0014 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0014 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0014 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0014 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0014 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0014 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0014 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0014 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0014 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0014 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0014 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0014 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0014 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0014 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0014 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0014 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0014 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0014 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0014 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0014 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0014 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0014 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0014 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0014 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0014 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0014 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0014 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0014 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0014 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0014 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0014 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0014 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0014 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0014 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0014 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0014 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0014 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0014 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0014 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0014 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0014 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0014 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0014 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0014 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0014 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0014 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0014 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0014 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0014 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0014 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0014 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0014 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0014 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0014 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0014 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0014 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0014 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0014 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0014 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0014 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0014 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0014 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0014 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0014 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0014 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0014 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0014 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0014 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0014 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0014 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0014 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0014 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0014 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0014 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0014 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0014 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0014 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0014 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0014 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0014 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0014 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0014 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0014 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0014 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0014 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0014 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0014 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0014 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0014 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0014 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0014 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0014 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0014 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0014 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0014 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0014 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0014 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0014 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0014 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0014 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0014 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0014 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0014 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0014 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0014 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0014 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0014 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0014 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0014 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0014 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0014 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0014 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0014 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0014 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0014 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0014 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0014 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0014 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0014 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0014 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0014 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0014 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0014 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0014 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0014 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0014 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0014 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0014 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0014 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0014 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0014 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0014 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0014 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0014 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0014 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0014 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0014 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0014 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0014 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0014 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0014 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0014 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0014 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0014 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0014 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0014 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0014 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0014 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0014 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0014 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0014 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0014 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0014 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0014 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0014 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0014 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0014 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0014 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0014 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0014 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0014 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0014 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0014 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0014 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0014 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0014 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0014 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0014 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0014 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0014 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0014 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0014 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0014 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0014 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0014 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0014 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0014 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0014 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0014 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0014 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0014 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0014 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0014 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0014 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0014 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0014 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0014 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0014 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0014 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0014 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0014 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0014 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0014 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0014 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0014 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0014 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0014 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0014 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0014 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0014 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0014 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0014 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0014 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0014 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0014 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0014 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0014 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0014 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0014 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0014 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0014 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0014 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0014 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0014 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0014 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0014 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0014 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0014 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0014 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0014 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0014 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0014 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0014 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0014 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0014 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0014 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0014 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0014 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0014 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0014 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0014 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0014 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0014 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0014 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0014 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0014 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0014 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0014 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0014 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0014 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0014 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0014 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0014 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0014 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0014 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0014 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0014 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0014 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0014 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0014 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0014 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0014 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0014 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0014 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0014 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0014 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0014 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0014 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0014 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0014 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0014 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0014 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0014 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0014 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0014 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0014 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0014 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0014 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0014 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0014 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0014 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0014 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0014 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0014 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0014 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0014 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0014 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0014 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0014 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0014 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0014 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0014 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0014 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0014 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0014 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0014 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0014 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0014 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0014 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0014 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0014 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0014 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0014 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0014 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0014 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0014 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0014 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0014 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0014 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0014 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0014 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0014 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0014 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0014 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0014 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0014 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0014 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0014 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0014 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0014 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0014 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0014 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0014 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0014 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0014 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0014 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0014 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0014 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0014 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0014 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0014 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0014 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0014 2.42871e-08 0)
IT09|T 0 T09  PWL(0 0 3.1e-12 0 6.1e-12 0.0007 9.1e-12 0 6.41e-11 0 6.71e-11 0.0007 7.01e-11 0 1.251e-10 0 1.281e-10 0.0007 1.311e-10 0 1.861e-10 0 1.891e-10 0.0007 1.921e-10 0 2.471e-10 0 2.501e-10 0.0007 2.531e-10 0 3.081e-10 0 3.111e-10 0.0007 3.141e-10 0 3.691e-10 0 3.721e-10 0.0007 3.751e-10 0 4.301e-10 0 4.331e-10 0.0007 4.361e-10 0 4.911e-10 0 4.941e-10 0.0007 4.971e-10 0 5.521e-10 0 5.551e-10 0.0007 5.581e-10 0 6.131e-10 0 6.161e-10 0.0007 6.191e-10 0 6.741e-10 0 6.771e-10 0.0007 6.801e-10 0 7.351e-10 0 7.381e-10 0.0007 7.411e-10 0 7.961e-10 0 7.991e-10 0.0007 8.021e-10 0 8.571e-10 0 8.601e-10 0.0007 8.631e-10 0 9.181e-10 0 9.211e-10 0.0007 9.241e-10 0 9.791e-10 0 9.821e-10 0.0007 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0007 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0007 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0007 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0007 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0007 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0007 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0007 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0007 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0007 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0007 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0007 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0007 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0007 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0007 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0007 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0007 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0007 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0007 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0007 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0007 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0007 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0007 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0007 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0007 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0007 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0007 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0007 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0007 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0007 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0007 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0007 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0007 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0007 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0007 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0007 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0007 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0007 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0007 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0007 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0007 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0007 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0007 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0007 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0007 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0007 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0007 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0007 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0007 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0007 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0007 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0007 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0007 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0007 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0007 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0007 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0007 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0007 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0007 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0007 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0007 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0007 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0007 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0007 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0007 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0007 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0007 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0007 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0007 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0007 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0007 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0007 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0007 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0007 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0007 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0007 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0007 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0007 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0007 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0007 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0007 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0007 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0007 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0007 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0007 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0007 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0007 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0007 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0007 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0007 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0007 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0007 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0007 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0007 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0007 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0007 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0007 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0007 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0007 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0007 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0007 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0007 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0007 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0007 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0007 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0007 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0007 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0007 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0007 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0007 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0007 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0007 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0007 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0007 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0007 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0007 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0007 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0007 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0007 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0007 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0007 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0007 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0007 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0007 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0007 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0007 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0007 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0007 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0007 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0007 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0007 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0007 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0007 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0007 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0007 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0007 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0007 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0007 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0007 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0007 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0007 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0007 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0007 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0007 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0007 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0007 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0007 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0007 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0007 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0007 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0007 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0007 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0007 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0007 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0007 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0007 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0007 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0007 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0007 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0007 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0007 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0007 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0007 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0007 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0007 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0007 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0007 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0007 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0007 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0007 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0007 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0007 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0007 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0007 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0007 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0007 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0007 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0007 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0007 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0007 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0007 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0007 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0007 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0007 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0007 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0007 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0007 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0007 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0007 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0007 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0007 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0007 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0007 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0007 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0007 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0007 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0007 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0007 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0007 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0007 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0007 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0007 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0007 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0007 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0007 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0007 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0007 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0007 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0007 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0007 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0007 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0007 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0007 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0007 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0007 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0007 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0007 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0007 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0007 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0007 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0007 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0007 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0007 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0007 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0007 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0007 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0007 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0007 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0007 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0007 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0007 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0007 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0007 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0007 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0007 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0007 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0007 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0007 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0007 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0007 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0007 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0007 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0007 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0007 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0007 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0007 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0007 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0007 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0007 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0007 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0007 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0007 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0007 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0007 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0007 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0007 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0007 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0007 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0007 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0007 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0007 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0007 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0007 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0007 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0007 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0007 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0007 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0007 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0007 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0007 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0007 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0007 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0007 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0007 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0007 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0007 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0007 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0007 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0007 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0007 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0007 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0007 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0007 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0007 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0007 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0007 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0007 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0007 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0007 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0007 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0007 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0007 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0007 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0007 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0007 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0007 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0007 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0007 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0007 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0007 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0007 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0007 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0007 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0007 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0007 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0007 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0007 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0007 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0007 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0007 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0007 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0007 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0007 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0007 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0007 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0007 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0007 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0007 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0007 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0007 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0007 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0007 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0007 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0007 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0007 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0007 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0007 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0007 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0007 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0007 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0007 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0007 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0007 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0007 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0007 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0007 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0007 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0007 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0007 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0007 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0007 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0007 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0007 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0007 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0007 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0007 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0007 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0007 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0007 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0007 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0007 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0007 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0007 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0007 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0007 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0007 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0007 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0007 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0007 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0007 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0007 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0007 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0007 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0007 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0007 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0007 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0007 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0007 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0007 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0007 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0007 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0007 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0007 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0007 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0007 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0007 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0007 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0007 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0007 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0007 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0007 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0007 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0007 2.42871e-08 0)
L_PG1_12|1 G1_1_TO1 _PG1_12|A1  2.067833848e-12
L_PG1_12|2 _PG1_12|A1 _PG1_12|A2  4.135667696e-12
L_PG1_12|3 _PG1_12|A3 _PG1_12|A4  8.271335392e-12
L_PG1_12|T T09 _PG1_12|T1  2.067833848e-12
L_PG1_12|4 _PG1_12|T1 _PG1_12|T2  4.135667696e-12
L_PG1_12|5 _PG1_12|A4 _PG1_12|Q1  4.135667696e-12
L_PG1_12|6 _PG1_12|Q1 G1_2  2.067833848e-12
IT10|T 0 T10  PWL(0 0 3.1e-12 0 6.1e-12 0.0014 9.1e-12 0 6.41e-11 0 6.71e-11 0.0014 7.01e-11 0 1.251e-10 0 1.281e-10 0.0014 1.311e-10 0 1.861e-10 0 1.891e-10 0.0014 1.921e-10 0 2.471e-10 0 2.501e-10 0.0014 2.531e-10 0 3.081e-10 0 3.111e-10 0.0014 3.141e-10 0 3.691e-10 0 3.721e-10 0.0014 3.751e-10 0 4.301e-10 0 4.331e-10 0.0014 4.361e-10 0 4.911e-10 0 4.941e-10 0.0014 4.971e-10 0 5.521e-10 0 5.551e-10 0.0014 5.581e-10 0 6.131e-10 0 6.161e-10 0.0014 6.191e-10 0 6.741e-10 0 6.771e-10 0.0014 6.801e-10 0 7.351e-10 0 7.381e-10 0.0014 7.411e-10 0 7.961e-10 0 7.991e-10 0.0014 8.021e-10 0 8.571e-10 0 8.601e-10 0.0014 8.631e-10 0 9.181e-10 0 9.211e-10 0.0014 9.241e-10 0 9.791e-10 0 9.821e-10 0.0014 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0014 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0014 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0014 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0014 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0014 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0014 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0014 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0014 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0014 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0014 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0014 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0014 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0014 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0014 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0014 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0014 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0014 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0014 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0014 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0014 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0014 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0014 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0014 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0014 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0014 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0014 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0014 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0014 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0014 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0014 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0014 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0014 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0014 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0014 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0014 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0014 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0014 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0014 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0014 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0014 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0014 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0014 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0014 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0014 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0014 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0014 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0014 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0014 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0014 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0014 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0014 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0014 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0014 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0014 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0014 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0014 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0014 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0014 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0014 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0014 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0014 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0014 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0014 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0014 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0014 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0014 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0014 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0014 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0014 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0014 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0014 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0014 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0014 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0014 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0014 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0014 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0014 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0014 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0014 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0014 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0014 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0014 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0014 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0014 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0014 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0014 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0014 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0014 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0014 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0014 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0014 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0014 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0014 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0014 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0014 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0014 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0014 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0014 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0014 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0014 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0014 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0014 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0014 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0014 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0014 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0014 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0014 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0014 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0014 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0014 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0014 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0014 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0014 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0014 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0014 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0014 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0014 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0014 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0014 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0014 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0014 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0014 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0014 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0014 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0014 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0014 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0014 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0014 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0014 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0014 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0014 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0014 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0014 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0014 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0014 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0014 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0014 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0014 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0014 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0014 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0014 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0014 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0014 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0014 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0014 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0014 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0014 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0014 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0014 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0014 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0014 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0014 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0014 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0014 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0014 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0014 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0014 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0014 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0014 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0014 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0014 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0014 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0014 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0014 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0014 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0014 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0014 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0014 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0014 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0014 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0014 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0014 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0014 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0014 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0014 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0014 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0014 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0014 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0014 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0014 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0014 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0014 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0014 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0014 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0014 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0014 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0014 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0014 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0014 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0014 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0014 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0014 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0014 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0014 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0014 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0014 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0014 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0014 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0014 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0014 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0014 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0014 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0014 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0014 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0014 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0014 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0014 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0014 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0014 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0014 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0014 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0014 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0014 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0014 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0014 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0014 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0014 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0014 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0014 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0014 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0014 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0014 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0014 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0014 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0014 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0014 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0014 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0014 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0014 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0014 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0014 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0014 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0014 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0014 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0014 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0014 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0014 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0014 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0014 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0014 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0014 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0014 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0014 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0014 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0014 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0014 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0014 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0014 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0014 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0014 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0014 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0014 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0014 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0014 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0014 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0014 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0014 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0014 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0014 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0014 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0014 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0014 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0014 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0014 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0014 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0014 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0014 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0014 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0014 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0014 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0014 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0014 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0014 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0014 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0014 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0014 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0014 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0014 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0014 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0014 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0014 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0014 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0014 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0014 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0014 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0014 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0014 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0014 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0014 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0014 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0014 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0014 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0014 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0014 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0014 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0014 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0014 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0014 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0014 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0014 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0014 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0014 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0014 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0014 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0014 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0014 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0014 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0014 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0014 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0014 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0014 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0014 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0014 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0014 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0014 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0014 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0014 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0014 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0014 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0014 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0014 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0014 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0014 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0014 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0014 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0014 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0014 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0014 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0014 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0014 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0014 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0014 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0014 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0014 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0014 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0014 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0014 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0014 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0014 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0014 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0014 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0014 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0014 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0014 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0014 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0014 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0014 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0014 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0014 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0014 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0014 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0014 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0014 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0014 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0014 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0014 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0014 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0014 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0014 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0014 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0014 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0014 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0014 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0014 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0014 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0014 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0014 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0014 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0014 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0014 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0014 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0014 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0014 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0014 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0014 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0014 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0014 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0014 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0014 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0014 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0014 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0014 2.42871e-08 0)
IT11|T 0 T11  PWL(0 0 3.1e-12 0 6.1e-12 0.0014 9.1e-12 0 6.41e-11 0 6.71e-11 0.0014 7.01e-11 0 1.251e-10 0 1.281e-10 0.0014 1.311e-10 0 1.861e-10 0 1.891e-10 0.0014 1.921e-10 0 2.471e-10 0 2.501e-10 0.0014 2.531e-10 0 3.081e-10 0 3.111e-10 0.0014 3.141e-10 0 3.691e-10 0 3.721e-10 0.0014 3.751e-10 0 4.301e-10 0 4.331e-10 0.0014 4.361e-10 0 4.911e-10 0 4.941e-10 0.0014 4.971e-10 0 5.521e-10 0 5.551e-10 0.0014 5.581e-10 0 6.131e-10 0 6.161e-10 0.0014 6.191e-10 0 6.741e-10 0 6.771e-10 0.0014 6.801e-10 0 7.351e-10 0 7.381e-10 0.0014 7.411e-10 0 7.961e-10 0 7.991e-10 0.0014 8.021e-10 0 8.571e-10 0 8.601e-10 0.0014 8.631e-10 0 9.181e-10 0 9.211e-10 0.0014 9.241e-10 0 9.791e-10 0 9.821e-10 0.0014 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0014 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0014 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0014 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0014 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0014 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0014 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0014 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0014 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0014 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0014 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0014 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0014 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0014 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0014 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0014 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0014 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0014 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0014 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0014 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0014 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0014 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0014 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0014 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0014 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0014 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0014 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0014 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0014 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0014 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0014 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0014 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0014 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0014 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0014 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0014 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0014 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0014 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0014 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0014 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0014 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0014 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0014 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0014 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0014 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0014 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0014 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0014 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0014 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0014 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0014 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0014 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0014 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0014 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0014 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0014 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0014 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0014 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0014 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0014 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0014 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0014 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0014 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0014 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0014 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0014 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0014 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0014 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0014 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0014 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0014 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0014 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0014 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0014 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0014 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0014 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0014 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0014 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0014 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0014 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0014 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0014 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0014 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0014 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0014 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0014 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0014 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0014 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0014 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0014 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0014 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0014 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0014 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0014 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0014 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0014 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0014 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0014 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0014 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0014 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0014 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0014 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0014 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0014 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0014 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0014 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0014 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0014 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0014 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0014 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0014 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0014 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0014 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0014 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0014 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0014 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0014 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0014 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0014 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0014 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0014 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0014 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0014 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0014 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0014 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0014 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0014 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0014 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0014 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0014 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0014 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0014 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0014 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0014 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0014 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0014 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0014 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0014 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0014 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0014 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0014 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0014 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0014 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0014 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0014 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0014 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0014 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0014 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0014 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0014 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0014 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0014 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0014 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0014 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0014 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0014 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0014 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0014 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0014 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0014 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0014 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0014 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0014 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0014 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0014 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0014 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0014 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0014 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0014 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0014 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0014 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0014 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0014 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0014 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0014 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0014 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0014 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0014 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0014 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0014 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0014 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0014 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0014 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0014 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0014 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0014 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0014 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0014 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0014 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0014 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0014 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0014 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0014 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0014 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0014 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0014 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0014 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0014 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0014 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0014 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0014 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0014 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0014 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0014 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0014 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0014 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0014 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0014 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0014 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0014 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0014 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0014 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0014 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0014 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0014 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0014 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0014 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0014 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0014 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0014 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0014 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0014 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0014 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0014 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0014 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0014 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0014 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0014 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0014 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0014 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0014 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0014 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0014 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0014 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0014 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0014 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0014 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0014 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0014 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0014 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0014 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0014 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0014 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0014 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0014 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0014 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0014 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0014 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0014 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0014 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0014 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0014 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0014 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0014 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0014 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0014 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0014 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0014 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0014 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0014 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0014 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0014 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0014 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0014 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0014 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0014 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0014 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0014 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0014 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0014 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0014 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0014 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0014 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0014 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0014 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0014 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0014 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0014 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0014 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0014 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0014 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0014 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0014 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0014 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0014 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0014 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0014 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0014 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0014 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0014 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0014 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0014 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0014 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0014 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0014 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0014 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0014 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0014 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0014 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0014 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0014 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0014 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0014 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0014 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0014 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0014 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0014 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0014 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0014 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0014 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0014 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0014 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0014 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0014 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0014 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0014 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0014 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0014 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0014 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0014 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0014 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0014 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0014 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0014 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0014 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0014 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0014 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0014 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0014 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0014 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0014 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0014 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0014 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0014 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0014 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0014 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0014 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0014 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0014 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0014 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0014 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0014 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0014 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0014 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0014 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0014 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0014 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0014 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0014 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0014 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0014 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0014 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0014 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0014 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0014 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0014 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0014 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0014 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0014 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0014 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0014 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0014 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0014 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0014 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0014 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0014 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0014 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0014 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0014 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0014 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0014 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0014 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0014 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0014 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0014 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0014 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0014 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0014 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0014 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0014 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0014 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0014 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0014 2.42871e-08 0)
ID11|T 0 D11  PWL(0 0 3.1e-12 0 6.1e-12 0.0007 9.1e-12 0 6.41e-11 0 6.71e-11 0.0007 7.01e-11 0 1.251e-10 0 1.281e-10 0.0007 1.311e-10 0 1.861e-10 0 1.891e-10 0.0007 1.921e-10 0 2.471e-10 0 2.501e-10 0.0007 2.531e-10 0 3.081e-10 0 3.111e-10 0.0007 3.141e-10 0 3.691e-10 0 3.721e-10 0.0007 3.751e-10 0 4.301e-10 0 4.331e-10 0.0007 4.361e-10 0 4.911e-10 0 4.941e-10 0.0007 4.971e-10 0 5.521e-10 0 5.551e-10 0.0007 5.581e-10 0 6.131e-10 0 6.161e-10 0.0007 6.191e-10 0 6.741e-10 0 6.771e-10 0.0007 6.801e-10 0 7.351e-10 0 7.381e-10 0.0007 7.411e-10 0 7.961e-10 0 7.991e-10 0.0007 8.021e-10 0 8.571e-10 0 8.601e-10 0.0007 8.631e-10 0 9.181e-10 0 9.211e-10 0.0007 9.241e-10 0 9.791e-10 0 9.821e-10 0.0007 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0007 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0007 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0007 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0007 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0007 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0007 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0007 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0007 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0007 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0007 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0007 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0007 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0007 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0007 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0007 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0007 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0007 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0007 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0007 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0007 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0007 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0007 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0007 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0007 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0007 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0007 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0007 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0007 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0007 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0007 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0007 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0007 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0007 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0007 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0007 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0007 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0007 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0007 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0007 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0007 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0007 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0007 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0007 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0007 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0007 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0007 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0007 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0007 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0007 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0007 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0007 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0007 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0007 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0007 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0007 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0007 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0007 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0007 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0007 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0007 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0007 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0007 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0007 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0007 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0007 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0007 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0007 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0007 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0007 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0007 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0007 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0007 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0007 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0007 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0007 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0007 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0007 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0007 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0007 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0007 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0007 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0007 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0007 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0007 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0007 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0007 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0007 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0007 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0007 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0007 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0007 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0007 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0007 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0007 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0007 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0007 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0007 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0007 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0007 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0007 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0007 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0007 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0007 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0007 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0007 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0007 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0007 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0007 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0007 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0007 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0007 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0007 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0007 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0007 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0007 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0007 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0007 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0007 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0007 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0007 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0007 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0007 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0007 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0007 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0007 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0007 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0007 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0007 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0007 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0007 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0007 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0007 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0007 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0007 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0007 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0007 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0007 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0007 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0007 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0007 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0007 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0007 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0007 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0007 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0007 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0007 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0007 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0007 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0007 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0007 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0007 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0007 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0007 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0007 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0007 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0007 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0007 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0007 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0007 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0007 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0007 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0007 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0007 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0007 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0007 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0007 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0007 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0007 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0007 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0007 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0007 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0007 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0007 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0007 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0007 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0007 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0007 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0007 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0007 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0007 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0007 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0007 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0007 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0007 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0007 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0007 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0007 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0007 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0007 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0007 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0007 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0007 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0007 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0007 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0007 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0007 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0007 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0007 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0007 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0007 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0007 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0007 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0007 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0007 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0007 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0007 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0007 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0007 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0007 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0007 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0007 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0007 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0007 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0007 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0007 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0007 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0007 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0007 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0007 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0007 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0007 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0007 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0007 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0007 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0007 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0007 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0007 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0007 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0007 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0007 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0007 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0007 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0007 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0007 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0007 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0007 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0007 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0007 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0007 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0007 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0007 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0007 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0007 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0007 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0007 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0007 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0007 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0007 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0007 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0007 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0007 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0007 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0007 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0007 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0007 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0007 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0007 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0007 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0007 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0007 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0007 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0007 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0007 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0007 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0007 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0007 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0007 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0007 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0007 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0007 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0007 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0007 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0007 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0007 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0007 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0007 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0007 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0007 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0007 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0007 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0007 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0007 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0007 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0007 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0007 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0007 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0007 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0007 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0007 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0007 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0007 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0007 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0007 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0007 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0007 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0007 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0007 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0007 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0007 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0007 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0007 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0007 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0007 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0007 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0007 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0007 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0007 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0007 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0007 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0007 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0007 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0007 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0007 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0007 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0007 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0007 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0007 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0007 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0007 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0007 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0007 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0007 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0007 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0007 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0007 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0007 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0007 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0007 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0007 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0007 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0007 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0007 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0007 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0007 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0007 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0007 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0007 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0007 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0007 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0007 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0007 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0007 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0007 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0007 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0007 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0007 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0007 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0007 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0007 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0007 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0007 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0007 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0007 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0007 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0007 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0007 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0007 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0007 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0007 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0007 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0007 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0007 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0007 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0007 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0007 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0007 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0007 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0007 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0007 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0007 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0007 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0007 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0007 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0007 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0007 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0007 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0007 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0007 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0007 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0007 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0007 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0007 2.42871e-08 0)
L_DFF_IP1_12|1 IP1_1_OUT_RX _DFF_IP1_12|A1  2.067833848e-12
L_DFF_IP1_12|2 _DFF_IP1_12|A1 _DFF_IP1_12|A2  4.135667696e-12
L_DFF_IP1_12|3 _DFF_IP1_12|A3 _DFF_IP1_12|A4  8.271335392e-12
L_DFF_IP1_12|T D11 _DFF_IP1_12|T1  2.067833848e-12
L_DFF_IP1_12|4 _DFF_IP1_12|T1 _DFF_IP1_12|T2  4.135667696e-12
L_DFF_IP1_12|5 _DFF_IP1_12|A4 _DFF_IP1_12|Q1  4.135667696e-12
L_DFF_IP1_12|6 _DFF_IP1_12|Q1 IP1_2_OUT  2.067833848e-12
ID12|T 0 D12  PWL(0 0 3.1e-12 0 6.1e-12 0.0007 9.1e-12 0 6.41e-11 0 6.71e-11 0.0007 7.01e-11 0 1.251e-10 0 1.281e-10 0.0007 1.311e-10 0 1.861e-10 0 1.891e-10 0.0007 1.921e-10 0 2.471e-10 0 2.501e-10 0.0007 2.531e-10 0 3.081e-10 0 3.111e-10 0.0007 3.141e-10 0 3.691e-10 0 3.721e-10 0.0007 3.751e-10 0 4.301e-10 0 4.331e-10 0.0007 4.361e-10 0 4.911e-10 0 4.941e-10 0.0007 4.971e-10 0 5.521e-10 0 5.551e-10 0.0007 5.581e-10 0 6.131e-10 0 6.161e-10 0.0007 6.191e-10 0 6.741e-10 0 6.771e-10 0.0007 6.801e-10 0 7.351e-10 0 7.381e-10 0.0007 7.411e-10 0 7.961e-10 0 7.991e-10 0.0007 8.021e-10 0 8.571e-10 0 8.601e-10 0.0007 8.631e-10 0 9.181e-10 0 9.211e-10 0.0007 9.241e-10 0 9.791e-10 0 9.821e-10 0.0007 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0007 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0007 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0007 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0007 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0007 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0007 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0007 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0007 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0007 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0007 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0007 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0007 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0007 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0007 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0007 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0007 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0007 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0007 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0007 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0007 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0007 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0007 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0007 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0007 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0007 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0007 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0007 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0007 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0007 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0007 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0007 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0007 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0007 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0007 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0007 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0007 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0007 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0007 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0007 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0007 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0007 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0007 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0007 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0007 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0007 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0007 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0007 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0007 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0007 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0007 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0007 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0007 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0007 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0007 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0007 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0007 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0007 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0007 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0007 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0007 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0007 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0007 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0007 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0007 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0007 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0007 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0007 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0007 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0007 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0007 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0007 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0007 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0007 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0007 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0007 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0007 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0007 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0007 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0007 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0007 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0007 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0007 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0007 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0007 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0007 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0007 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0007 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0007 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0007 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0007 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0007 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0007 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0007 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0007 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0007 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0007 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0007 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0007 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0007 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0007 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0007 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0007 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0007 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0007 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0007 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0007 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0007 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0007 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0007 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0007 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0007 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0007 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0007 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0007 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0007 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0007 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0007 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0007 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0007 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0007 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0007 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0007 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0007 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0007 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0007 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0007 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0007 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0007 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0007 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0007 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0007 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0007 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0007 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0007 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0007 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0007 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0007 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0007 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0007 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0007 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0007 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0007 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0007 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0007 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0007 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0007 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0007 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0007 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0007 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0007 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0007 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0007 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0007 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0007 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0007 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0007 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0007 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0007 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0007 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0007 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0007 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0007 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0007 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0007 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0007 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0007 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0007 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0007 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0007 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0007 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0007 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0007 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0007 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0007 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0007 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0007 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0007 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0007 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0007 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0007 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0007 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0007 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0007 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0007 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0007 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0007 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0007 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0007 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0007 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0007 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0007 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0007 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0007 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0007 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0007 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0007 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0007 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0007 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0007 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0007 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0007 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0007 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0007 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0007 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0007 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0007 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0007 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0007 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0007 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0007 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0007 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0007 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0007 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0007 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0007 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0007 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0007 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0007 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0007 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0007 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0007 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0007 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0007 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0007 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0007 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0007 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0007 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0007 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0007 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0007 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0007 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0007 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0007 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0007 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0007 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0007 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0007 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0007 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0007 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0007 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0007 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0007 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0007 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0007 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0007 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0007 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0007 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0007 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0007 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0007 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0007 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0007 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0007 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0007 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0007 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0007 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0007 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0007 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0007 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0007 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0007 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0007 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0007 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0007 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0007 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0007 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0007 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0007 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0007 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0007 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0007 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0007 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0007 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0007 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0007 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0007 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0007 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0007 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0007 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0007 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0007 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0007 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0007 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0007 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0007 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0007 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0007 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0007 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0007 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0007 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0007 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0007 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0007 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0007 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0007 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0007 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0007 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0007 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0007 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0007 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0007 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0007 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0007 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0007 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0007 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0007 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0007 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0007 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0007 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0007 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0007 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0007 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0007 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0007 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0007 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0007 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0007 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0007 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0007 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0007 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0007 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0007 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0007 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0007 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0007 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0007 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0007 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0007 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0007 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0007 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0007 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0007 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0007 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0007 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0007 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0007 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0007 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0007 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0007 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0007 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0007 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0007 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0007 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0007 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0007 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0007 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0007 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0007 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0007 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0007 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0007 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0007 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0007 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0007 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0007 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0007 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0007 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0007 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0007 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0007 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0007 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0007 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0007 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0007 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0007 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0007 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0007 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0007 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0007 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0007 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0007 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0007 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0007 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0007 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0007 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0007 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0007 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0007 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0007 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0007 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0007 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0007 2.42871e-08 0)
L_DFF_IP2_12|1 IP2_1_OUT_RX _DFF_IP2_12|A1  2.067833848e-12
L_DFF_IP2_12|2 _DFF_IP2_12|A1 _DFF_IP2_12|A2  4.135667696e-12
L_DFF_IP2_12|3 _DFF_IP2_12|A3 _DFF_IP2_12|A4  8.271335392e-12
L_DFF_IP2_12|T D12 _DFF_IP2_12|T1  2.067833848e-12
L_DFF_IP2_12|4 _DFF_IP2_12|T1 _DFF_IP2_12|T2  4.135667696e-12
L_DFF_IP2_12|5 _DFF_IP2_12|A4 _DFF_IP2_12|Q1  4.135667696e-12
L_DFF_IP2_12|6 _DFF_IP2_12|Q1 IP2_2_OUT  2.067833848e-12
ID13|T 0 D13  PWL(0 0 3.1e-12 0 6.1e-12 0.0007 9.1e-12 0 6.41e-11 0 6.71e-11 0.0007 7.01e-11 0 1.251e-10 0 1.281e-10 0.0007 1.311e-10 0 1.861e-10 0 1.891e-10 0.0007 1.921e-10 0 2.471e-10 0 2.501e-10 0.0007 2.531e-10 0 3.081e-10 0 3.111e-10 0.0007 3.141e-10 0 3.691e-10 0 3.721e-10 0.0007 3.751e-10 0 4.301e-10 0 4.331e-10 0.0007 4.361e-10 0 4.911e-10 0 4.941e-10 0.0007 4.971e-10 0 5.521e-10 0 5.551e-10 0.0007 5.581e-10 0 6.131e-10 0 6.161e-10 0.0007 6.191e-10 0 6.741e-10 0 6.771e-10 0.0007 6.801e-10 0 7.351e-10 0 7.381e-10 0.0007 7.411e-10 0 7.961e-10 0 7.991e-10 0.0007 8.021e-10 0 8.571e-10 0 8.601e-10 0.0007 8.631e-10 0 9.181e-10 0 9.211e-10 0.0007 9.241e-10 0 9.791e-10 0 9.821e-10 0.0007 9.851e-10 0 1.0401e-09 0 1.0431e-09 0.0007 1.0461e-09 0 1.1011e-09 0 1.1041e-09 0.0007 1.1071e-09 0 1.1621e-09 0 1.1651e-09 0.0007 1.1681e-09 0 1.2231e-09 0 1.2261e-09 0.0007 1.2291e-09 0 1.2841e-09 0 1.2871e-09 0.0007 1.2901e-09 0 1.3451e-09 0 1.3481e-09 0.0007 1.3511e-09 0 1.4061e-09 0 1.4091e-09 0.0007 1.4121e-09 0 1.4671e-09 0 1.4701e-09 0.0007 1.4731e-09 0 1.5281e-09 0 1.5311e-09 0.0007 1.5341e-09 0 1.5891e-09 0 1.5921e-09 0.0007 1.5951e-09 0 1.6501e-09 0 1.6531e-09 0.0007 1.6561e-09 0 1.7111e-09 0 1.7141e-09 0.0007 1.7171e-09 0 1.7721e-09 0 1.7751e-09 0.0007 1.7781e-09 0 1.8331e-09 0 1.8361e-09 0.0007 1.8391e-09 0 1.8941e-09 0 1.8971e-09 0.0007 1.9001e-09 0 1.9551e-09 0 1.9581e-09 0.0007 1.9611e-09 0 2.0161e-09 0 2.0191e-09 0.0007 2.0221e-09 0 2.0771e-09 0 2.0801e-09 0.0007 2.0831e-09 0 2.1381e-09 0 2.1411e-09 0.0007 2.1441e-09 0 2.1991e-09 0 2.2021e-09 0.0007 2.2051e-09 0 2.2601e-09 0 2.2631e-09 0.0007 2.2661e-09 0 2.3211e-09 0 2.3241e-09 0.0007 2.3271e-09 0 2.3821e-09 0 2.3851e-09 0.0007 2.3881e-09 0 2.4431e-09 0 2.4461e-09 0.0007 2.4491e-09 0 2.5041e-09 0 2.5071e-09 0.0007 2.5101e-09 0 2.5651e-09 0 2.5681e-09 0.0007 2.5711e-09 0 2.6261e-09 0 2.6291e-09 0.0007 2.6321e-09 0 2.6871e-09 0 2.6901e-09 0.0007 2.6931e-09 0 2.7481e-09 0 2.7511e-09 0.0007 2.7541e-09 0 2.8091e-09 0 2.8121e-09 0.0007 2.8151e-09 0 2.8701e-09 0 2.8731e-09 0.0007 2.8761e-09 0 2.9311e-09 0 2.9341e-09 0.0007 2.9371e-09 0 2.9921e-09 0 2.9951e-09 0.0007 2.9981e-09 0 3.0531e-09 0 3.0561e-09 0.0007 3.0591e-09 0 3.1141e-09 0 3.1171e-09 0.0007 3.1201e-09 0 3.1751e-09 0 3.1781e-09 0.0007 3.1811e-09 0 3.2361e-09 0 3.2391e-09 0.0007 3.2421e-09 0 3.2971e-09 0 3.3001e-09 0.0007 3.3031e-09 0 3.3581e-09 0 3.3611e-09 0.0007 3.3641e-09 0 3.4191e-09 0 3.4221e-09 0.0007 3.4251e-09 0 3.4801e-09 0 3.4831e-09 0.0007 3.4861e-09 0 3.5411e-09 0 3.5441e-09 0.0007 3.5471e-09 0 3.6021e-09 0 3.6051e-09 0.0007 3.6081e-09 0 3.6631e-09 0 3.6661e-09 0.0007 3.6691e-09 0 3.7241e-09 0 3.7271e-09 0.0007 3.7301e-09 0 3.7851e-09 0 3.7881e-09 0.0007 3.7911e-09 0 3.8461e-09 0 3.8491e-09 0.0007 3.8521e-09 0 3.9071e-09 0 3.9101e-09 0.0007 3.9131e-09 0 3.9681e-09 0 3.9711e-09 0.0007 3.9741e-09 0 4.0291e-09 0 4.0321e-09 0.0007 4.0351e-09 0 4.0901e-09 0 4.0931e-09 0.0007 4.0961e-09 0 4.1511e-09 0 4.1541e-09 0.0007 4.1571e-09 0 4.2121e-09 0 4.2151e-09 0.0007 4.2181e-09 0 4.2731e-09 0 4.2761e-09 0.0007 4.2791e-09 0 4.3341e-09 0 4.3371e-09 0.0007 4.3401e-09 0 4.3951e-09 0 4.3981e-09 0.0007 4.4011e-09 0 4.4561e-09 0 4.4591e-09 0.0007 4.4621e-09 0 4.5171e-09 0 4.5201e-09 0.0007 4.5231e-09 0 4.5781e-09 0 4.5811e-09 0.0007 4.5841e-09 0 4.6391e-09 0 4.6421e-09 0.0007 4.6451e-09 0 4.7001e-09 0 4.7031e-09 0.0007 4.7061e-09 0 4.7611e-09 0 4.7641e-09 0.0007 4.7671e-09 0 4.8221e-09 0 4.8251e-09 0.0007 4.8281e-09 0 4.8831e-09 0 4.8861e-09 0.0007 4.8891e-09 0 4.9441e-09 0 4.9471e-09 0.0007 4.9501e-09 0 5.0051e-09 0 5.0081e-09 0.0007 5.0111e-09 0 5.0661e-09 0 5.0691e-09 0.0007 5.0721e-09 0 5.1271e-09 0 5.1301e-09 0.0007 5.1331e-09 0 5.1881e-09 0 5.1911e-09 0.0007 5.1941e-09 0 5.2491e-09 0 5.2521e-09 0.0007 5.2551e-09 0 5.3101e-09 0 5.3131e-09 0.0007 5.3161e-09 0 5.3711e-09 0 5.3741e-09 0.0007 5.3771e-09 0 5.4321e-09 0 5.4351e-09 0.0007 5.4381e-09 0 5.4931e-09 0 5.4961e-09 0.0007 5.4991e-09 0 5.5541e-09 0 5.5571e-09 0.0007 5.5601e-09 0 5.6151e-09 0 5.6181e-09 0.0007 5.6211e-09 0 5.6761e-09 0 5.6791e-09 0.0007 5.6821e-09 0 5.7371e-09 0 5.7401e-09 0.0007 5.7431e-09 0 5.7981e-09 0 5.8011e-09 0.0007 5.8041e-09 0 5.8591e-09 0 5.8621e-09 0.0007 5.8651e-09 0 5.9201e-09 0 5.9231e-09 0.0007 5.9261e-09 0 5.9811e-09 0 5.9841e-09 0.0007 5.9871e-09 0 6.0421e-09 0 6.0451e-09 0.0007 6.0481e-09 0 6.1031e-09 0 6.1061e-09 0.0007 6.1091e-09 0 6.1641e-09 0 6.1671e-09 0.0007 6.1701e-09 0 6.2251e-09 0 6.2281e-09 0.0007 6.2311e-09 0 6.2861e-09 0 6.2891e-09 0.0007 6.2921e-09 0 6.3471e-09 0 6.3501e-09 0.0007 6.3531e-09 0 6.4081e-09 0 6.4111e-09 0.0007 6.4141e-09 0 6.4691e-09 0 6.4721e-09 0.0007 6.4751e-09 0 6.5301e-09 0 6.5331e-09 0.0007 6.5361e-09 0 6.5911e-09 0 6.5941e-09 0.0007 6.5971e-09 0 6.6521e-09 0 6.6551e-09 0.0007 6.6581e-09 0 6.7131e-09 0 6.7161e-09 0.0007 6.7191e-09 0 6.7741e-09 0 6.7771e-09 0.0007 6.7801e-09 0 6.8351e-09 0 6.8381e-09 0.0007 6.8411e-09 0 6.8961e-09 0 6.8991e-09 0.0007 6.9021e-09 0 6.9571e-09 0 6.9601e-09 0.0007 6.9631e-09 0 7.0181e-09 0 7.0211e-09 0.0007 7.0241e-09 0 7.0791e-09 0 7.0821e-09 0.0007 7.0851e-09 0 7.1401e-09 0 7.1431e-09 0.0007 7.1461e-09 0 7.2011e-09 0 7.2041e-09 0.0007 7.2071e-09 0 7.2621e-09 0 7.2651e-09 0.0007 7.2681e-09 0 7.3231e-09 0 7.3261e-09 0.0007 7.3291e-09 0 7.3841e-09 0 7.3871e-09 0.0007 7.3901e-09 0 7.4451e-09 0 7.4481e-09 0.0007 7.4511e-09 0 7.5061e-09 0 7.5091e-09 0.0007 7.5121e-09 0 7.5671e-09 0 7.5701e-09 0.0007 7.5731e-09 0 7.6281e-09 0 7.6311e-09 0.0007 7.6341e-09 0 7.6891e-09 0 7.6921e-09 0.0007 7.6951e-09 0 7.7501e-09 0 7.7531e-09 0.0007 7.7561e-09 0 7.8111e-09 0 7.8141e-09 0.0007 7.8171e-09 0 7.8721e-09 0 7.8751e-09 0.0007 7.8781e-09 0 7.9331e-09 0 7.9361e-09 0.0007 7.9391e-09 0 7.9941e-09 0 7.9971e-09 0.0007 8.0001e-09 0 8.0551e-09 0 8.0581e-09 0.0007 8.0611e-09 0 8.1161e-09 0 8.1191e-09 0.0007 8.1221e-09 0 8.1771e-09 0 8.1801e-09 0.0007 8.1831e-09 0 8.2381e-09 0 8.2411e-09 0.0007 8.2441e-09 0 8.2991e-09 0 8.3021e-09 0.0007 8.3051e-09 0 8.3601e-09 0 8.3631e-09 0.0007 8.3661e-09 0 8.4211e-09 0 8.4241e-09 0.0007 8.4271e-09 0 8.4821e-09 0 8.4851e-09 0.0007 8.4881e-09 0 8.5431e-09 0 8.5461e-09 0.0007 8.5491e-09 0 8.6041e-09 0 8.6071e-09 0.0007 8.6101e-09 0 8.6651e-09 0 8.6681e-09 0.0007 8.6711e-09 0 8.7261e-09 0 8.7291e-09 0.0007 8.7321e-09 0 8.7871e-09 0 8.7901e-09 0.0007 8.7931e-09 0 8.8481e-09 0 8.8511e-09 0.0007 8.8541e-09 0 8.9091e-09 0 8.9121e-09 0.0007 8.9151e-09 0 8.9701e-09 0 8.9731e-09 0.0007 8.9761e-09 0 9.0311e-09 0 9.0341e-09 0.0007 9.0371e-09 0 9.0921e-09 0 9.0951e-09 0.0007 9.0981e-09 0 9.1531e-09 0 9.1561e-09 0.0007 9.1591e-09 0 9.2141e-09 0 9.2171e-09 0.0007 9.2201e-09 0 9.2751e-09 0 9.2781e-09 0.0007 9.2811e-09 0 9.3361e-09 0 9.3391e-09 0.0007 9.3421e-09 0 9.3971e-09 0 9.4001e-09 0.0007 9.4031e-09 0 9.4581e-09 0 9.4611e-09 0.0007 9.4641e-09 0 9.5191e-09 0 9.5221e-09 0.0007 9.5251e-09 0 9.5801e-09 0 9.5831e-09 0.0007 9.5861e-09 0 9.6411e-09 0 9.6441e-09 0.0007 9.6471e-09 0 9.7021e-09 0 9.7051e-09 0.0007 9.7081e-09 0 9.7631e-09 0 9.7661e-09 0.0007 9.7691e-09 0 9.8241e-09 0 9.8271e-09 0.0007 9.8301e-09 0 9.8851e-09 0 9.8881e-09 0.0007 9.8911e-09 0 9.9461e-09 0 9.9491e-09 0.0007 9.9521e-09 0 1.00071e-08 0 1.00101e-08 0.0007 1.00131e-08 0 1.00681e-08 0 1.00711e-08 0.0007 1.00741e-08 0 1.01291e-08 0 1.01321e-08 0.0007 1.01351e-08 0 1.01901e-08 0 1.01931e-08 0.0007 1.01961e-08 0 1.02511e-08 0 1.02541e-08 0.0007 1.02571e-08 0 1.03121e-08 0 1.03151e-08 0.0007 1.03181e-08 0 1.03731e-08 0 1.03761e-08 0.0007 1.03791e-08 0 1.04341e-08 0 1.04371e-08 0.0007 1.04401e-08 0 1.04951e-08 0 1.04981e-08 0.0007 1.05011e-08 0 1.05561e-08 0 1.05591e-08 0.0007 1.05621e-08 0 1.06171e-08 0 1.06201e-08 0.0007 1.06231e-08 0 1.06781e-08 0 1.06811e-08 0.0007 1.06841e-08 0 1.07391e-08 0 1.07421e-08 0.0007 1.07451e-08 0 1.08001e-08 0 1.08031e-08 0.0007 1.08061e-08 0 1.08611e-08 0 1.08641e-08 0.0007 1.08671e-08 0 1.09221e-08 0 1.09251e-08 0.0007 1.09281e-08 0 1.09831e-08 0 1.09861e-08 0.0007 1.09891e-08 0 1.10441e-08 0 1.10471e-08 0.0007 1.10501e-08 0 1.11051e-08 0 1.11081e-08 0.0007 1.11111e-08 0 1.11661e-08 0 1.11691e-08 0.0007 1.11721e-08 0 1.12271e-08 0 1.12301e-08 0.0007 1.12331e-08 0 1.12881e-08 0 1.12911e-08 0.0007 1.12941e-08 0 1.13491e-08 0 1.13521e-08 0.0007 1.13551e-08 0 1.14101e-08 0 1.14131e-08 0.0007 1.14161e-08 0 1.14711e-08 0 1.14741e-08 0.0007 1.14771e-08 0 1.15321e-08 0 1.15351e-08 0.0007 1.15381e-08 0 1.15931e-08 0 1.15961e-08 0.0007 1.15991e-08 0 1.16541e-08 0 1.16571e-08 0.0007 1.16601e-08 0 1.17151e-08 0 1.17181e-08 0.0007 1.17211e-08 0 1.17761e-08 0 1.17791e-08 0.0007 1.17821e-08 0 1.18371e-08 0 1.18401e-08 0.0007 1.18431e-08 0 1.18981e-08 0 1.19011e-08 0.0007 1.19041e-08 0 1.19591e-08 0 1.19621e-08 0.0007 1.19651e-08 0 1.20201e-08 0 1.20231e-08 0.0007 1.20261e-08 0 1.20811e-08 0 1.20841e-08 0.0007 1.20871e-08 0 1.21421e-08 0 1.21451e-08 0.0007 1.21481e-08 0 1.22031e-08 0 1.22061e-08 0.0007 1.22091e-08 0 1.22641e-08 0 1.22671e-08 0.0007 1.22701e-08 0 1.23251e-08 0 1.23281e-08 0.0007 1.23311e-08 0 1.23861e-08 0 1.23891e-08 0.0007 1.23921e-08 0 1.24471e-08 0 1.24501e-08 0.0007 1.24531e-08 0 1.25081e-08 0 1.25111e-08 0.0007 1.25141e-08 0 1.25691e-08 0 1.25721e-08 0.0007 1.25751e-08 0 1.26301e-08 0 1.26331e-08 0.0007 1.26361e-08 0 1.26911e-08 0 1.26941e-08 0.0007 1.26971e-08 0 1.27521e-08 0 1.27551e-08 0.0007 1.27581e-08 0 1.28131e-08 0 1.28161e-08 0.0007 1.28191e-08 0 1.28741e-08 0 1.28771e-08 0.0007 1.28801e-08 0 1.29351e-08 0 1.29381e-08 0.0007 1.29411e-08 0 1.29961e-08 0 1.29991e-08 0.0007 1.30021e-08 0 1.30571e-08 0 1.30601e-08 0.0007 1.30631e-08 0 1.31181e-08 0 1.31211e-08 0.0007 1.31241e-08 0 1.31791e-08 0 1.31821e-08 0.0007 1.31851e-08 0 1.32401e-08 0 1.32431e-08 0.0007 1.32461e-08 0 1.33011e-08 0 1.33041e-08 0.0007 1.33071e-08 0 1.33621e-08 0 1.33651e-08 0.0007 1.33681e-08 0 1.34231e-08 0 1.34261e-08 0.0007 1.34291e-08 0 1.34841e-08 0 1.34871e-08 0.0007 1.34901e-08 0 1.35451e-08 0 1.35481e-08 0.0007 1.35511e-08 0 1.36061e-08 0 1.36091e-08 0.0007 1.36121e-08 0 1.36671e-08 0 1.36701e-08 0.0007 1.36731e-08 0 1.37281e-08 0 1.37311e-08 0.0007 1.37341e-08 0 1.37891e-08 0 1.37921e-08 0.0007 1.37951e-08 0 1.38501e-08 0 1.38531e-08 0.0007 1.38561e-08 0 1.39111e-08 0 1.39141e-08 0.0007 1.39171e-08 0 1.39721e-08 0 1.39751e-08 0.0007 1.39781e-08 0 1.40331e-08 0 1.40361e-08 0.0007 1.40391e-08 0 1.40941e-08 0 1.40971e-08 0.0007 1.41001e-08 0 1.41551e-08 0 1.41581e-08 0.0007 1.41611e-08 0 1.42161e-08 0 1.42191e-08 0.0007 1.42221e-08 0 1.42771e-08 0 1.42801e-08 0.0007 1.42831e-08 0 1.43381e-08 0 1.43411e-08 0.0007 1.43441e-08 0 1.43991e-08 0 1.44021e-08 0.0007 1.44051e-08 0 1.44601e-08 0 1.44631e-08 0.0007 1.44661e-08 0 1.45211e-08 0 1.45241e-08 0.0007 1.45271e-08 0 1.45821e-08 0 1.45851e-08 0.0007 1.45881e-08 0 1.46431e-08 0 1.46461e-08 0.0007 1.46491e-08 0 1.47041e-08 0 1.47071e-08 0.0007 1.47101e-08 0 1.47651e-08 0 1.47681e-08 0.0007 1.47711e-08 0 1.48261e-08 0 1.48291e-08 0.0007 1.48321e-08 0 1.48871e-08 0 1.48901e-08 0.0007 1.48931e-08 0 1.49481e-08 0 1.49511e-08 0.0007 1.49541e-08 0 1.50091e-08 0 1.50121e-08 0.0007 1.50151e-08 0 1.50701e-08 0 1.50731e-08 0.0007 1.50761e-08 0 1.51311e-08 0 1.51341e-08 0.0007 1.51371e-08 0 1.51921e-08 0 1.51951e-08 0.0007 1.51981e-08 0 1.52531e-08 0 1.52561e-08 0.0007 1.52591e-08 0 1.53141e-08 0 1.53171e-08 0.0007 1.53201e-08 0 1.53751e-08 0 1.53781e-08 0.0007 1.53811e-08 0 1.54361e-08 0 1.54391e-08 0.0007 1.54421e-08 0 1.54971e-08 0 1.55001e-08 0.0007 1.55031e-08 0 1.55581e-08 0 1.55611e-08 0.0007 1.55641e-08 0 1.56191e-08 0 1.56221e-08 0.0007 1.56251e-08 0 1.56801e-08 0 1.56831e-08 0.0007 1.56861e-08 0 1.57411e-08 0 1.57441e-08 0.0007 1.57471e-08 0 1.58021e-08 0 1.58051e-08 0.0007 1.58081e-08 0 1.58631e-08 0 1.58661e-08 0.0007 1.58691e-08 0 1.59241e-08 0 1.59271e-08 0.0007 1.59301e-08 0 1.59851e-08 0 1.59881e-08 0.0007 1.59911e-08 0 1.60461e-08 0 1.60491e-08 0.0007 1.60521e-08 0 1.61071e-08 0 1.61101e-08 0.0007 1.61131e-08 0 1.61681e-08 0 1.61711e-08 0.0007 1.61741e-08 0 1.62291e-08 0 1.62321e-08 0.0007 1.62351e-08 0 1.62901e-08 0 1.62931e-08 0.0007 1.62961e-08 0 1.63511e-08 0 1.63541e-08 0.0007 1.63571e-08 0 1.64121e-08 0 1.64151e-08 0.0007 1.64181e-08 0 1.64731e-08 0 1.64761e-08 0.0007 1.64791e-08 0 1.65341e-08 0 1.65371e-08 0.0007 1.65401e-08 0 1.65951e-08 0 1.65981e-08 0.0007 1.66011e-08 0 1.66561e-08 0 1.66591e-08 0.0007 1.66621e-08 0 1.67171e-08 0 1.67201e-08 0.0007 1.67231e-08 0 1.67781e-08 0 1.67811e-08 0.0007 1.67841e-08 0 1.68391e-08 0 1.68421e-08 0.0007 1.68451e-08 0 1.69001e-08 0 1.69031e-08 0.0007 1.69061e-08 0 1.69611e-08 0 1.69641e-08 0.0007 1.69671e-08 0 1.70221e-08 0 1.70251e-08 0.0007 1.70281e-08 0 1.70831e-08 0 1.70861e-08 0.0007 1.70891e-08 0 1.71441e-08 0 1.71471e-08 0.0007 1.71501e-08 0 1.72051e-08 0 1.72081e-08 0.0007 1.72111e-08 0 1.72661e-08 0 1.72691e-08 0.0007 1.72721e-08 0 1.73271e-08 0 1.73301e-08 0.0007 1.73331e-08 0 1.73881e-08 0 1.73911e-08 0.0007 1.73941e-08 0 1.74491e-08 0 1.74521e-08 0.0007 1.74551e-08 0 1.75101e-08 0 1.75131e-08 0.0007 1.75161e-08 0 1.75711e-08 0 1.75741e-08 0.0007 1.75771e-08 0 1.76321e-08 0 1.76351e-08 0.0007 1.76381e-08 0 1.76931e-08 0 1.76961e-08 0.0007 1.76991e-08 0 1.77541e-08 0 1.77571e-08 0.0007 1.77601e-08 0 1.78151e-08 0 1.78181e-08 0.0007 1.78211e-08 0 1.78761e-08 0 1.78791e-08 0.0007 1.78821e-08 0 1.79371e-08 0 1.79401e-08 0.0007 1.79431e-08 0 1.79981e-08 0 1.80011e-08 0.0007 1.80041e-08 0 1.80591e-08 0 1.80621e-08 0.0007 1.80651e-08 0 1.81201e-08 0 1.81231e-08 0.0007 1.81261e-08 0 1.81811e-08 0 1.81841e-08 0.0007 1.81871e-08 0 1.82421e-08 0 1.82451e-08 0.0007 1.82481e-08 0 1.83031e-08 0 1.83061e-08 0.0007 1.83091e-08 0 1.83641e-08 0 1.83671e-08 0.0007 1.83701e-08 0 1.84251e-08 0 1.84281e-08 0.0007 1.84311e-08 0 1.84861e-08 0 1.84891e-08 0.0007 1.84921e-08 0 1.85471e-08 0 1.85501e-08 0.0007 1.85531e-08 0 1.86081e-08 0 1.86111e-08 0.0007 1.86141e-08 0 1.86691e-08 0 1.86721e-08 0.0007 1.86751e-08 0 1.87301e-08 0 1.87331e-08 0.0007 1.87361e-08 0 1.87911e-08 0 1.87941e-08 0.0007 1.87971e-08 0 1.88521e-08 0 1.88551e-08 0.0007 1.88581e-08 0 1.89131e-08 0 1.89161e-08 0.0007 1.89191e-08 0 1.89741e-08 0 1.89771e-08 0.0007 1.89801e-08 0 1.90351e-08 0 1.90381e-08 0.0007 1.90411e-08 0 1.90961e-08 0 1.90991e-08 0.0007 1.91021e-08 0 1.91571e-08 0 1.91601e-08 0.0007 1.91631e-08 0 1.92181e-08 0 1.92211e-08 0.0007 1.92241e-08 0 1.92791e-08 0 1.92821e-08 0.0007 1.92851e-08 0 1.93401e-08 0 1.93431e-08 0.0007 1.93461e-08 0 1.94011e-08 0 1.94041e-08 0.0007 1.94071e-08 0 1.94621e-08 0 1.94651e-08 0.0007 1.94681e-08 0 1.95231e-08 0 1.95261e-08 0.0007 1.95291e-08 0 1.95841e-08 0 1.95871e-08 0.0007 1.95901e-08 0 1.96451e-08 0 1.96481e-08 0.0007 1.96511e-08 0 1.97061e-08 0 1.97091e-08 0.0007 1.97121e-08 0 1.97671e-08 0 1.97701e-08 0.0007 1.97731e-08 0 1.98281e-08 0 1.98311e-08 0.0007 1.98341e-08 0 1.98891e-08 0 1.98921e-08 0.0007 1.98951e-08 0 1.99501e-08 0 1.99531e-08 0.0007 1.99561e-08 0 2.00111e-08 0 2.00141e-08 0.0007 2.00171e-08 0 2.00721e-08 0 2.00751e-08 0.0007 2.00781e-08 0 2.01331e-08 0 2.01361e-08 0.0007 2.01391e-08 0 2.01941e-08 0 2.01971e-08 0.0007 2.02001e-08 0 2.02551e-08 0 2.02581e-08 0.0007 2.02611e-08 0 2.03161e-08 0 2.03191e-08 0.0007 2.03221e-08 0 2.03771e-08 0 2.03801e-08 0.0007 2.03831e-08 0 2.04381e-08 0 2.04411e-08 0.0007 2.04441e-08 0 2.04991e-08 0 2.05021e-08 0.0007 2.05051e-08 0 2.05601e-08 0 2.05631e-08 0.0007 2.05661e-08 0 2.06211e-08 0 2.06241e-08 0.0007 2.06271e-08 0 2.06821e-08 0 2.06851e-08 0.0007 2.06881e-08 0 2.07431e-08 0 2.07461e-08 0.0007 2.07491e-08 0 2.08041e-08 0 2.08071e-08 0.0007 2.08101e-08 0 2.08651e-08 0 2.08681e-08 0.0007 2.08711e-08 0 2.09261e-08 0 2.09291e-08 0.0007 2.09321e-08 0 2.09871e-08 0 2.09901e-08 0.0007 2.09931e-08 0 2.10481e-08 0 2.10511e-08 0.0007 2.10541e-08 0 2.11091e-08 0 2.11121e-08 0.0007 2.11151e-08 0 2.11701e-08 0 2.11731e-08 0.0007 2.11761e-08 0 2.12311e-08 0 2.12341e-08 0.0007 2.12371e-08 0 2.12921e-08 0 2.12951e-08 0.0007 2.12981e-08 0 2.13531e-08 0 2.13561e-08 0.0007 2.13591e-08 0 2.14141e-08 0 2.14171e-08 0.0007 2.14201e-08 0 2.14751e-08 0 2.14781e-08 0.0007 2.14811e-08 0 2.15361e-08 0 2.15391e-08 0.0007 2.15421e-08 0 2.15971e-08 0 2.16001e-08 0.0007 2.16031e-08 0 2.16581e-08 0 2.16611e-08 0.0007 2.16641e-08 0 2.17191e-08 0 2.17221e-08 0.0007 2.17251e-08 0 2.17801e-08 0 2.17831e-08 0.0007 2.17861e-08 0 2.18411e-08 0 2.18441e-08 0.0007 2.18471e-08 0 2.19021e-08 0 2.19051e-08 0.0007 2.19081e-08 0 2.19631e-08 0 2.19661e-08 0.0007 2.19691e-08 0 2.20241e-08 0 2.20271e-08 0.0007 2.20301e-08 0 2.20851e-08 0 2.20881e-08 0.0007 2.20911e-08 0 2.21461e-08 0 2.21491e-08 0.0007 2.21521e-08 0 2.22071e-08 0 2.22101e-08 0.0007 2.22131e-08 0 2.22681e-08 0 2.22711e-08 0.0007 2.22741e-08 0 2.23291e-08 0 2.23321e-08 0.0007 2.23351e-08 0 2.23901e-08 0 2.23931e-08 0.0007 2.23961e-08 0 2.24511e-08 0 2.24541e-08 0.0007 2.24571e-08 0 2.25121e-08 0 2.25151e-08 0.0007 2.25181e-08 0 2.25731e-08 0 2.25761e-08 0.0007 2.25791e-08 0 2.26341e-08 0 2.26371e-08 0.0007 2.26401e-08 0 2.26951e-08 0 2.26981e-08 0.0007 2.27011e-08 0 2.27561e-08 0 2.27591e-08 0.0007 2.27621e-08 0 2.28171e-08 0 2.28201e-08 0.0007 2.28231e-08 0 2.28781e-08 0 2.28811e-08 0.0007 2.28841e-08 0 2.29391e-08 0 2.29421e-08 0.0007 2.29451e-08 0 2.30001e-08 0 2.30031e-08 0.0007 2.30061e-08 0 2.30611e-08 0 2.30641e-08 0.0007 2.30671e-08 0 2.31221e-08 0 2.31251e-08 0.0007 2.31281e-08 0 2.31831e-08 0 2.31861e-08 0.0007 2.31891e-08 0 2.32441e-08 0 2.32471e-08 0.0007 2.32501e-08 0 2.33051e-08 0 2.33081e-08 0.0007 2.33111e-08 0 2.33661e-08 0 2.33691e-08 0.0007 2.33721e-08 0 2.34271e-08 0 2.34301e-08 0.0007 2.34331e-08 0 2.34881e-08 0 2.34911e-08 0.0007 2.34941e-08 0 2.35491e-08 0 2.35521e-08 0.0007 2.35551e-08 0 2.36101e-08 0 2.36131e-08 0.0007 2.36161e-08 0 2.36711e-08 0 2.36741e-08 0.0007 2.36771e-08 0 2.37321e-08 0 2.37351e-08 0.0007 2.37381e-08 0 2.37931e-08 0 2.37961e-08 0.0007 2.37991e-08 0 2.38541e-08 0 2.38571e-08 0.0007 2.38601e-08 0 2.39151e-08 0 2.39181e-08 0.0007 2.39211e-08 0 2.39761e-08 0 2.39791e-08 0.0007 2.39821e-08 0 2.40371e-08 0 2.40401e-08 0.0007 2.40431e-08 0 2.40981e-08 0 2.41011e-08 0.0007 2.41041e-08 0 2.41591e-08 0 2.41621e-08 0.0007 2.41651e-08 0 2.42201e-08 0 2.42231e-08 0.0007 2.42261e-08 0 2.42811e-08 0 2.42841e-08 0.0007 2.42871e-08 0)
L_DFF_IP3_12|1 IP3_1_OUT_RX _DFF_IP3_12|A1  2.067833848e-12
L_DFF_IP3_12|2 _DFF_IP3_12|A1 _DFF_IP3_12|A2  4.135667696e-12
L_DFF_IP3_12|3 _DFF_IP3_12|A3 _DFF_IP3_12|A4  8.271335392e-12
L_DFF_IP3_12|T D13 _DFF_IP3_12|T1  2.067833848e-12
L_DFF_IP3_12|4 _DFF_IP3_12|T1 _DFF_IP3_12|T2  4.135667696e-12
L_DFF_IP3_12|5 _DFF_IP3_12|A4 _DFF_IP3_12|Q1  4.135667696e-12
L_DFF_IP3_12|6 _DFF_IP3_12|Q1 IP3_2_OUT  2.067833848e-12
IT12|T 0 T12  PWL(0 0 5e-14 0 3.05e-12 0.0007 6.05e-12 0 6.105e-11 0 6.405e-11 0.0007 6.705e-11 0 1.2205e-10 0 1.2505e-10 0.0007 1.2805e-10 0 1.8305e-10 0 1.8605e-10 0.0007 1.8905e-10 0 2.4405e-10 0 2.4705e-10 0.0007 2.5005e-10 0 3.0505e-10 0 3.0805e-10 0.0007 3.1105e-10 0 3.6605e-10 0 3.6905e-10 0.0007 3.7205e-10 0 4.2705e-10 0 4.3005e-10 0.0007 4.3305e-10 0 4.8805e-10 0 4.9105e-10 0.0007 4.9405e-10 0 5.4905e-10 0 5.5205e-10 0.0007 5.5505e-10 0 6.1005e-10 0 6.1305e-10 0.0007 6.1605e-10 0 6.7105e-10 0 6.7405e-10 0.0007 6.7705e-10 0 7.3205e-10 0 7.3505e-10 0.0007 7.3805e-10 0 7.9305e-10 0 7.9605e-10 0.0007 7.9905e-10 0 8.5405e-10 0 8.5705e-10 0.0007 8.6005e-10 0 9.1505e-10 0 9.1805e-10 0.0007 9.2105e-10 0 9.7605e-10 0 9.7905e-10 0.0007 9.8205e-10 0 1.03705e-09 0 1.04005e-09 0.0007 1.04305e-09 0 1.09805e-09 0 1.10105e-09 0.0007 1.10405e-09 0 1.15905e-09 0 1.16205e-09 0.0007 1.16505e-09 0 1.22005e-09 0 1.22305e-09 0.0007 1.22605e-09 0 1.28105e-09 0 1.28405e-09 0.0007 1.28705e-09 0 1.34205e-09 0 1.34505e-09 0.0007 1.34805e-09 0 1.40305e-09 0 1.40605e-09 0.0007 1.40905e-09 0 1.46405e-09 0 1.46705e-09 0.0007 1.47005e-09 0 1.52505e-09 0 1.52805e-09 0.0007 1.53105e-09 0 1.58605e-09 0 1.58905e-09 0.0007 1.59205e-09 0 1.64705e-09 0 1.65005e-09 0.0007 1.65305e-09 0 1.70805e-09 0 1.71105e-09 0.0007 1.71405e-09 0 1.76905e-09 0 1.77205e-09 0.0007 1.77505e-09 0 1.83005e-09 0 1.83305e-09 0.0007 1.83605e-09 0 1.89105e-09 0 1.89405e-09 0.0007 1.89705e-09 0 1.95205e-09 0 1.95505e-09 0.0007 1.95805e-09 0 2.01305e-09 0 2.01605e-09 0.0007 2.01905e-09 0 2.07405e-09 0 2.07705e-09 0.0007 2.08005e-09 0 2.13505e-09 0 2.13805e-09 0.0007 2.14105e-09 0 2.19605e-09 0 2.19905e-09 0.0007 2.20205e-09 0 2.25705e-09 0 2.26005e-09 0.0007 2.26305e-09 0 2.31805e-09 0 2.32105e-09 0.0007 2.32405e-09 0 2.37905e-09 0 2.38205e-09 0.0007 2.38505e-09 0 2.44005e-09 0 2.44305e-09 0.0007 2.44605e-09 0 2.50105e-09 0 2.50405e-09 0.0007 2.50705e-09 0 2.56205e-09 0 2.56505e-09 0.0007 2.56805e-09 0 2.62305e-09 0 2.62605e-09 0.0007 2.62905e-09 0 2.68405e-09 0 2.68705e-09 0.0007 2.69005e-09 0 2.74505e-09 0 2.74805e-09 0.0007 2.75105e-09 0 2.80605e-09 0 2.80905e-09 0.0007 2.81205e-09 0 2.86705e-09 0 2.87005e-09 0.0007 2.87305e-09 0 2.92805e-09 0 2.93105e-09 0.0007 2.93405e-09 0 2.98905e-09 0 2.99205e-09 0.0007 2.99505e-09 0 3.05005e-09 0 3.05305e-09 0.0007 3.05605e-09 0 3.11105e-09 0 3.11405e-09 0.0007 3.11705e-09 0 3.17205e-09 0 3.17505e-09 0.0007 3.17805e-09 0 3.23305e-09 0 3.23605e-09 0.0007 3.23905e-09 0 3.29405e-09 0 3.29705e-09 0.0007 3.30005e-09 0 3.35505e-09 0 3.35805e-09 0.0007 3.36105e-09 0 3.41605e-09 0 3.41905e-09 0.0007 3.42205e-09 0 3.47705e-09 0 3.48005e-09 0.0007 3.48305e-09 0 3.53805e-09 0 3.54105e-09 0.0007 3.54405e-09 0 3.59905e-09 0 3.60205e-09 0.0007 3.60505e-09 0 3.66005e-09 0 3.66305e-09 0.0007 3.66605e-09 0 3.72105e-09 0 3.72405e-09 0.0007 3.72705e-09 0 3.78205e-09 0 3.78505e-09 0.0007 3.78805e-09 0 3.84305e-09 0 3.84605e-09 0.0007 3.84905e-09 0 3.90405e-09 0 3.90705e-09 0.0007 3.91005e-09 0 3.96505e-09 0 3.96805e-09 0.0007 3.97105e-09 0 4.02605e-09 0 4.02905e-09 0.0007 4.03205e-09 0 4.08705e-09 0 4.09005e-09 0.0007 4.09305e-09 0 4.14805e-09 0 4.15105e-09 0.0007 4.15405e-09 0 4.20905e-09 0 4.21205e-09 0.0007 4.21505e-09 0 4.27005e-09 0 4.27305e-09 0.0007 4.27605e-09 0 4.33105e-09 0 4.33405e-09 0.0007 4.33705e-09 0 4.39205e-09 0 4.39505e-09 0.0007 4.39805e-09 0 4.45305e-09 0 4.45605e-09 0.0007 4.45905e-09 0 4.51405e-09 0 4.51705e-09 0.0007 4.52005e-09 0 4.57505e-09 0 4.57805e-09 0.0007 4.58105e-09 0 4.63605e-09 0 4.63905e-09 0.0007 4.64205e-09 0 4.69705e-09 0 4.70005e-09 0.0007 4.70305e-09 0 4.75805e-09 0 4.76105e-09 0.0007 4.76405e-09 0 4.81905e-09 0 4.82205e-09 0.0007 4.82505e-09 0 4.88005e-09 0 4.88305e-09 0.0007 4.88605e-09 0 4.94105e-09 0 4.94405e-09 0.0007 4.94705e-09 0 5.00205e-09 0 5.00505e-09 0.0007 5.00805e-09 0 5.06305e-09 0 5.06605e-09 0.0007 5.06905e-09 0 5.12405e-09 0 5.12705e-09 0.0007 5.13005e-09 0 5.18505e-09 0 5.18805e-09 0.0007 5.19105e-09 0 5.24605e-09 0 5.24905e-09 0.0007 5.25205e-09 0 5.30705e-09 0 5.31005e-09 0.0007 5.31305e-09 0 5.36805e-09 0 5.37105e-09 0.0007 5.37405e-09 0 5.42905e-09 0 5.43205e-09 0.0007 5.43505e-09 0 5.49005e-09 0 5.49305e-09 0.0007 5.49605e-09 0 5.55105e-09 0 5.55405e-09 0.0007 5.55705e-09 0 5.61205e-09 0 5.61505e-09 0.0007 5.61805e-09 0 5.67305e-09 0 5.67605e-09 0.0007 5.67905e-09 0 5.73405e-09 0 5.73705e-09 0.0007 5.74005e-09 0 5.79505e-09 0 5.79805e-09 0.0007 5.80105e-09 0 5.85605e-09 0 5.85905e-09 0.0007 5.86205e-09 0 5.91705e-09 0 5.92005e-09 0.0007 5.92305e-09 0 5.97805e-09 0 5.98105e-09 0.0007 5.98405e-09 0 6.03905e-09 0 6.04205e-09 0.0007 6.04505e-09 0 6.10005e-09 0 6.10305e-09 0.0007 6.10605e-09 0 6.16105e-09 0 6.16405e-09 0.0007 6.16705e-09 0 6.22205e-09 0 6.22505e-09 0.0007 6.22805e-09 0 6.28305e-09 0 6.28605e-09 0.0007 6.28905e-09 0 6.34405e-09 0 6.34705e-09 0.0007 6.35005e-09 0 6.40505e-09 0 6.40805e-09 0.0007 6.41105e-09 0 6.46605e-09 0 6.46905e-09 0.0007 6.47205e-09 0 6.52705e-09 0 6.53005e-09 0.0007 6.53305e-09 0 6.58805e-09 0 6.59105e-09 0.0007 6.59405e-09 0 6.64905e-09 0 6.65205e-09 0.0007 6.65505e-09 0 6.71005e-09 0 6.71305e-09 0.0007 6.71605e-09 0 6.77105e-09 0 6.77405e-09 0.0007 6.77705e-09 0 6.83205e-09 0 6.83505e-09 0.0007 6.83805e-09 0 6.89305e-09 0 6.89605e-09 0.0007 6.89905e-09 0 6.95405e-09 0 6.95705e-09 0.0007 6.96005e-09 0 7.01505e-09 0 7.01805e-09 0.0007 7.02105e-09 0 7.07605e-09 0 7.07905e-09 0.0007 7.08205e-09 0 7.13705e-09 0 7.14005e-09 0.0007 7.14305e-09 0 7.19805e-09 0 7.20105e-09 0.0007 7.20405e-09 0 7.25905e-09 0 7.26205e-09 0.0007 7.26505e-09 0 7.32005e-09 0 7.32305e-09 0.0007 7.32605e-09 0 7.38105e-09 0 7.38405e-09 0.0007 7.38705e-09 0 7.44205e-09 0 7.44505e-09 0.0007 7.44805e-09 0 7.50305e-09 0 7.50605e-09 0.0007 7.50905e-09 0 7.56405e-09 0 7.56705e-09 0.0007 7.57005e-09 0 7.62505e-09 0 7.62805e-09 0.0007 7.63105e-09 0 7.68605e-09 0 7.68905e-09 0.0007 7.69205e-09 0 7.74705e-09 0 7.75005e-09 0.0007 7.75305e-09 0 7.80805e-09 0 7.81105e-09 0.0007 7.81405e-09 0 7.86905e-09 0 7.87205e-09 0.0007 7.87505e-09 0 7.93005e-09 0 7.93305e-09 0.0007 7.93605e-09 0 7.99105e-09 0 7.99405e-09 0.0007 7.99705e-09 0 8.05205e-09 0 8.05505e-09 0.0007 8.05805e-09 0 8.11305e-09 0 8.11605e-09 0.0007 8.11905e-09 0 8.17405e-09 0 8.17705e-09 0.0007 8.18005e-09 0 8.23505e-09 0 8.23805e-09 0.0007 8.24105e-09 0 8.29605e-09 0 8.29905e-09 0.0007 8.30205e-09 0 8.35705e-09 0 8.36005e-09 0.0007 8.36305e-09 0 8.41805e-09 0 8.42105e-09 0.0007 8.42405e-09 0 8.47905e-09 0 8.48205e-09 0.0007 8.48505e-09 0 8.54005e-09 0 8.54305e-09 0.0007 8.54605e-09 0 8.60105e-09 0 8.60405e-09 0.0007 8.60705e-09 0 8.66205e-09 0 8.66505e-09 0.0007 8.66805e-09 0 8.72305e-09 0 8.72605e-09 0.0007 8.72905e-09 0 8.78405e-09 0 8.78705e-09 0.0007 8.79005e-09 0 8.84505e-09 0 8.84805e-09 0.0007 8.85105e-09 0 8.90605e-09 0 8.90905e-09 0.0007 8.91205e-09 0 8.96705e-09 0 8.97005e-09 0.0007 8.97305e-09 0 9.02805e-09 0 9.03105e-09 0.0007 9.03405e-09 0 9.08905e-09 0 9.09205e-09 0.0007 9.09505e-09 0 9.15005e-09 0 9.15305e-09 0.0007 9.15605e-09 0 9.21105e-09 0 9.21405e-09 0.0007 9.21705e-09 0 9.27205e-09 0 9.27505e-09 0.0007 9.27805e-09 0 9.33305e-09 0 9.33605e-09 0.0007 9.33905e-09 0 9.39405e-09 0 9.39705e-09 0.0007 9.40005e-09 0 9.45505e-09 0 9.45805e-09 0.0007 9.46105e-09 0 9.51605e-09 0 9.51905e-09 0.0007 9.52205e-09 0 9.57705e-09 0 9.58005e-09 0.0007 9.58305e-09 0 9.63805e-09 0 9.64105e-09 0.0007 9.64405e-09 0 9.69905e-09 0 9.70205e-09 0.0007 9.70505e-09 0 9.76005e-09 0 9.76305e-09 0.0007 9.76605e-09 0 9.82105e-09 0 9.82405e-09 0.0007 9.82705e-09 0 9.88205e-09 0 9.88505e-09 0.0007 9.88805e-09 0 9.94305e-09 0 9.94605e-09 0.0007 9.94905e-09 0 1.0004e-08 0 1.0007e-08 0.0007 1.001e-08 0 1.0065e-08 0 1.0068e-08 0.0007 1.0071e-08 0 1.0126e-08 0 1.0129e-08 0.0007 1.0132e-08 0 1.0187e-08 0 1.019e-08 0.0007 1.01931e-08 0 1.0248e-08 0 1.0251e-08 0.0007 1.0254e-08 0 1.0309e-08 0 1.0312e-08 0.0007 1.0315e-08 0 1.037e-08 0 1.0373e-08 0.0007 1.0376e-08 0 1.0431e-08 0 1.0434e-08 0.0007 1.0437e-08 0 1.0492e-08 0 1.0495e-08 0.0007 1.0498e-08 0 1.0553e-08 0 1.0556e-08 0.0007 1.0559e-08 0 1.0614e-08 0 1.0617e-08 0.0007 1.062e-08 0 1.0675e-08 0 1.0678e-08 0.0007 1.0681e-08 0 1.0736e-08 0 1.0739e-08 0.0007 1.0742e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0858e-08 0 1.0861e-08 0.0007 1.0864e-08 0 1.0919e-08 0 1.0922e-08 0.0007 1.0925e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.1041e-08 0 1.1044e-08 0.0007 1.1047e-08 0 1.1102e-08 0 1.1105e-08 0.0007 1.1108e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1224e-08 0 1.1227e-08 0.0007 1.123e-08 0 1.1285e-08 0 1.1288e-08 0.0007 1.1291e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1468e-08 0 1.1471e-08 0.0007 1.1474e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.159e-08 0 1.1593e-08 0.0007 1.1596e-08 0 1.1651e-08 0 1.1654e-08 0.0007 1.1657e-08 0 1.1712e-08 0 1.1715e-08 0.0007 1.1718e-08 0 1.1773e-08 0 1.1776e-08 0.0007 1.1779e-08 0 1.1834e-08 0 1.1837e-08 0.0007 1.184e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.1956e-08 0 1.1959e-08 0.0007 1.1962e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2078e-08 0 1.2081e-08 0.0007 1.2084e-08 0 1.2139e-08 0 1.2142e-08 0.0007 1.2145e-08 0 1.22e-08 0 1.2203e-08 0.0007 1.2206e-08 0 1.2261e-08 0 1.2264e-08 0.0007 1.2267e-08 0 1.2322e-08 0 1.2325e-08 0.0007 1.2328e-08 0 1.2383e-08 0 1.2386e-08 0.0007 1.2389e-08 0 1.2444e-08 0 1.2447e-08 0.0007 1.245e-08 0 1.2505e-08 0 1.2508e-08 0.0007 1.2511e-08 0 1.2566e-08 0 1.2569e-08 0.0007 1.2572e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2688e-08 0 1.2691e-08 0.0007 1.2694e-08 0 1.2749e-08 0 1.2752e-08 0.0007 1.2755e-08 0 1.281e-08 0 1.2813e-08 0.0007 1.2816e-08 0 1.2871e-08 0 1.2874e-08 0.0007 1.2877e-08 0 1.2932e-08 0 1.2935e-08 0.0007 1.2938e-08 0 1.2993e-08 0 1.2996e-08 0.0007 1.2999e-08 0 1.3054e-08 0 1.3057e-08 0.0007 1.306e-08 0 1.3115e-08 0 1.3118e-08 0.0007 1.3121e-08 0 1.3176e-08 0 1.3179e-08 0.0007 1.3182e-08 0 1.3237e-08 0 1.324e-08 0.0007 1.3243e-08 0 1.3298e-08 0 1.3301e-08 0.0007 1.3304e-08 0 1.3359e-08 0 1.3362e-08 0.0007 1.3365e-08 0 1.342e-08 0 1.3423e-08 0.0007 1.3426e-08 0 1.3481e-08 0 1.3484e-08 0.0007 1.3487e-08 0 1.3542e-08 0 1.3545e-08 0.0007 1.3548e-08 0 1.3603e-08 0 1.3606e-08 0.0007 1.3609e-08 0 1.3664e-08 0 1.3667e-08 0.0007 1.367e-08 0 1.3725e-08 0 1.3728e-08 0.0007 1.3731e-08 0 1.3786e-08 0 1.3789e-08 0.0007 1.3792e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.3908e-08 0 1.3911e-08 0.0007 1.3914e-08 0 1.3969e-08 0 1.3972e-08 0.0007 1.3975e-08 0 1.403e-08 0 1.4033e-08 0.0007 1.4036e-08 0 1.4091e-08 0 1.4094e-08 0.0007 1.4097e-08 0 1.4152e-08 0 1.4155e-08 0.0007 1.4158e-08 0 1.4213e-08 0 1.4216e-08 0.0007 1.4219e-08 0 1.4274e-08 0 1.4277e-08 0.0007 1.428e-08 0 1.4335e-08 0 1.4338e-08 0.0007 1.4341e-08 0 1.4396e-08 0 1.4399e-08 0.0007 1.4402e-08 0 1.4457e-08 0 1.446e-08 0.0007 1.4463e-08 0 1.4518e-08 0 1.4521e-08 0.0007 1.4524e-08 0 1.4579e-08 0 1.4582e-08 0.0007 1.4585e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.4701e-08 0 1.4704e-08 0.0007 1.4707e-08 0 1.4762e-08 0 1.4765e-08 0.0007 1.4768e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4884e-08 0 1.4887e-08 0.0007 1.489e-08 0 1.4945e-08 0 1.4948e-08 0.0007 1.4951e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5067e-08 0 1.507e-08 0.0007 1.5073e-08 0 1.5128e-08 0 1.5131e-08 0.0007 1.5134e-08 0 1.5189e-08 0 1.5192e-08 0.0007 1.5195e-08 0 1.52501e-08 0 1.52531e-08 0.0007 1.52561e-08 0 1.5311e-08 0 1.53141e-08 0.0007 1.53171e-08 0 1.5372e-08 0 1.5375e-08 0.0007 1.5378e-08 0 1.5433e-08 0 1.5436e-08 0.0007 1.5439e-08 0 1.5494e-08 0 1.5497e-08 0.0007 1.55e-08 0 1.5555e-08 0 1.5558e-08 0.0007 1.5561e-08 0 1.5616e-08 0 1.5619e-08 0.0007 1.5622e-08 0 1.5677e-08 0 1.568e-08 0.0007 1.5683e-08 0 1.5738e-08 0 1.5741e-08 0.0007 1.5744e-08 0 1.5799e-08 0 1.5802e-08 0.0007 1.5805e-08 0 1.586e-08 0 1.5863e-08 0.0007 1.5866e-08 0 1.59211e-08 0 1.59241e-08 0.0007 1.59271e-08 0 1.5982e-08 0 1.5985e-08 0.0007 1.59881e-08 0 1.6043e-08 0 1.6046e-08 0.0007 1.6049e-08 0 1.6104e-08 0 1.6107e-08 0.0007 1.611e-08 0 1.6165e-08 0 1.6168e-08 0.0007 1.6171e-08 0 1.6226e-08 0 1.6229e-08 0.0007 1.6232e-08 0 1.6287e-08 0 1.629e-08 0.0007 1.6293e-08 0 1.6348e-08 0 1.6351e-08 0.0007 1.6354e-08 0 1.6409e-08 0 1.6412e-08 0.0007 1.6415e-08 0 1.647e-08 0 1.6473e-08 0.0007 1.6476e-08 0 1.65311e-08 0 1.65341e-08 0.0007 1.65371e-08 0 1.65921e-08 0 1.65951e-08 0.0007 1.65981e-08 0 1.6653e-08 0 1.6656e-08 0.0007 1.6659e-08 0 1.6714e-08 0 1.6717e-08 0.0007 1.672e-08 0 1.6775e-08 0 1.6778e-08 0.0007 1.6781e-08 0 1.6836e-08 0 1.6839e-08 0.0007 1.6842e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6958e-08 0 1.6961e-08 0.0007 1.6964e-08 0 1.7019e-08 0 1.7022e-08 0.0007 1.7025e-08 0 1.708e-08 0 1.7083e-08 0.0007 1.7086e-08 0 1.7141e-08 0 1.7144e-08 0.0007 1.7147e-08 0 1.72021e-08 0 1.72051e-08 0.0007 1.72081e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.72691e-08 0 1.7324e-08 0 1.7327e-08 0.0007 1.733e-08 0 1.7385e-08 0 1.7388e-08 0.0007 1.7391e-08 0 1.7446e-08 0 1.7449e-08 0.0007 1.7452e-08 0 1.7507e-08 0 1.751e-08 0.0007 1.7513e-08 0 1.7568e-08 0 1.7571e-08 0.0007 1.7574e-08 0 1.7629e-08 0 1.7632e-08 0.0007 1.7635e-08 0 1.769e-08 0 1.7693e-08 0.0007 1.7696e-08 0 1.7751e-08 0 1.7754e-08 0.0007 1.7757e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.78731e-08 0 1.78761e-08 0.0007 1.78791e-08 0 1.7934e-08 0 1.7937e-08 0.0007 1.794e-08 0 1.7995e-08 0 1.7998e-08 0.0007 1.8001e-08 0 1.8056e-08 0 1.8059e-08 0.0007 1.8062e-08 0 1.8117e-08 0 1.812e-08 0.0007 1.8123e-08 0 1.8178e-08 0 1.8181e-08 0.0007 1.8184e-08 0 1.8239e-08 0 1.8242e-08 0.0007 1.8245e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.8361e-08 0 1.8364e-08 0.0007 1.8367e-08 0 1.8422e-08 0 1.8425e-08 0.0007 1.8428e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8544e-08 0 1.8547e-08 0.0007 1.85501e-08 0 1.8605e-08 0 1.8608e-08 0.0007 1.8611e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8727e-08 0 1.873e-08 0.0007 1.8733e-08 0 1.8788e-08 0 1.8791e-08 0.0007 1.8794e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.891e-08 0 1.8913e-08 0.0007 1.8916e-08 0 1.8971e-08 0 1.8974e-08 0.0007 1.8977e-08 0 1.9032e-08 0 1.9035e-08 0.0007 1.9038e-08 0 1.9093e-08 0 1.9096e-08 0.0007 1.9099e-08 0 1.91541e-08 0 1.91571e-08 0.0007 1.91601e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9276e-08 0 1.9279e-08 0.0007 1.9282e-08 0 1.9337e-08 0 1.934e-08 0.0007 1.9343e-08 0 1.9398e-08 0 1.9401e-08 0.0007 1.9404e-08 0 1.9459e-08 0 1.9462e-08 0.0007 1.9465e-08 0 1.952e-08 0 1.9523e-08 0.0007 1.9526e-08 0 1.9581e-08 0 1.9584e-08 0.0007 1.9587e-08 0 1.9642e-08 0 1.9645e-08 0.0007 1.9648e-08 0 1.9703e-08 0 1.9706e-08 0.0007 1.9709e-08 0 1.9764e-08 0 1.9767e-08 0.0007 1.977e-08 0 1.9825e-08 0 1.9828e-08 0.0007 1.98311e-08 0 1.9886e-08 0 1.9889e-08 0.0007 1.9892e-08 0 1.9947e-08 0 1.995e-08 0.0007 1.9953e-08 0 2.0008e-08 0 2.0011e-08 0.0007 2.0014e-08 0 2.0069e-08 0 2.0072e-08 0.0007 2.0075e-08 0 2.013e-08 0 2.0133e-08 0.0007 2.0136e-08 0 2.0191e-08 0 2.0194e-08 0.0007 2.0197e-08 0 2.0252e-08 0 2.0255e-08 0.0007 2.0258e-08 0 2.0313e-08 0 2.0316e-08 0.0007 2.0319e-08 0 2.0374e-08 0 2.0377e-08 0.0007 2.038e-08 0 2.04351e-08 0 2.04381e-08 0.0007 2.04411e-08 0 2.0496e-08 0 2.0499e-08 0.0007 2.0502e-08 0 2.0557e-08 0 2.056e-08 0.0007 2.0563e-08 0 2.0618e-08 0 2.0621e-08 0.0007 2.0624e-08 0 2.0679e-08 0 2.0682e-08 0.0007 2.0685e-08 0 2.074e-08 0 2.0743e-08 0.0007 2.0746e-08 0 2.0801e-08 0 2.0804e-08 0.0007 2.0807e-08 0 2.0862e-08 0 2.0865e-08 0.0007 2.0868e-08 0 2.0923e-08 0 2.0926e-08 0.0007 2.0929e-08 0 2.0984e-08 0 2.0987e-08 0.0007 2.099e-08 0 2.1045e-08 0 2.1048e-08 0.0007 2.1051e-08 0 2.1106e-08 0 2.11091e-08 0.0007 2.11121e-08 0 2.1167e-08 0 2.117e-08 0.0007 2.1173e-08 0 2.1228e-08 0 2.1231e-08 0.0007 2.1234e-08 0 2.1289e-08 0 2.1292e-08 0.0007 2.1295e-08 0 2.135e-08 0 2.1353e-08 0.0007 2.1356e-08 0 2.1411e-08 0 2.1414e-08 0.0007 2.1417e-08 0 2.1472e-08 0 2.1475e-08 0.0007 2.1478e-08 0 2.1533e-08 0 2.1536e-08 0.0007 2.1539e-08 0 2.1594e-08 0 2.1597e-08 0.0007 2.16e-08 0 2.1655e-08 0 2.1658e-08 0.0007 2.1661e-08 0 2.1716e-08 0 2.1719e-08 0.0007 2.1722e-08 0 2.1777e-08 0 2.178e-08 0.0007 2.1783e-08 0 2.1838e-08 0 2.1841e-08 0.0007 2.1844e-08 0 2.1899e-08 0 2.1902e-08 0.0007 2.1905e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.2021e-08 0 2.2024e-08 0.0007 2.2027e-08 0 2.2082e-08 0 2.2085e-08 0.0007 2.2088e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2204e-08 0 2.2207e-08 0.0007 2.221e-08 0 2.2265e-08 0 2.2268e-08 0.0007 2.2271e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2448e-08 0 2.2451e-08 0.0007 2.2454e-08 0 2.2509e-08 0 2.2512e-08 0.0007 2.2515e-08 0 2.257e-08 0 2.2573e-08 0.0007 2.2576e-08 0 2.2631e-08 0 2.2634e-08 0.0007 2.2637e-08 0 2.2692e-08 0 2.2695e-08 0.0007 2.2698e-08 0 2.2753e-08 0 2.2756e-08 0.0007 2.2759e-08 0 2.2814e-08 0 2.2817e-08 0.0007 2.282e-08 0 2.2875e-08 0 2.2878e-08 0.0007 2.2881e-08 0 2.2936e-08 0 2.2939e-08 0.0007 2.2942e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3058e-08 0 2.3061e-08 0.0007 2.3064e-08 0 2.3119e-08 0 2.3122e-08 0.0007 2.3125e-08 0 2.318e-08 0 2.3183e-08 0.0007 2.3186e-08 0 2.3241e-08 0 2.3244e-08 0.0007 2.3247e-08 0 2.3302e-08 0 2.3305e-08 0.0007 2.3308e-08 0 2.3363e-08 0 2.3366e-08 0.0007 2.3369e-08 0 2.3424e-08 0 2.3427e-08 0.0007 2.343e-08 0 2.3485e-08 0 2.3488e-08 0.0007 2.3491e-08 0 2.3546e-08 0 2.3549e-08 0.0007 2.3552e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3668e-08 0 2.3671e-08 0.0007 2.3674e-08 0 2.3729e-08 0 2.3732e-08 0.0007 2.3735e-08 0 2.379e-08 0 2.3793e-08 0.0007 2.3796e-08 0 2.3851e-08 0 2.3854e-08 0.0007 2.3857e-08 0 2.3912e-08 0 2.3915e-08 0.0007 2.3918e-08 0 2.3973e-08 0 2.3976e-08 0.0007 2.3979e-08 0 2.4034e-08 0 2.4037e-08 0.0007 2.404e-08 0 2.4095e-08 0 2.4098e-08 0.0007 2.4101e-08 0 2.4156e-08 0 2.4159e-08 0.0007 2.4162e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4278e-08 0 2.4281e-08 0.0007 2.4284e-08 0)
L_S0|1 P0_2_RX _S0|A1  2.067833848e-12
L_S0|2 _S0|A1 _S0|A2  4.135667696e-12
L_S0|3 _S0|A3 _S0|A4  8.271335392e-12
L_S0|T T12 _S0|T1  2.067833848e-12
L_S0|4 _S0|T1 _S0|T2  4.135667696e-12
L_S0|5 _S0|A4 _S0|Q1  4.135667696e-12
L_S0|6 _S0|Q1 S0  2.067833848e-12
IT13|T 0 T13  PWL(0 0 5e-14 0 3.05e-12 0.0007 6.05e-12 0 6.105e-11 0 6.405e-11 0.0007 6.705e-11 0 1.2205e-10 0 1.2505e-10 0.0007 1.2805e-10 0 1.8305e-10 0 1.8605e-10 0.0007 1.8905e-10 0 2.4405e-10 0 2.4705e-10 0.0007 2.5005e-10 0 3.0505e-10 0 3.0805e-10 0.0007 3.1105e-10 0 3.6605e-10 0 3.6905e-10 0.0007 3.7205e-10 0 4.2705e-10 0 4.3005e-10 0.0007 4.3305e-10 0 4.8805e-10 0 4.9105e-10 0.0007 4.9405e-10 0 5.4905e-10 0 5.5205e-10 0.0007 5.5505e-10 0 6.1005e-10 0 6.1305e-10 0.0007 6.1605e-10 0 6.7105e-10 0 6.7405e-10 0.0007 6.7705e-10 0 7.3205e-10 0 7.3505e-10 0.0007 7.3805e-10 0 7.9305e-10 0 7.9605e-10 0.0007 7.9905e-10 0 8.5405e-10 0 8.5705e-10 0.0007 8.6005e-10 0 9.1505e-10 0 9.1805e-10 0.0007 9.2105e-10 0 9.7605e-10 0 9.7905e-10 0.0007 9.8205e-10 0 1.03705e-09 0 1.04005e-09 0.0007 1.04305e-09 0 1.09805e-09 0 1.10105e-09 0.0007 1.10405e-09 0 1.15905e-09 0 1.16205e-09 0.0007 1.16505e-09 0 1.22005e-09 0 1.22305e-09 0.0007 1.22605e-09 0 1.28105e-09 0 1.28405e-09 0.0007 1.28705e-09 0 1.34205e-09 0 1.34505e-09 0.0007 1.34805e-09 0 1.40305e-09 0 1.40605e-09 0.0007 1.40905e-09 0 1.46405e-09 0 1.46705e-09 0.0007 1.47005e-09 0 1.52505e-09 0 1.52805e-09 0.0007 1.53105e-09 0 1.58605e-09 0 1.58905e-09 0.0007 1.59205e-09 0 1.64705e-09 0 1.65005e-09 0.0007 1.65305e-09 0 1.70805e-09 0 1.71105e-09 0.0007 1.71405e-09 0 1.76905e-09 0 1.77205e-09 0.0007 1.77505e-09 0 1.83005e-09 0 1.83305e-09 0.0007 1.83605e-09 0 1.89105e-09 0 1.89405e-09 0.0007 1.89705e-09 0 1.95205e-09 0 1.95505e-09 0.0007 1.95805e-09 0 2.01305e-09 0 2.01605e-09 0.0007 2.01905e-09 0 2.07405e-09 0 2.07705e-09 0.0007 2.08005e-09 0 2.13505e-09 0 2.13805e-09 0.0007 2.14105e-09 0 2.19605e-09 0 2.19905e-09 0.0007 2.20205e-09 0 2.25705e-09 0 2.26005e-09 0.0007 2.26305e-09 0 2.31805e-09 0 2.32105e-09 0.0007 2.32405e-09 0 2.37905e-09 0 2.38205e-09 0.0007 2.38505e-09 0 2.44005e-09 0 2.44305e-09 0.0007 2.44605e-09 0 2.50105e-09 0 2.50405e-09 0.0007 2.50705e-09 0 2.56205e-09 0 2.56505e-09 0.0007 2.56805e-09 0 2.62305e-09 0 2.62605e-09 0.0007 2.62905e-09 0 2.68405e-09 0 2.68705e-09 0.0007 2.69005e-09 0 2.74505e-09 0 2.74805e-09 0.0007 2.75105e-09 0 2.80605e-09 0 2.80905e-09 0.0007 2.81205e-09 0 2.86705e-09 0 2.87005e-09 0.0007 2.87305e-09 0 2.92805e-09 0 2.93105e-09 0.0007 2.93405e-09 0 2.98905e-09 0 2.99205e-09 0.0007 2.99505e-09 0 3.05005e-09 0 3.05305e-09 0.0007 3.05605e-09 0 3.11105e-09 0 3.11405e-09 0.0007 3.11705e-09 0 3.17205e-09 0 3.17505e-09 0.0007 3.17805e-09 0 3.23305e-09 0 3.23605e-09 0.0007 3.23905e-09 0 3.29405e-09 0 3.29705e-09 0.0007 3.30005e-09 0 3.35505e-09 0 3.35805e-09 0.0007 3.36105e-09 0 3.41605e-09 0 3.41905e-09 0.0007 3.42205e-09 0 3.47705e-09 0 3.48005e-09 0.0007 3.48305e-09 0 3.53805e-09 0 3.54105e-09 0.0007 3.54405e-09 0 3.59905e-09 0 3.60205e-09 0.0007 3.60505e-09 0 3.66005e-09 0 3.66305e-09 0.0007 3.66605e-09 0 3.72105e-09 0 3.72405e-09 0.0007 3.72705e-09 0 3.78205e-09 0 3.78505e-09 0.0007 3.78805e-09 0 3.84305e-09 0 3.84605e-09 0.0007 3.84905e-09 0 3.90405e-09 0 3.90705e-09 0.0007 3.91005e-09 0 3.96505e-09 0 3.96805e-09 0.0007 3.97105e-09 0 4.02605e-09 0 4.02905e-09 0.0007 4.03205e-09 0 4.08705e-09 0 4.09005e-09 0.0007 4.09305e-09 0 4.14805e-09 0 4.15105e-09 0.0007 4.15405e-09 0 4.20905e-09 0 4.21205e-09 0.0007 4.21505e-09 0 4.27005e-09 0 4.27305e-09 0.0007 4.27605e-09 0 4.33105e-09 0 4.33405e-09 0.0007 4.33705e-09 0 4.39205e-09 0 4.39505e-09 0.0007 4.39805e-09 0 4.45305e-09 0 4.45605e-09 0.0007 4.45905e-09 0 4.51405e-09 0 4.51705e-09 0.0007 4.52005e-09 0 4.57505e-09 0 4.57805e-09 0.0007 4.58105e-09 0 4.63605e-09 0 4.63905e-09 0.0007 4.64205e-09 0 4.69705e-09 0 4.70005e-09 0.0007 4.70305e-09 0 4.75805e-09 0 4.76105e-09 0.0007 4.76405e-09 0 4.81905e-09 0 4.82205e-09 0.0007 4.82505e-09 0 4.88005e-09 0 4.88305e-09 0.0007 4.88605e-09 0 4.94105e-09 0 4.94405e-09 0.0007 4.94705e-09 0 5.00205e-09 0 5.00505e-09 0.0007 5.00805e-09 0 5.06305e-09 0 5.06605e-09 0.0007 5.06905e-09 0 5.12405e-09 0 5.12705e-09 0.0007 5.13005e-09 0 5.18505e-09 0 5.18805e-09 0.0007 5.19105e-09 0 5.24605e-09 0 5.24905e-09 0.0007 5.25205e-09 0 5.30705e-09 0 5.31005e-09 0.0007 5.31305e-09 0 5.36805e-09 0 5.37105e-09 0.0007 5.37405e-09 0 5.42905e-09 0 5.43205e-09 0.0007 5.43505e-09 0 5.49005e-09 0 5.49305e-09 0.0007 5.49605e-09 0 5.55105e-09 0 5.55405e-09 0.0007 5.55705e-09 0 5.61205e-09 0 5.61505e-09 0.0007 5.61805e-09 0 5.67305e-09 0 5.67605e-09 0.0007 5.67905e-09 0 5.73405e-09 0 5.73705e-09 0.0007 5.74005e-09 0 5.79505e-09 0 5.79805e-09 0.0007 5.80105e-09 0 5.85605e-09 0 5.85905e-09 0.0007 5.86205e-09 0 5.91705e-09 0 5.92005e-09 0.0007 5.92305e-09 0 5.97805e-09 0 5.98105e-09 0.0007 5.98405e-09 0 6.03905e-09 0 6.04205e-09 0.0007 6.04505e-09 0 6.10005e-09 0 6.10305e-09 0.0007 6.10605e-09 0 6.16105e-09 0 6.16405e-09 0.0007 6.16705e-09 0 6.22205e-09 0 6.22505e-09 0.0007 6.22805e-09 0 6.28305e-09 0 6.28605e-09 0.0007 6.28905e-09 0 6.34405e-09 0 6.34705e-09 0.0007 6.35005e-09 0 6.40505e-09 0 6.40805e-09 0.0007 6.41105e-09 0 6.46605e-09 0 6.46905e-09 0.0007 6.47205e-09 0 6.52705e-09 0 6.53005e-09 0.0007 6.53305e-09 0 6.58805e-09 0 6.59105e-09 0.0007 6.59405e-09 0 6.64905e-09 0 6.65205e-09 0.0007 6.65505e-09 0 6.71005e-09 0 6.71305e-09 0.0007 6.71605e-09 0 6.77105e-09 0 6.77405e-09 0.0007 6.77705e-09 0 6.83205e-09 0 6.83505e-09 0.0007 6.83805e-09 0 6.89305e-09 0 6.89605e-09 0.0007 6.89905e-09 0 6.95405e-09 0 6.95705e-09 0.0007 6.96005e-09 0 7.01505e-09 0 7.01805e-09 0.0007 7.02105e-09 0 7.07605e-09 0 7.07905e-09 0.0007 7.08205e-09 0 7.13705e-09 0 7.14005e-09 0.0007 7.14305e-09 0 7.19805e-09 0 7.20105e-09 0.0007 7.20405e-09 0 7.25905e-09 0 7.26205e-09 0.0007 7.26505e-09 0 7.32005e-09 0 7.32305e-09 0.0007 7.32605e-09 0 7.38105e-09 0 7.38405e-09 0.0007 7.38705e-09 0 7.44205e-09 0 7.44505e-09 0.0007 7.44805e-09 0 7.50305e-09 0 7.50605e-09 0.0007 7.50905e-09 0 7.56405e-09 0 7.56705e-09 0.0007 7.57005e-09 0 7.62505e-09 0 7.62805e-09 0.0007 7.63105e-09 0 7.68605e-09 0 7.68905e-09 0.0007 7.69205e-09 0 7.74705e-09 0 7.75005e-09 0.0007 7.75305e-09 0 7.80805e-09 0 7.81105e-09 0.0007 7.81405e-09 0 7.86905e-09 0 7.87205e-09 0.0007 7.87505e-09 0 7.93005e-09 0 7.93305e-09 0.0007 7.93605e-09 0 7.99105e-09 0 7.99405e-09 0.0007 7.99705e-09 0 8.05205e-09 0 8.05505e-09 0.0007 8.05805e-09 0 8.11305e-09 0 8.11605e-09 0.0007 8.11905e-09 0 8.17405e-09 0 8.17705e-09 0.0007 8.18005e-09 0 8.23505e-09 0 8.23805e-09 0.0007 8.24105e-09 0 8.29605e-09 0 8.29905e-09 0.0007 8.30205e-09 0 8.35705e-09 0 8.36005e-09 0.0007 8.36305e-09 0 8.41805e-09 0 8.42105e-09 0.0007 8.42405e-09 0 8.47905e-09 0 8.48205e-09 0.0007 8.48505e-09 0 8.54005e-09 0 8.54305e-09 0.0007 8.54605e-09 0 8.60105e-09 0 8.60405e-09 0.0007 8.60705e-09 0 8.66205e-09 0 8.66505e-09 0.0007 8.66805e-09 0 8.72305e-09 0 8.72605e-09 0.0007 8.72905e-09 0 8.78405e-09 0 8.78705e-09 0.0007 8.79005e-09 0 8.84505e-09 0 8.84805e-09 0.0007 8.85105e-09 0 8.90605e-09 0 8.90905e-09 0.0007 8.91205e-09 0 8.96705e-09 0 8.97005e-09 0.0007 8.97305e-09 0 9.02805e-09 0 9.03105e-09 0.0007 9.03405e-09 0 9.08905e-09 0 9.09205e-09 0.0007 9.09505e-09 0 9.15005e-09 0 9.15305e-09 0.0007 9.15605e-09 0 9.21105e-09 0 9.21405e-09 0.0007 9.21705e-09 0 9.27205e-09 0 9.27505e-09 0.0007 9.27805e-09 0 9.33305e-09 0 9.33605e-09 0.0007 9.33905e-09 0 9.39405e-09 0 9.39705e-09 0.0007 9.40005e-09 0 9.45505e-09 0 9.45805e-09 0.0007 9.46105e-09 0 9.51605e-09 0 9.51905e-09 0.0007 9.52205e-09 0 9.57705e-09 0 9.58005e-09 0.0007 9.58305e-09 0 9.63805e-09 0 9.64105e-09 0.0007 9.64405e-09 0 9.69905e-09 0 9.70205e-09 0.0007 9.70505e-09 0 9.76005e-09 0 9.76305e-09 0.0007 9.76605e-09 0 9.82105e-09 0 9.82405e-09 0.0007 9.82705e-09 0 9.88205e-09 0 9.88505e-09 0.0007 9.88805e-09 0 9.94305e-09 0 9.94605e-09 0.0007 9.94905e-09 0 1.0004e-08 0 1.0007e-08 0.0007 1.001e-08 0 1.0065e-08 0 1.0068e-08 0.0007 1.0071e-08 0 1.0126e-08 0 1.0129e-08 0.0007 1.0132e-08 0 1.0187e-08 0 1.019e-08 0.0007 1.01931e-08 0 1.0248e-08 0 1.0251e-08 0.0007 1.0254e-08 0 1.0309e-08 0 1.0312e-08 0.0007 1.0315e-08 0 1.037e-08 0 1.0373e-08 0.0007 1.0376e-08 0 1.0431e-08 0 1.0434e-08 0.0007 1.0437e-08 0 1.0492e-08 0 1.0495e-08 0.0007 1.0498e-08 0 1.0553e-08 0 1.0556e-08 0.0007 1.0559e-08 0 1.0614e-08 0 1.0617e-08 0.0007 1.062e-08 0 1.0675e-08 0 1.0678e-08 0.0007 1.0681e-08 0 1.0736e-08 0 1.0739e-08 0.0007 1.0742e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0858e-08 0 1.0861e-08 0.0007 1.0864e-08 0 1.0919e-08 0 1.0922e-08 0.0007 1.0925e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.1041e-08 0 1.1044e-08 0.0007 1.1047e-08 0 1.1102e-08 0 1.1105e-08 0.0007 1.1108e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1224e-08 0 1.1227e-08 0.0007 1.123e-08 0 1.1285e-08 0 1.1288e-08 0.0007 1.1291e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1468e-08 0 1.1471e-08 0.0007 1.1474e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.159e-08 0 1.1593e-08 0.0007 1.1596e-08 0 1.1651e-08 0 1.1654e-08 0.0007 1.1657e-08 0 1.1712e-08 0 1.1715e-08 0.0007 1.1718e-08 0 1.1773e-08 0 1.1776e-08 0.0007 1.1779e-08 0 1.1834e-08 0 1.1837e-08 0.0007 1.184e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.1956e-08 0 1.1959e-08 0.0007 1.1962e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2078e-08 0 1.2081e-08 0.0007 1.2084e-08 0 1.2139e-08 0 1.2142e-08 0.0007 1.2145e-08 0 1.22e-08 0 1.2203e-08 0.0007 1.2206e-08 0 1.2261e-08 0 1.2264e-08 0.0007 1.2267e-08 0 1.2322e-08 0 1.2325e-08 0.0007 1.2328e-08 0 1.2383e-08 0 1.2386e-08 0.0007 1.2389e-08 0 1.2444e-08 0 1.2447e-08 0.0007 1.245e-08 0 1.2505e-08 0 1.2508e-08 0.0007 1.2511e-08 0 1.2566e-08 0 1.2569e-08 0.0007 1.2572e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2688e-08 0 1.2691e-08 0.0007 1.2694e-08 0 1.2749e-08 0 1.2752e-08 0.0007 1.2755e-08 0 1.281e-08 0 1.2813e-08 0.0007 1.2816e-08 0 1.2871e-08 0 1.2874e-08 0.0007 1.2877e-08 0 1.2932e-08 0 1.2935e-08 0.0007 1.2938e-08 0 1.2993e-08 0 1.2996e-08 0.0007 1.2999e-08 0 1.3054e-08 0 1.3057e-08 0.0007 1.306e-08 0 1.3115e-08 0 1.3118e-08 0.0007 1.3121e-08 0 1.3176e-08 0 1.3179e-08 0.0007 1.3182e-08 0 1.3237e-08 0 1.324e-08 0.0007 1.3243e-08 0 1.3298e-08 0 1.3301e-08 0.0007 1.3304e-08 0 1.3359e-08 0 1.3362e-08 0.0007 1.3365e-08 0 1.342e-08 0 1.3423e-08 0.0007 1.3426e-08 0 1.3481e-08 0 1.3484e-08 0.0007 1.3487e-08 0 1.3542e-08 0 1.3545e-08 0.0007 1.3548e-08 0 1.3603e-08 0 1.3606e-08 0.0007 1.3609e-08 0 1.3664e-08 0 1.3667e-08 0.0007 1.367e-08 0 1.3725e-08 0 1.3728e-08 0.0007 1.3731e-08 0 1.3786e-08 0 1.3789e-08 0.0007 1.3792e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.3908e-08 0 1.3911e-08 0.0007 1.3914e-08 0 1.3969e-08 0 1.3972e-08 0.0007 1.3975e-08 0 1.403e-08 0 1.4033e-08 0.0007 1.4036e-08 0 1.4091e-08 0 1.4094e-08 0.0007 1.4097e-08 0 1.4152e-08 0 1.4155e-08 0.0007 1.4158e-08 0 1.4213e-08 0 1.4216e-08 0.0007 1.4219e-08 0 1.4274e-08 0 1.4277e-08 0.0007 1.428e-08 0 1.4335e-08 0 1.4338e-08 0.0007 1.4341e-08 0 1.4396e-08 0 1.4399e-08 0.0007 1.4402e-08 0 1.4457e-08 0 1.446e-08 0.0007 1.4463e-08 0 1.4518e-08 0 1.4521e-08 0.0007 1.4524e-08 0 1.4579e-08 0 1.4582e-08 0.0007 1.4585e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.4701e-08 0 1.4704e-08 0.0007 1.4707e-08 0 1.4762e-08 0 1.4765e-08 0.0007 1.4768e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4884e-08 0 1.4887e-08 0.0007 1.489e-08 0 1.4945e-08 0 1.4948e-08 0.0007 1.4951e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5067e-08 0 1.507e-08 0.0007 1.5073e-08 0 1.5128e-08 0 1.5131e-08 0.0007 1.5134e-08 0 1.5189e-08 0 1.5192e-08 0.0007 1.5195e-08 0 1.52501e-08 0 1.52531e-08 0.0007 1.52561e-08 0 1.5311e-08 0 1.53141e-08 0.0007 1.53171e-08 0 1.5372e-08 0 1.5375e-08 0.0007 1.5378e-08 0 1.5433e-08 0 1.5436e-08 0.0007 1.5439e-08 0 1.5494e-08 0 1.5497e-08 0.0007 1.55e-08 0 1.5555e-08 0 1.5558e-08 0.0007 1.5561e-08 0 1.5616e-08 0 1.5619e-08 0.0007 1.5622e-08 0 1.5677e-08 0 1.568e-08 0.0007 1.5683e-08 0 1.5738e-08 0 1.5741e-08 0.0007 1.5744e-08 0 1.5799e-08 0 1.5802e-08 0.0007 1.5805e-08 0 1.586e-08 0 1.5863e-08 0.0007 1.5866e-08 0 1.59211e-08 0 1.59241e-08 0.0007 1.59271e-08 0 1.5982e-08 0 1.5985e-08 0.0007 1.59881e-08 0 1.6043e-08 0 1.6046e-08 0.0007 1.6049e-08 0 1.6104e-08 0 1.6107e-08 0.0007 1.611e-08 0 1.6165e-08 0 1.6168e-08 0.0007 1.6171e-08 0 1.6226e-08 0 1.6229e-08 0.0007 1.6232e-08 0 1.6287e-08 0 1.629e-08 0.0007 1.6293e-08 0 1.6348e-08 0 1.6351e-08 0.0007 1.6354e-08 0 1.6409e-08 0 1.6412e-08 0.0007 1.6415e-08 0 1.647e-08 0 1.6473e-08 0.0007 1.6476e-08 0 1.65311e-08 0 1.65341e-08 0.0007 1.65371e-08 0 1.65921e-08 0 1.65951e-08 0.0007 1.65981e-08 0 1.6653e-08 0 1.6656e-08 0.0007 1.6659e-08 0 1.6714e-08 0 1.6717e-08 0.0007 1.672e-08 0 1.6775e-08 0 1.6778e-08 0.0007 1.6781e-08 0 1.6836e-08 0 1.6839e-08 0.0007 1.6842e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6958e-08 0 1.6961e-08 0.0007 1.6964e-08 0 1.7019e-08 0 1.7022e-08 0.0007 1.7025e-08 0 1.708e-08 0 1.7083e-08 0.0007 1.7086e-08 0 1.7141e-08 0 1.7144e-08 0.0007 1.7147e-08 0 1.72021e-08 0 1.72051e-08 0.0007 1.72081e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.72691e-08 0 1.7324e-08 0 1.7327e-08 0.0007 1.733e-08 0 1.7385e-08 0 1.7388e-08 0.0007 1.7391e-08 0 1.7446e-08 0 1.7449e-08 0.0007 1.7452e-08 0 1.7507e-08 0 1.751e-08 0.0007 1.7513e-08 0 1.7568e-08 0 1.7571e-08 0.0007 1.7574e-08 0 1.7629e-08 0 1.7632e-08 0.0007 1.7635e-08 0 1.769e-08 0 1.7693e-08 0.0007 1.7696e-08 0 1.7751e-08 0 1.7754e-08 0.0007 1.7757e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.78731e-08 0 1.78761e-08 0.0007 1.78791e-08 0 1.7934e-08 0 1.7937e-08 0.0007 1.794e-08 0 1.7995e-08 0 1.7998e-08 0.0007 1.8001e-08 0 1.8056e-08 0 1.8059e-08 0.0007 1.8062e-08 0 1.8117e-08 0 1.812e-08 0.0007 1.8123e-08 0 1.8178e-08 0 1.8181e-08 0.0007 1.8184e-08 0 1.8239e-08 0 1.8242e-08 0.0007 1.8245e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.8361e-08 0 1.8364e-08 0.0007 1.8367e-08 0 1.8422e-08 0 1.8425e-08 0.0007 1.8428e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8544e-08 0 1.8547e-08 0.0007 1.85501e-08 0 1.8605e-08 0 1.8608e-08 0.0007 1.8611e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8727e-08 0 1.873e-08 0.0007 1.8733e-08 0 1.8788e-08 0 1.8791e-08 0.0007 1.8794e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.891e-08 0 1.8913e-08 0.0007 1.8916e-08 0 1.8971e-08 0 1.8974e-08 0.0007 1.8977e-08 0 1.9032e-08 0 1.9035e-08 0.0007 1.9038e-08 0 1.9093e-08 0 1.9096e-08 0.0007 1.9099e-08 0 1.91541e-08 0 1.91571e-08 0.0007 1.91601e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9276e-08 0 1.9279e-08 0.0007 1.9282e-08 0 1.9337e-08 0 1.934e-08 0.0007 1.9343e-08 0 1.9398e-08 0 1.9401e-08 0.0007 1.9404e-08 0 1.9459e-08 0 1.9462e-08 0.0007 1.9465e-08 0 1.952e-08 0 1.9523e-08 0.0007 1.9526e-08 0 1.9581e-08 0 1.9584e-08 0.0007 1.9587e-08 0 1.9642e-08 0 1.9645e-08 0.0007 1.9648e-08 0 1.9703e-08 0 1.9706e-08 0.0007 1.9709e-08 0 1.9764e-08 0 1.9767e-08 0.0007 1.977e-08 0 1.9825e-08 0 1.9828e-08 0.0007 1.98311e-08 0 1.9886e-08 0 1.9889e-08 0.0007 1.9892e-08 0 1.9947e-08 0 1.995e-08 0.0007 1.9953e-08 0 2.0008e-08 0 2.0011e-08 0.0007 2.0014e-08 0 2.0069e-08 0 2.0072e-08 0.0007 2.0075e-08 0 2.013e-08 0 2.0133e-08 0.0007 2.0136e-08 0 2.0191e-08 0 2.0194e-08 0.0007 2.0197e-08 0 2.0252e-08 0 2.0255e-08 0.0007 2.0258e-08 0 2.0313e-08 0 2.0316e-08 0.0007 2.0319e-08 0 2.0374e-08 0 2.0377e-08 0.0007 2.038e-08 0 2.04351e-08 0 2.04381e-08 0.0007 2.04411e-08 0 2.0496e-08 0 2.0499e-08 0.0007 2.0502e-08 0 2.0557e-08 0 2.056e-08 0.0007 2.0563e-08 0 2.0618e-08 0 2.0621e-08 0.0007 2.0624e-08 0 2.0679e-08 0 2.0682e-08 0.0007 2.0685e-08 0 2.074e-08 0 2.0743e-08 0.0007 2.0746e-08 0 2.0801e-08 0 2.0804e-08 0.0007 2.0807e-08 0 2.0862e-08 0 2.0865e-08 0.0007 2.0868e-08 0 2.0923e-08 0 2.0926e-08 0.0007 2.0929e-08 0 2.0984e-08 0 2.0987e-08 0.0007 2.099e-08 0 2.1045e-08 0 2.1048e-08 0.0007 2.1051e-08 0 2.1106e-08 0 2.11091e-08 0.0007 2.11121e-08 0 2.1167e-08 0 2.117e-08 0.0007 2.1173e-08 0 2.1228e-08 0 2.1231e-08 0.0007 2.1234e-08 0 2.1289e-08 0 2.1292e-08 0.0007 2.1295e-08 0 2.135e-08 0 2.1353e-08 0.0007 2.1356e-08 0 2.1411e-08 0 2.1414e-08 0.0007 2.1417e-08 0 2.1472e-08 0 2.1475e-08 0.0007 2.1478e-08 0 2.1533e-08 0 2.1536e-08 0.0007 2.1539e-08 0 2.1594e-08 0 2.1597e-08 0.0007 2.16e-08 0 2.1655e-08 0 2.1658e-08 0.0007 2.1661e-08 0 2.1716e-08 0 2.1719e-08 0.0007 2.1722e-08 0 2.1777e-08 0 2.178e-08 0.0007 2.1783e-08 0 2.1838e-08 0 2.1841e-08 0.0007 2.1844e-08 0 2.1899e-08 0 2.1902e-08 0.0007 2.1905e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.2021e-08 0 2.2024e-08 0.0007 2.2027e-08 0 2.2082e-08 0 2.2085e-08 0.0007 2.2088e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2204e-08 0 2.2207e-08 0.0007 2.221e-08 0 2.2265e-08 0 2.2268e-08 0.0007 2.2271e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2448e-08 0 2.2451e-08 0.0007 2.2454e-08 0 2.2509e-08 0 2.2512e-08 0.0007 2.2515e-08 0 2.257e-08 0 2.2573e-08 0.0007 2.2576e-08 0 2.2631e-08 0 2.2634e-08 0.0007 2.2637e-08 0 2.2692e-08 0 2.2695e-08 0.0007 2.2698e-08 0 2.2753e-08 0 2.2756e-08 0.0007 2.2759e-08 0 2.2814e-08 0 2.2817e-08 0.0007 2.282e-08 0 2.2875e-08 0 2.2878e-08 0.0007 2.2881e-08 0 2.2936e-08 0 2.2939e-08 0.0007 2.2942e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3058e-08 0 2.3061e-08 0.0007 2.3064e-08 0 2.3119e-08 0 2.3122e-08 0.0007 2.3125e-08 0 2.318e-08 0 2.3183e-08 0.0007 2.3186e-08 0 2.3241e-08 0 2.3244e-08 0.0007 2.3247e-08 0 2.3302e-08 0 2.3305e-08 0.0007 2.3308e-08 0 2.3363e-08 0 2.3366e-08 0.0007 2.3369e-08 0 2.3424e-08 0 2.3427e-08 0.0007 2.343e-08 0 2.3485e-08 0 2.3488e-08 0.0007 2.3491e-08 0 2.3546e-08 0 2.3549e-08 0.0007 2.3552e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3668e-08 0 2.3671e-08 0.0007 2.3674e-08 0 2.3729e-08 0 2.3732e-08 0.0007 2.3735e-08 0 2.379e-08 0 2.3793e-08 0.0007 2.3796e-08 0 2.3851e-08 0 2.3854e-08 0.0007 2.3857e-08 0 2.3912e-08 0 2.3915e-08 0.0007 2.3918e-08 0 2.3973e-08 0 2.3976e-08 0.0007 2.3979e-08 0 2.4034e-08 0 2.4037e-08 0.0007 2.404e-08 0 2.4095e-08 0 2.4098e-08 0.0007 2.4101e-08 0 2.4156e-08 0 2.4159e-08 0.0007 2.4162e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4278e-08 0 2.4281e-08 0.0007 2.4284e-08 0)
L_S1|A1 G0_2_RX _S1|A1  2.067833848e-12
L_S1|A2 _S1|A1 _S1|A2  4.135667696e-12
L_S1|A3 _S1|A3 _S1|AB  8.271335392e-12
L_S1|B1 IP1_2_OUT_RX _S1|B1  2.067833848e-12
L_S1|B2 _S1|B1 _S1|B2  4.135667696e-12
L_S1|B3 _S1|B3 _S1|AB  8.271335392e-12
L_S1|T1 T13 _S1|T1  2.067833848e-12
L_S1|T2 _S1|T1 _S1|T2  4.135667696e-12
L_S1|Q2 _S1|ABTQ _S1|Q1  4.135667696e-12
L_S1|Q1 _S1|Q1 S1  2.067833848e-12
IT14|T 0 T14  PWL(0 0 5e-14 0 3.05e-12 0.0007 6.05e-12 0 6.105e-11 0 6.405e-11 0.0007 6.705e-11 0 1.2205e-10 0 1.2505e-10 0.0007 1.2805e-10 0 1.8305e-10 0 1.8605e-10 0.0007 1.8905e-10 0 2.4405e-10 0 2.4705e-10 0.0007 2.5005e-10 0 3.0505e-10 0 3.0805e-10 0.0007 3.1105e-10 0 3.6605e-10 0 3.6905e-10 0.0007 3.7205e-10 0 4.2705e-10 0 4.3005e-10 0.0007 4.3305e-10 0 4.8805e-10 0 4.9105e-10 0.0007 4.9405e-10 0 5.4905e-10 0 5.5205e-10 0.0007 5.5505e-10 0 6.1005e-10 0 6.1305e-10 0.0007 6.1605e-10 0 6.7105e-10 0 6.7405e-10 0.0007 6.7705e-10 0 7.3205e-10 0 7.3505e-10 0.0007 7.3805e-10 0 7.9305e-10 0 7.9605e-10 0.0007 7.9905e-10 0 8.5405e-10 0 8.5705e-10 0.0007 8.6005e-10 0 9.1505e-10 0 9.1805e-10 0.0007 9.2105e-10 0 9.7605e-10 0 9.7905e-10 0.0007 9.8205e-10 0 1.03705e-09 0 1.04005e-09 0.0007 1.04305e-09 0 1.09805e-09 0 1.10105e-09 0.0007 1.10405e-09 0 1.15905e-09 0 1.16205e-09 0.0007 1.16505e-09 0 1.22005e-09 0 1.22305e-09 0.0007 1.22605e-09 0 1.28105e-09 0 1.28405e-09 0.0007 1.28705e-09 0 1.34205e-09 0 1.34505e-09 0.0007 1.34805e-09 0 1.40305e-09 0 1.40605e-09 0.0007 1.40905e-09 0 1.46405e-09 0 1.46705e-09 0.0007 1.47005e-09 0 1.52505e-09 0 1.52805e-09 0.0007 1.53105e-09 0 1.58605e-09 0 1.58905e-09 0.0007 1.59205e-09 0 1.64705e-09 0 1.65005e-09 0.0007 1.65305e-09 0 1.70805e-09 0 1.71105e-09 0.0007 1.71405e-09 0 1.76905e-09 0 1.77205e-09 0.0007 1.77505e-09 0 1.83005e-09 0 1.83305e-09 0.0007 1.83605e-09 0 1.89105e-09 0 1.89405e-09 0.0007 1.89705e-09 0 1.95205e-09 0 1.95505e-09 0.0007 1.95805e-09 0 2.01305e-09 0 2.01605e-09 0.0007 2.01905e-09 0 2.07405e-09 0 2.07705e-09 0.0007 2.08005e-09 0 2.13505e-09 0 2.13805e-09 0.0007 2.14105e-09 0 2.19605e-09 0 2.19905e-09 0.0007 2.20205e-09 0 2.25705e-09 0 2.26005e-09 0.0007 2.26305e-09 0 2.31805e-09 0 2.32105e-09 0.0007 2.32405e-09 0 2.37905e-09 0 2.38205e-09 0.0007 2.38505e-09 0 2.44005e-09 0 2.44305e-09 0.0007 2.44605e-09 0 2.50105e-09 0 2.50405e-09 0.0007 2.50705e-09 0 2.56205e-09 0 2.56505e-09 0.0007 2.56805e-09 0 2.62305e-09 0 2.62605e-09 0.0007 2.62905e-09 0 2.68405e-09 0 2.68705e-09 0.0007 2.69005e-09 0 2.74505e-09 0 2.74805e-09 0.0007 2.75105e-09 0 2.80605e-09 0 2.80905e-09 0.0007 2.81205e-09 0 2.86705e-09 0 2.87005e-09 0.0007 2.87305e-09 0 2.92805e-09 0 2.93105e-09 0.0007 2.93405e-09 0 2.98905e-09 0 2.99205e-09 0.0007 2.99505e-09 0 3.05005e-09 0 3.05305e-09 0.0007 3.05605e-09 0 3.11105e-09 0 3.11405e-09 0.0007 3.11705e-09 0 3.17205e-09 0 3.17505e-09 0.0007 3.17805e-09 0 3.23305e-09 0 3.23605e-09 0.0007 3.23905e-09 0 3.29405e-09 0 3.29705e-09 0.0007 3.30005e-09 0 3.35505e-09 0 3.35805e-09 0.0007 3.36105e-09 0 3.41605e-09 0 3.41905e-09 0.0007 3.42205e-09 0 3.47705e-09 0 3.48005e-09 0.0007 3.48305e-09 0 3.53805e-09 0 3.54105e-09 0.0007 3.54405e-09 0 3.59905e-09 0 3.60205e-09 0.0007 3.60505e-09 0 3.66005e-09 0 3.66305e-09 0.0007 3.66605e-09 0 3.72105e-09 0 3.72405e-09 0.0007 3.72705e-09 0 3.78205e-09 0 3.78505e-09 0.0007 3.78805e-09 0 3.84305e-09 0 3.84605e-09 0.0007 3.84905e-09 0 3.90405e-09 0 3.90705e-09 0.0007 3.91005e-09 0 3.96505e-09 0 3.96805e-09 0.0007 3.97105e-09 0 4.02605e-09 0 4.02905e-09 0.0007 4.03205e-09 0 4.08705e-09 0 4.09005e-09 0.0007 4.09305e-09 0 4.14805e-09 0 4.15105e-09 0.0007 4.15405e-09 0 4.20905e-09 0 4.21205e-09 0.0007 4.21505e-09 0 4.27005e-09 0 4.27305e-09 0.0007 4.27605e-09 0 4.33105e-09 0 4.33405e-09 0.0007 4.33705e-09 0 4.39205e-09 0 4.39505e-09 0.0007 4.39805e-09 0 4.45305e-09 0 4.45605e-09 0.0007 4.45905e-09 0 4.51405e-09 0 4.51705e-09 0.0007 4.52005e-09 0 4.57505e-09 0 4.57805e-09 0.0007 4.58105e-09 0 4.63605e-09 0 4.63905e-09 0.0007 4.64205e-09 0 4.69705e-09 0 4.70005e-09 0.0007 4.70305e-09 0 4.75805e-09 0 4.76105e-09 0.0007 4.76405e-09 0 4.81905e-09 0 4.82205e-09 0.0007 4.82505e-09 0 4.88005e-09 0 4.88305e-09 0.0007 4.88605e-09 0 4.94105e-09 0 4.94405e-09 0.0007 4.94705e-09 0 5.00205e-09 0 5.00505e-09 0.0007 5.00805e-09 0 5.06305e-09 0 5.06605e-09 0.0007 5.06905e-09 0 5.12405e-09 0 5.12705e-09 0.0007 5.13005e-09 0 5.18505e-09 0 5.18805e-09 0.0007 5.19105e-09 0 5.24605e-09 0 5.24905e-09 0.0007 5.25205e-09 0 5.30705e-09 0 5.31005e-09 0.0007 5.31305e-09 0 5.36805e-09 0 5.37105e-09 0.0007 5.37405e-09 0 5.42905e-09 0 5.43205e-09 0.0007 5.43505e-09 0 5.49005e-09 0 5.49305e-09 0.0007 5.49605e-09 0 5.55105e-09 0 5.55405e-09 0.0007 5.55705e-09 0 5.61205e-09 0 5.61505e-09 0.0007 5.61805e-09 0 5.67305e-09 0 5.67605e-09 0.0007 5.67905e-09 0 5.73405e-09 0 5.73705e-09 0.0007 5.74005e-09 0 5.79505e-09 0 5.79805e-09 0.0007 5.80105e-09 0 5.85605e-09 0 5.85905e-09 0.0007 5.86205e-09 0 5.91705e-09 0 5.92005e-09 0.0007 5.92305e-09 0 5.97805e-09 0 5.98105e-09 0.0007 5.98405e-09 0 6.03905e-09 0 6.04205e-09 0.0007 6.04505e-09 0 6.10005e-09 0 6.10305e-09 0.0007 6.10605e-09 0 6.16105e-09 0 6.16405e-09 0.0007 6.16705e-09 0 6.22205e-09 0 6.22505e-09 0.0007 6.22805e-09 0 6.28305e-09 0 6.28605e-09 0.0007 6.28905e-09 0 6.34405e-09 0 6.34705e-09 0.0007 6.35005e-09 0 6.40505e-09 0 6.40805e-09 0.0007 6.41105e-09 0 6.46605e-09 0 6.46905e-09 0.0007 6.47205e-09 0 6.52705e-09 0 6.53005e-09 0.0007 6.53305e-09 0 6.58805e-09 0 6.59105e-09 0.0007 6.59405e-09 0 6.64905e-09 0 6.65205e-09 0.0007 6.65505e-09 0 6.71005e-09 0 6.71305e-09 0.0007 6.71605e-09 0 6.77105e-09 0 6.77405e-09 0.0007 6.77705e-09 0 6.83205e-09 0 6.83505e-09 0.0007 6.83805e-09 0 6.89305e-09 0 6.89605e-09 0.0007 6.89905e-09 0 6.95405e-09 0 6.95705e-09 0.0007 6.96005e-09 0 7.01505e-09 0 7.01805e-09 0.0007 7.02105e-09 0 7.07605e-09 0 7.07905e-09 0.0007 7.08205e-09 0 7.13705e-09 0 7.14005e-09 0.0007 7.14305e-09 0 7.19805e-09 0 7.20105e-09 0.0007 7.20405e-09 0 7.25905e-09 0 7.26205e-09 0.0007 7.26505e-09 0 7.32005e-09 0 7.32305e-09 0.0007 7.32605e-09 0 7.38105e-09 0 7.38405e-09 0.0007 7.38705e-09 0 7.44205e-09 0 7.44505e-09 0.0007 7.44805e-09 0 7.50305e-09 0 7.50605e-09 0.0007 7.50905e-09 0 7.56405e-09 0 7.56705e-09 0.0007 7.57005e-09 0 7.62505e-09 0 7.62805e-09 0.0007 7.63105e-09 0 7.68605e-09 0 7.68905e-09 0.0007 7.69205e-09 0 7.74705e-09 0 7.75005e-09 0.0007 7.75305e-09 0 7.80805e-09 0 7.81105e-09 0.0007 7.81405e-09 0 7.86905e-09 0 7.87205e-09 0.0007 7.87505e-09 0 7.93005e-09 0 7.93305e-09 0.0007 7.93605e-09 0 7.99105e-09 0 7.99405e-09 0.0007 7.99705e-09 0 8.05205e-09 0 8.05505e-09 0.0007 8.05805e-09 0 8.11305e-09 0 8.11605e-09 0.0007 8.11905e-09 0 8.17405e-09 0 8.17705e-09 0.0007 8.18005e-09 0 8.23505e-09 0 8.23805e-09 0.0007 8.24105e-09 0 8.29605e-09 0 8.29905e-09 0.0007 8.30205e-09 0 8.35705e-09 0 8.36005e-09 0.0007 8.36305e-09 0 8.41805e-09 0 8.42105e-09 0.0007 8.42405e-09 0 8.47905e-09 0 8.48205e-09 0.0007 8.48505e-09 0 8.54005e-09 0 8.54305e-09 0.0007 8.54605e-09 0 8.60105e-09 0 8.60405e-09 0.0007 8.60705e-09 0 8.66205e-09 0 8.66505e-09 0.0007 8.66805e-09 0 8.72305e-09 0 8.72605e-09 0.0007 8.72905e-09 0 8.78405e-09 0 8.78705e-09 0.0007 8.79005e-09 0 8.84505e-09 0 8.84805e-09 0.0007 8.85105e-09 0 8.90605e-09 0 8.90905e-09 0.0007 8.91205e-09 0 8.96705e-09 0 8.97005e-09 0.0007 8.97305e-09 0 9.02805e-09 0 9.03105e-09 0.0007 9.03405e-09 0 9.08905e-09 0 9.09205e-09 0.0007 9.09505e-09 0 9.15005e-09 0 9.15305e-09 0.0007 9.15605e-09 0 9.21105e-09 0 9.21405e-09 0.0007 9.21705e-09 0 9.27205e-09 0 9.27505e-09 0.0007 9.27805e-09 0 9.33305e-09 0 9.33605e-09 0.0007 9.33905e-09 0 9.39405e-09 0 9.39705e-09 0.0007 9.40005e-09 0 9.45505e-09 0 9.45805e-09 0.0007 9.46105e-09 0 9.51605e-09 0 9.51905e-09 0.0007 9.52205e-09 0 9.57705e-09 0 9.58005e-09 0.0007 9.58305e-09 0 9.63805e-09 0 9.64105e-09 0.0007 9.64405e-09 0 9.69905e-09 0 9.70205e-09 0.0007 9.70505e-09 0 9.76005e-09 0 9.76305e-09 0.0007 9.76605e-09 0 9.82105e-09 0 9.82405e-09 0.0007 9.82705e-09 0 9.88205e-09 0 9.88505e-09 0.0007 9.88805e-09 0 9.94305e-09 0 9.94605e-09 0.0007 9.94905e-09 0 1.0004e-08 0 1.0007e-08 0.0007 1.001e-08 0 1.0065e-08 0 1.0068e-08 0.0007 1.0071e-08 0 1.0126e-08 0 1.0129e-08 0.0007 1.0132e-08 0 1.0187e-08 0 1.019e-08 0.0007 1.01931e-08 0 1.0248e-08 0 1.0251e-08 0.0007 1.0254e-08 0 1.0309e-08 0 1.0312e-08 0.0007 1.0315e-08 0 1.037e-08 0 1.0373e-08 0.0007 1.0376e-08 0 1.0431e-08 0 1.0434e-08 0.0007 1.0437e-08 0 1.0492e-08 0 1.0495e-08 0.0007 1.0498e-08 0 1.0553e-08 0 1.0556e-08 0.0007 1.0559e-08 0 1.0614e-08 0 1.0617e-08 0.0007 1.062e-08 0 1.0675e-08 0 1.0678e-08 0.0007 1.0681e-08 0 1.0736e-08 0 1.0739e-08 0.0007 1.0742e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0858e-08 0 1.0861e-08 0.0007 1.0864e-08 0 1.0919e-08 0 1.0922e-08 0.0007 1.0925e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.1041e-08 0 1.1044e-08 0.0007 1.1047e-08 0 1.1102e-08 0 1.1105e-08 0.0007 1.1108e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1224e-08 0 1.1227e-08 0.0007 1.123e-08 0 1.1285e-08 0 1.1288e-08 0.0007 1.1291e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1468e-08 0 1.1471e-08 0.0007 1.1474e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.159e-08 0 1.1593e-08 0.0007 1.1596e-08 0 1.1651e-08 0 1.1654e-08 0.0007 1.1657e-08 0 1.1712e-08 0 1.1715e-08 0.0007 1.1718e-08 0 1.1773e-08 0 1.1776e-08 0.0007 1.1779e-08 0 1.1834e-08 0 1.1837e-08 0.0007 1.184e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.1956e-08 0 1.1959e-08 0.0007 1.1962e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2078e-08 0 1.2081e-08 0.0007 1.2084e-08 0 1.2139e-08 0 1.2142e-08 0.0007 1.2145e-08 0 1.22e-08 0 1.2203e-08 0.0007 1.2206e-08 0 1.2261e-08 0 1.2264e-08 0.0007 1.2267e-08 0 1.2322e-08 0 1.2325e-08 0.0007 1.2328e-08 0 1.2383e-08 0 1.2386e-08 0.0007 1.2389e-08 0 1.2444e-08 0 1.2447e-08 0.0007 1.245e-08 0 1.2505e-08 0 1.2508e-08 0.0007 1.2511e-08 0 1.2566e-08 0 1.2569e-08 0.0007 1.2572e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2688e-08 0 1.2691e-08 0.0007 1.2694e-08 0 1.2749e-08 0 1.2752e-08 0.0007 1.2755e-08 0 1.281e-08 0 1.2813e-08 0.0007 1.2816e-08 0 1.2871e-08 0 1.2874e-08 0.0007 1.2877e-08 0 1.2932e-08 0 1.2935e-08 0.0007 1.2938e-08 0 1.2993e-08 0 1.2996e-08 0.0007 1.2999e-08 0 1.3054e-08 0 1.3057e-08 0.0007 1.306e-08 0 1.3115e-08 0 1.3118e-08 0.0007 1.3121e-08 0 1.3176e-08 0 1.3179e-08 0.0007 1.3182e-08 0 1.3237e-08 0 1.324e-08 0.0007 1.3243e-08 0 1.3298e-08 0 1.3301e-08 0.0007 1.3304e-08 0 1.3359e-08 0 1.3362e-08 0.0007 1.3365e-08 0 1.342e-08 0 1.3423e-08 0.0007 1.3426e-08 0 1.3481e-08 0 1.3484e-08 0.0007 1.3487e-08 0 1.3542e-08 0 1.3545e-08 0.0007 1.3548e-08 0 1.3603e-08 0 1.3606e-08 0.0007 1.3609e-08 0 1.3664e-08 0 1.3667e-08 0.0007 1.367e-08 0 1.3725e-08 0 1.3728e-08 0.0007 1.3731e-08 0 1.3786e-08 0 1.3789e-08 0.0007 1.3792e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.3908e-08 0 1.3911e-08 0.0007 1.3914e-08 0 1.3969e-08 0 1.3972e-08 0.0007 1.3975e-08 0 1.403e-08 0 1.4033e-08 0.0007 1.4036e-08 0 1.4091e-08 0 1.4094e-08 0.0007 1.4097e-08 0 1.4152e-08 0 1.4155e-08 0.0007 1.4158e-08 0 1.4213e-08 0 1.4216e-08 0.0007 1.4219e-08 0 1.4274e-08 0 1.4277e-08 0.0007 1.428e-08 0 1.4335e-08 0 1.4338e-08 0.0007 1.4341e-08 0 1.4396e-08 0 1.4399e-08 0.0007 1.4402e-08 0 1.4457e-08 0 1.446e-08 0.0007 1.4463e-08 0 1.4518e-08 0 1.4521e-08 0.0007 1.4524e-08 0 1.4579e-08 0 1.4582e-08 0.0007 1.4585e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.4701e-08 0 1.4704e-08 0.0007 1.4707e-08 0 1.4762e-08 0 1.4765e-08 0.0007 1.4768e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4884e-08 0 1.4887e-08 0.0007 1.489e-08 0 1.4945e-08 0 1.4948e-08 0.0007 1.4951e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5067e-08 0 1.507e-08 0.0007 1.5073e-08 0 1.5128e-08 0 1.5131e-08 0.0007 1.5134e-08 0 1.5189e-08 0 1.5192e-08 0.0007 1.5195e-08 0 1.52501e-08 0 1.52531e-08 0.0007 1.52561e-08 0 1.5311e-08 0 1.53141e-08 0.0007 1.53171e-08 0 1.5372e-08 0 1.5375e-08 0.0007 1.5378e-08 0 1.5433e-08 0 1.5436e-08 0.0007 1.5439e-08 0 1.5494e-08 0 1.5497e-08 0.0007 1.55e-08 0 1.5555e-08 0 1.5558e-08 0.0007 1.5561e-08 0 1.5616e-08 0 1.5619e-08 0.0007 1.5622e-08 0 1.5677e-08 0 1.568e-08 0.0007 1.5683e-08 0 1.5738e-08 0 1.5741e-08 0.0007 1.5744e-08 0 1.5799e-08 0 1.5802e-08 0.0007 1.5805e-08 0 1.586e-08 0 1.5863e-08 0.0007 1.5866e-08 0 1.59211e-08 0 1.59241e-08 0.0007 1.59271e-08 0 1.5982e-08 0 1.5985e-08 0.0007 1.59881e-08 0 1.6043e-08 0 1.6046e-08 0.0007 1.6049e-08 0 1.6104e-08 0 1.6107e-08 0.0007 1.611e-08 0 1.6165e-08 0 1.6168e-08 0.0007 1.6171e-08 0 1.6226e-08 0 1.6229e-08 0.0007 1.6232e-08 0 1.6287e-08 0 1.629e-08 0.0007 1.6293e-08 0 1.6348e-08 0 1.6351e-08 0.0007 1.6354e-08 0 1.6409e-08 0 1.6412e-08 0.0007 1.6415e-08 0 1.647e-08 0 1.6473e-08 0.0007 1.6476e-08 0 1.65311e-08 0 1.65341e-08 0.0007 1.65371e-08 0 1.65921e-08 0 1.65951e-08 0.0007 1.65981e-08 0 1.6653e-08 0 1.6656e-08 0.0007 1.6659e-08 0 1.6714e-08 0 1.6717e-08 0.0007 1.672e-08 0 1.6775e-08 0 1.6778e-08 0.0007 1.6781e-08 0 1.6836e-08 0 1.6839e-08 0.0007 1.6842e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6958e-08 0 1.6961e-08 0.0007 1.6964e-08 0 1.7019e-08 0 1.7022e-08 0.0007 1.7025e-08 0 1.708e-08 0 1.7083e-08 0.0007 1.7086e-08 0 1.7141e-08 0 1.7144e-08 0.0007 1.7147e-08 0 1.72021e-08 0 1.72051e-08 0.0007 1.72081e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.72691e-08 0 1.7324e-08 0 1.7327e-08 0.0007 1.733e-08 0 1.7385e-08 0 1.7388e-08 0.0007 1.7391e-08 0 1.7446e-08 0 1.7449e-08 0.0007 1.7452e-08 0 1.7507e-08 0 1.751e-08 0.0007 1.7513e-08 0 1.7568e-08 0 1.7571e-08 0.0007 1.7574e-08 0 1.7629e-08 0 1.7632e-08 0.0007 1.7635e-08 0 1.769e-08 0 1.7693e-08 0.0007 1.7696e-08 0 1.7751e-08 0 1.7754e-08 0.0007 1.7757e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.78731e-08 0 1.78761e-08 0.0007 1.78791e-08 0 1.7934e-08 0 1.7937e-08 0.0007 1.794e-08 0 1.7995e-08 0 1.7998e-08 0.0007 1.8001e-08 0 1.8056e-08 0 1.8059e-08 0.0007 1.8062e-08 0 1.8117e-08 0 1.812e-08 0.0007 1.8123e-08 0 1.8178e-08 0 1.8181e-08 0.0007 1.8184e-08 0 1.8239e-08 0 1.8242e-08 0.0007 1.8245e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.8361e-08 0 1.8364e-08 0.0007 1.8367e-08 0 1.8422e-08 0 1.8425e-08 0.0007 1.8428e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8544e-08 0 1.8547e-08 0.0007 1.85501e-08 0 1.8605e-08 0 1.8608e-08 0.0007 1.8611e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8727e-08 0 1.873e-08 0.0007 1.8733e-08 0 1.8788e-08 0 1.8791e-08 0.0007 1.8794e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.891e-08 0 1.8913e-08 0.0007 1.8916e-08 0 1.8971e-08 0 1.8974e-08 0.0007 1.8977e-08 0 1.9032e-08 0 1.9035e-08 0.0007 1.9038e-08 0 1.9093e-08 0 1.9096e-08 0.0007 1.9099e-08 0 1.91541e-08 0 1.91571e-08 0.0007 1.91601e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9276e-08 0 1.9279e-08 0.0007 1.9282e-08 0 1.9337e-08 0 1.934e-08 0.0007 1.9343e-08 0 1.9398e-08 0 1.9401e-08 0.0007 1.9404e-08 0 1.9459e-08 0 1.9462e-08 0.0007 1.9465e-08 0 1.952e-08 0 1.9523e-08 0.0007 1.9526e-08 0 1.9581e-08 0 1.9584e-08 0.0007 1.9587e-08 0 1.9642e-08 0 1.9645e-08 0.0007 1.9648e-08 0 1.9703e-08 0 1.9706e-08 0.0007 1.9709e-08 0 1.9764e-08 0 1.9767e-08 0.0007 1.977e-08 0 1.9825e-08 0 1.9828e-08 0.0007 1.98311e-08 0 1.9886e-08 0 1.9889e-08 0.0007 1.9892e-08 0 1.9947e-08 0 1.995e-08 0.0007 1.9953e-08 0 2.0008e-08 0 2.0011e-08 0.0007 2.0014e-08 0 2.0069e-08 0 2.0072e-08 0.0007 2.0075e-08 0 2.013e-08 0 2.0133e-08 0.0007 2.0136e-08 0 2.0191e-08 0 2.0194e-08 0.0007 2.0197e-08 0 2.0252e-08 0 2.0255e-08 0.0007 2.0258e-08 0 2.0313e-08 0 2.0316e-08 0.0007 2.0319e-08 0 2.0374e-08 0 2.0377e-08 0.0007 2.038e-08 0 2.04351e-08 0 2.04381e-08 0.0007 2.04411e-08 0 2.0496e-08 0 2.0499e-08 0.0007 2.0502e-08 0 2.0557e-08 0 2.056e-08 0.0007 2.0563e-08 0 2.0618e-08 0 2.0621e-08 0.0007 2.0624e-08 0 2.0679e-08 0 2.0682e-08 0.0007 2.0685e-08 0 2.074e-08 0 2.0743e-08 0.0007 2.0746e-08 0 2.0801e-08 0 2.0804e-08 0.0007 2.0807e-08 0 2.0862e-08 0 2.0865e-08 0.0007 2.0868e-08 0 2.0923e-08 0 2.0926e-08 0.0007 2.0929e-08 0 2.0984e-08 0 2.0987e-08 0.0007 2.099e-08 0 2.1045e-08 0 2.1048e-08 0.0007 2.1051e-08 0 2.1106e-08 0 2.11091e-08 0.0007 2.11121e-08 0 2.1167e-08 0 2.117e-08 0.0007 2.1173e-08 0 2.1228e-08 0 2.1231e-08 0.0007 2.1234e-08 0 2.1289e-08 0 2.1292e-08 0.0007 2.1295e-08 0 2.135e-08 0 2.1353e-08 0.0007 2.1356e-08 0 2.1411e-08 0 2.1414e-08 0.0007 2.1417e-08 0 2.1472e-08 0 2.1475e-08 0.0007 2.1478e-08 0 2.1533e-08 0 2.1536e-08 0.0007 2.1539e-08 0 2.1594e-08 0 2.1597e-08 0.0007 2.16e-08 0 2.1655e-08 0 2.1658e-08 0.0007 2.1661e-08 0 2.1716e-08 0 2.1719e-08 0.0007 2.1722e-08 0 2.1777e-08 0 2.178e-08 0.0007 2.1783e-08 0 2.1838e-08 0 2.1841e-08 0.0007 2.1844e-08 0 2.1899e-08 0 2.1902e-08 0.0007 2.1905e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.2021e-08 0 2.2024e-08 0.0007 2.2027e-08 0 2.2082e-08 0 2.2085e-08 0.0007 2.2088e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2204e-08 0 2.2207e-08 0.0007 2.221e-08 0 2.2265e-08 0 2.2268e-08 0.0007 2.2271e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2448e-08 0 2.2451e-08 0.0007 2.2454e-08 0 2.2509e-08 0 2.2512e-08 0.0007 2.2515e-08 0 2.257e-08 0 2.2573e-08 0.0007 2.2576e-08 0 2.2631e-08 0 2.2634e-08 0.0007 2.2637e-08 0 2.2692e-08 0 2.2695e-08 0.0007 2.2698e-08 0 2.2753e-08 0 2.2756e-08 0.0007 2.2759e-08 0 2.2814e-08 0 2.2817e-08 0.0007 2.282e-08 0 2.2875e-08 0 2.2878e-08 0.0007 2.2881e-08 0 2.2936e-08 0 2.2939e-08 0.0007 2.2942e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3058e-08 0 2.3061e-08 0.0007 2.3064e-08 0 2.3119e-08 0 2.3122e-08 0.0007 2.3125e-08 0 2.318e-08 0 2.3183e-08 0.0007 2.3186e-08 0 2.3241e-08 0 2.3244e-08 0.0007 2.3247e-08 0 2.3302e-08 0 2.3305e-08 0.0007 2.3308e-08 0 2.3363e-08 0 2.3366e-08 0.0007 2.3369e-08 0 2.3424e-08 0 2.3427e-08 0.0007 2.343e-08 0 2.3485e-08 0 2.3488e-08 0.0007 2.3491e-08 0 2.3546e-08 0 2.3549e-08 0.0007 2.3552e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3668e-08 0 2.3671e-08 0.0007 2.3674e-08 0 2.3729e-08 0 2.3732e-08 0.0007 2.3735e-08 0 2.379e-08 0 2.3793e-08 0.0007 2.3796e-08 0 2.3851e-08 0 2.3854e-08 0.0007 2.3857e-08 0 2.3912e-08 0 2.3915e-08 0.0007 2.3918e-08 0 2.3973e-08 0 2.3976e-08 0.0007 2.3979e-08 0 2.4034e-08 0 2.4037e-08 0.0007 2.404e-08 0 2.4095e-08 0 2.4098e-08 0.0007 2.4101e-08 0 2.4156e-08 0 2.4159e-08 0.0007 2.4162e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4278e-08 0 2.4281e-08 0.0007 2.4284e-08 0)
L_S2|A1 G1_2_RX _S2|A1  2.067833848e-12
L_S2|A2 _S2|A1 _S2|A2  4.135667696e-12
L_S2|A3 _S2|A3 _S2|AB  8.271335392e-12
L_S2|B1 IP2_2_OUT_RX _S2|B1  2.067833848e-12
L_S2|B2 _S2|B1 _S2|B2  4.135667696e-12
L_S2|B3 _S2|B3 _S2|AB  8.271335392e-12
L_S2|T1 T14 _S2|T1  2.067833848e-12
L_S2|T2 _S2|T1 _S2|T2  4.135667696e-12
L_S2|Q2 _S2|ABTQ _S2|Q1  4.135667696e-12
L_S2|Q1 _S2|Q1 S2  2.067833848e-12
IT15|T 0 T15  PWL(0 0 5e-14 0 3.05e-12 0.0007 6.05e-12 0 6.105e-11 0 6.405e-11 0.0007 6.705e-11 0 1.2205e-10 0 1.2505e-10 0.0007 1.2805e-10 0 1.8305e-10 0 1.8605e-10 0.0007 1.8905e-10 0 2.4405e-10 0 2.4705e-10 0.0007 2.5005e-10 0 3.0505e-10 0 3.0805e-10 0.0007 3.1105e-10 0 3.6605e-10 0 3.6905e-10 0.0007 3.7205e-10 0 4.2705e-10 0 4.3005e-10 0.0007 4.3305e-10 0 4.8805e-10 0 4.9105e-10 0.0007 4.9405e-10 0 5.4905e-10 0 5.5205e-10 0.0007 5.5505e-10 0 6.1005e-10 0 6.1305e-10 0.0007 6.1605e-10 0 6.7105e-10 0 6.7405e-10 0.0007 6.7705e-10 0 7.3205e-10 0 7.3505e-10 0.0007 7.3805e-10 0 7.9305e-10 0 7.9605e-10 0.0007 7.9905e-10 0 8.5405e-10 0 8.5705e-10 0.0007 8.6005e-10 0 9.1505e-10 0 9.1805e-10 0.0007 9.2105e-10 0 9.7605e-10 0 9.7905e-10 0.0007 9.8205e-10 0 1.03705e-09 0 1.04005e-09 0.0007 1.04305e-09 0 1.09805e-09 0 1.10105e-09 0.0007 1.10405e-09 0 1.15905e-09 0 1.16205e-09 0.0007 1.16505e-09 0 1.22005e-09 0 1.22305e-09 0.0007 1.22605e-09 0 1.28105e-09 0 1.28405e-09 0.0007 1.28705e-09 0 1.34205e-09 0 1.34505e-09 0.0007 1.34805e-09 0 1.40305e-09 0 1.40605e-09 0.0007 1.40905e-09 0 1.46405e-09 0 1.46705e-09 0.0007 1.47005e-09 0 1.52505e-09 0 1.52805e-09 0.0007 1.53105e-09 0 1.58605e-09 0 1.58905e-09 0.0007 1.59205e-09 0 1.64705e-09 0 1.65005e-09 0.0007 1.65305e-09 0 1.70805e-09 0 1.71105e-09 0.0007 1.71405e-09 0 1.76905e-09 0 1.77205e-09 0.0007 1.77505e-09 0 1.83005e-09 0 1.83305e-09 0.0007 1.83605e-09 0 1.89105e-09 0 1.89405e-09 0.0007 1.89705e-09 0 1.95205e-09 0 1.95505e-09 0.0007 1.95805e-09 0 2.01305e-09 0 2.01605e-09 0.0007 2.01905e-09 0 2.07405e-09 0 2.07705e-09 0.0007 2.08005e-09 0 2.13505e-09 0 2.13805e-09 0.0007 2.14105e-09 0 2.19605e-09 0 2.19905e-09 0.0007 2.20205e-09 0 2.25705e-09 0 2.26005e-09 0.0007 2.26305e-09 0 2.31805e-09 0 2.32105e-09 0.0007 2.32405e-09 0 2.37905e-09 0 2.38205e-09 0.0007 2.38505e-09 0 2.44005e-09 0 2.44305e-09 0.0007 2.44605e-09 0 2.50105e-09 0 2.50405e-09 0.0007 2.50705e-09 0 2.56205e-09 0 2.56505e-09 0.0007 2.56805e-09 0 2.62305e-09 0 2.62605e-09 0.0007 2.62905e-09 0 2.68405e-09 0 2.68705e-09 0.0007 2.69005e-09 0 2.74505e-09 0 2.74805e-09 0.0007 2.75105e-09 0 2.80605e-09 0 2.80905e-09 0.0007 2.81205e-09 0 2.86705e-09 0 2.87005e-09 0.0007 2.87305e-09 0 2.92805e-09 0 2.93105e-09 0.0007 2.93405e-09 0 2.98905e-09 0 2.99205e-09 0.0007 2.99505e-09 0 3.05005e-09 0 3.05305e-09 0.0007 3.05605e-09 0 3.11105e-09 0 3.11405e-09 0.0007 3.11705e-09 0 3.17205e-09 0 3.17505e-09 0.0007 3.17805e-09 0 3.23305e-09 0 3.23605e-09 0.0007 3.23905e-09 0 3.29405e-09 0 3.29705e-09 0.0007 3.30005e-09 0 3.35505e-09 0 3.35805e-09 0.0007 3.36105e-09 0 3.41605e-09 0 3.41905e-09 0.0007 3.42205e-09 0 3.47705e-09 0 3.48005e-09 0.0007 3.48305e-09 0 3.53805e-09 0 3.54105e-09 0.0007 3.54405e-09 0 3.59905e-09 0 3.60205e-09 0.0007 3.60505e-09 0 3.66005e-09 0 3.66305e-09 0.0007 3.66605e-09 0 3.72105e-09 0 3.72405e-09 0.0007 3.72705e-09 0 3.78205e-09 0 3.78505e-09 0.0007 3.78805e-09 0 3.84305e-09 0 3.84605e-09 0.0007 3.84905e-09 0 3.90405e-09 0 3.90705e-09 0.0007 3.91005e-09 0 3.96505e-09 0 3.96805e-09 0.0007 3.97105e-09 0 4.02605e-09 0 4.02905e-09 0.0007 4.03205e-09 0 4.08705e-09 0 4.09005e-09 0.0007 4.09305e-09 0 4.14805e-09 0 4.15105e-09 0.0007 4.15405e-09 0 4.20905e-09 0 4.21205e-09 0.0007 4.21505e-09 0 4.27005e-09 0 4.27305e-09 0.0007 4.27605e-09 0 4.33105e-09 0 4.33405e-09 0.0007 4.33705e-09 0 4.39205e-09 0 4.39505e-09 0.0007 4.39805e-09 0 4.45305e-09 0 4.45605e-09 0.0007 4.45905e-09 0 4.51405e-09 0 4.51705e-09 0.0007 4.52005e-09 0 4.57505e-09 0 4.57805e-09 0.0007 4.58105e-09 0 4.63605e-09 0 4.63905e-09 0.0007 4.64205e-09 0 4.69705e-09 0 4.70005e-09 0.0007 4.70305e-09 0 4.75805e-09 0 4.76105e-09 0.0007 4.76405e-09 0 4.81905e-09 0 4.82205e-09 0.0007 4.82505e-09 0 4.88005e-09 0 4.88305e-09 0.0007 4.88605e-09 0 4.94105e-09 0 4.94405e-09 0.0007 4.94705e-09 0 5.00205e-09 0 5.00505e-09 0.0007 5.00805e-09 0 5.06305e-09 0 5.06605e-09 0.0007 5.06905e-09 0 5.12405e-09 0 5.12705e-09 0.0007 5.13005e-09 0 5.18505e-09 0 5.18805e-09 0.0007 5.19105e-09 0 5.24605e-09 0 5.24905e-09 0.0007 5.25205e-09 0 5.30705e-09 0 5.31005e-09 0.0007 5.31305e-09 0 5.36805e-09 0 5.37105e-09 0.0007 5.37405e-09 0 5.42905e-09 0 5.43205e-09 0.0007 5.43505e-09 0 5.49005e-09 0 5.49305e-09 0.0007 5.49605e-09 0 5.55105e-09 0 5.55405e-09 0.0007 5.55705e-09 0 5.61205e-09 0 5.61505e-09 0.0007 5.61805e-09 0 5.67305e-09 0 5.67605e-09 0.0007 5.67905e-09 0 5.73405e-09 0 5.73705e-09 0.0007 5.74005e-09 0 5.79505e-09 0 5.79805e-09 0.0007 5.80105e-09 0 5.85605e-09 0 5.85905e-09 0.0007 5.86205e-09 0 5.91705e-09 0 5.92005e-09 0.0007 5.92305e-09 0 5.97805e-09 0 5.98105e-09 0.0007 5.98405e-09 0 6.03905e-09 0 6.04205e-09 0.0007 6.04505e-09 0 6.10005e-09 0 6.10305e-09 0.0007 6.10605e-09 0 6.16105e-09 0 6.16405e-09 0.0007 6.16705e-09 0 6.22205e-09 0 6.22505e-09 0.0007 6.22805e-09 0 6.28305e-09 0 6.28605e-09 0.0007 6.28905e-09 0 6.34405e-09 0 6.34705e-09 0.0007 6.35005e-09 0 6.40505e-09 0 6.40805e-09 0.0007 6.41105e-09 0 6.46605e-09 0 6.46905e-09 0.0007 6.47205e-09 0 6.52705e-09 0 6.53005e-09 0.0007 6.53305e-09 0 6.58805e-09 0 6.59105e-09 0.0007 6.59405e-09 0 6.64905e-09 0 6.65205e-09 0.0007 6.65505e-09 0 6.71005e-09 0 6.71305e-09 0.0007 6.71605e-09 0 6.77105e-09 0 6.77405e-09 0.0007 6.77705e-09 0 6.83205e-09 0 6.83505e-09 0.0007 6.83805e-09 0 6.89305e-09 0 6.89605e-09 0.0007 6.89905e-09 0 6.95405e-09 0 6.95705e-09 0.0007 6.96005e-09 0 7.01505e-09 0 7.01805e-09 0.0007 7.02105e-09 0 7.07605e-09 0 7.07905e-09 0.0007 7.08205e-09 0 7.13705e-09 0 7.14005e-09 0.0007 7.14305e-09 0 7.19805e-09 0 7.20105e-09 0.0007 7.20405e-09 0 7.25905e-09 0 7.26205e-09 0.0007 7.26505e-09 0 7.32005e-09 0 7.32305e-09 0.0007 7.32605e-09 0 7.38105e-09 0 7.38405e-09 0.0007 7.38705e-09 0 7.44205e-09 0 7.44505e-09 0.0007 7.44805e-09 0 7.50305e-09 0 7.50605e-09 0.0007 7.50905e-09 0 7.56405e-09 0 7.56705e-09 0.0007 7.57005e-09 0 7.62505e-09 0 7.62805e-09 0.0007 7.63105e-09 0 7.68605e-09 0 7.68905e-09 0.0007 7.69205e-09 0 7.74705e-09 0 7.75005e-09 0.0007 7.75305e-09 0 7.80805e-09 0 7.81105e-09 0.0007 7.81405e-09 0 7.86905e-09 0 7.87205e-09 0.0007 7.87505e-09 0 7.93005e-09 0 7.93305e-09 0.0007 7.93605e-09 0 7.99105e-09 0 7.99405e-09 0.0007 7.99705e-09 0 8.05205e-09 0 8.05505e-09 0.0007 8.05805e-09 0 8.11305e-09 0 8.11605e-09 0.0007 8.11905e-09 0 8.17405e-09 0 8.17705e-09 0.0007 8.18005e-09 0 8.23505e-09 0 8.23805e-09 0.0007 8.24105e-09 0 8.29605e-09 0 8.29905e-09 0.0007 8.30205e-09 0 8.35705e-09 0 8.36005e-09 0.0007 8.36305e-09 0 8.41805e-09 0 8.42105e-09 0.0007 8.42405e-09 0 8.47905e-09 0 8.48205e-09 0.0007 8.48505e-09 0 8.54005e-09 0 8.54305e-09 0.0007 8.54605e-09 0 8.60105e-09 0 8.60405e-09 0.0007 8.60705e-09 0 8.66205e-09 0 8.66505e-09 0.0007 8.66805e-09 0 8.72305e-09 0 8.72605e-09 0.0007 8.72905e-09 0 8.78405e-09 0 8.78705e-09 0.0007 8.79005e-09 0 8.84505e-09 0 8.84805e-09 0.0007 8.85105e-09 0 8.90605e-09 0 8.90905e-09 0.0007 8.91205e-09 0 8.96705e-09 0 8.97005e-09 0.0007 8.97305e-09 0 9.02805e-09 0 9.03105e-09 0.0007 9.03405e-09 0 9.08905e-09 0 9.09205e-09 0.0007 9.09505e-09 0 9.15005e-09 0 9.15305e-09 0.0007 9.15605e-09 0 9.21105e-09 0 9.21405e-09 0.0007 9.21705e-09 0 9.27205e-09 0 9.27505e-09 0.0007 9.27805e-09 0 9.33305e-09 0 9.33605e-09 0.0007 9.33905e-09 0 9.39405e-09 0 9.39705e-09 0.0007 9.40005e-09 0 9.45505e-09 0 9.45805e-09 0.0007 9.46105e-09 0 9.51605e-09 0 9.51905e-09 0.0007 9.52205e-09 0 9.57705e-09 0 9.58005e-09 0.0007 9.58305e-09 0 9.63805e-09 0 9.64105e-09 0.0007 9.64405e-09 0 9.69905e-09 0 9.70205e-09 0.0007 9.70505e-09 0 9.76005e-09 0 9.76305e-09 0.0007 9.76605e-09 0 9.82105e-09 0 9.82405e-09 0.0007 9.82705e-09 0 9.88205e-09 0 9.88505e-09 0.0007 9.88805e-09 0 9.94305e-09 0 9.94605e-09 0.0007 9.94905e-09 0 1.0004e-08 0 1.0007e-08 0.0007 1.001e-08 0 1.0065e-08 0 1.0068e-08 0.0007 1.0071e-08 0 1.0126e-08 0 1.0129e-08 0.0007 1.0132e-08 0 1.0187e-08 0 1.019e-08 0.0007 1.01931e-08 0 1.0248e-08 0 1.0251e-08 0.0007 1.0254e-08 0 1.0309e-08 0 1.0312e-08 0.0007 1.0315e-08 0 1.037e-08 0 1.0373e-08 0.0007 1.0376e-08 0 1.0431e-08 0 1.0434e-08 0.0007 1.0437e-08 0 1.0492e-08 0 1.0495e-08 0.0007 1.0498e-08 0 1.0553e-08 0 1.0556e-08 0.0007 1.0559e-08 0 1.0614e-08 0 1.0617e-08 0.0007 1.062e-08 0 1.0675e-08 0 1.0678e-08 0.0007 1.0681e-08 0 1.0736e-08 0 1.0739e-08 0.0007 1.0742e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0858e-08 0 1.0861e-08 0.0007 1.0864e-08 0 1.0919e-08 0 1.0922e-08 0.0007 1.0925e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.1041e-08 0 1.1044e-08 0.0007 1.1047e-08 0 1.1102e-08 0 1.1105e-08 0.0007 1.1108e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1224e-08 0 1.1227e-08 0.0007 1.123e-08 0 1.1285e-08 0 1.1288e-08 0.0007 1.1291e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1468e-08 0 1.1471e-08 0.0007 1.1474e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.159e-08 0 1.1593e-08 0.0007 1.1596e-08 0 1.1651e-08 0 1.1654e-08 0.0007 1.1657e-08 0 1.1712e-08 0 1.1715e-08 0.0007 1.1718e-08 0 1.1773e-08 0 1.1776e-08 0.0007 1.1779e-08 0 1.1834e-08 0 1.1837e-08 0.0007 1.184e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.1956e-08 0 1.1959e-08 0.0007 1.1962e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2078e-08 0 1.2081e-08 0.0007 1.2084e-08 0 1.2139e-08 0 1.2142e-08 0.0007 1.2145e-08 0 1.22e-08 0 1.2203e-08 0.0007 1.2206e-08 0 1.2261e-08 0 1.2264e-08 0.0007 1.2267e-08 0 1.2322e-08 0 1.2325e-08 0.0007 1.2328e-08 0 1.2383e-08 0 1.2386e-08 0.0007 1.2389e-08 0 1.2444e-08 0 1.2447e-08 0.0007 1.245e-08 0 1.2505e-08 0 1.2508e-08 0.0007 1.2511e-08 0 1.2566e-08 0 1.2569e-08 0.0007 1.2572e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2688e-08 0 1.2691e-08 0.0007 1.2694e-08 0 1.2749e-08 0 1.2752e-08 0.0007 1.2755e-08 0 1.281e-08 0 1.2813e-08 0.0007 1.2816e-08 0 1.2871e-08 0 1.2874e-08 0.0007 1.2877e-08 0 1.2932e-08 0 1.2935e-08 0.0007 1.2938e-08 0 1.2993e-08 0 1.2996e-08 0.0007 1.2999e-08 0 1.3054e-08 0 1.3057e-08 0.0007 1.306e-08 0 1.3115e-08 0 1.3118e-08 0.0007 1.3121e-08 0 1.3176e-08 0 1.3179e-08 0.0007 1.3182e-08 0 1.3237e-08 0 1.324e-08 0.0007 1.3243e-08 0 1.3298e-08 0 1.3301e-08 0.0007 1.3304e-08 0 1.3359e-08 0 1.3362e-08 0.0007 1.3365e-08 0 1.342e-08 0 1.3423e-08 0.0007 1.3426e-08 0 1.3481e-08 0 1.3484e-08 0.0007 1.3487e-08 0 1.3542e-08 0 1.3545e-08 0.0007 1.3548e-08 0 1.3603e-08 0 1.3606e-08 0.0007 1.3609e-08 0 1.3664e-08 0 1.3667e-08 0.0007 1.367e-08 0 1.3725e-08 0 1.3728e-08 0.0007 1.3731e-08 0 1.3786e-08 0 1.3789e-08 0.0007 1.3792e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.3908e-08 0 1.3911e-08 0.0007 1.3914e-08 0 1.3969e-08 0 1.3972e-08 0.0007 1.3975e-08 0 1.403e-08 0 1.4033e-08 0.0007 1.4036e-08 0 1.4091e-08 0 1.4094e-08 0.0007 1.4097e-08 0 1.4152e-08 0 1.4155e-08 0.0007 1.4158e-08 0 1.4213e-08 0 1.4216e-08 0.0007 1.4219e-08 0 1.4274e-08 0 1.4277e-08 0.0007 1.428e-08 0 1.4335e-08 0 1.4338e-08 0.0007 1.4341e-08 0 1.4396e-08 0 1.4399e-08 0.0007 1.4402e-08 0 1.4457e-08 0 1.446e-08 0.0007 1.4463e-08 0 1.4518e-08 0 1.4521e-08 0.0007 1.4524e-08 0 1.4579e-08 0 1.4582e-08 0.0007 1.4585e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.4701e-08 0 1.4704e-08 0.0007 1.4707e-08 0 1.4762e-08 0 1.4765e-08 0.0007 1.4768e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4884e-08 0 1.4887e-08 0.0007 1.489e-08 0 1.4945e-08 0 1.4948e-08 0.0007 1.4951e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5067e-08 0 1.507e-08 0.0007 1.5073e-08 0 1.5128e-08 0 1.5131e-08 0.0007 1.5134e-08 0 1.5189e-08 0 1.5192e-08 0.0007 1.5195e-08 0 1.52501e-08 0 1.52531e-08 0.0007 1.52561e-08 0 1.5311e-08 0 1.53141e-08 0.0007 1.53171e-08 0 1.5372e-08 0 1.5375e-08 0.0007 1.5378e-08 0 1.5433e-08 0 1.5436e-08 0.0007 1.5439e-08 0 1.5494e-08 0 1.5497e-08 0.0007 1.55e-08 0 1.5555e-08 0 1.5558e-08 0.0007 1.5561e-08 0 1.5616e-08 0 1.5619e-08 0.0007 1.5622e-08 0 1.5677e-08 0 1.568e-08 0.0007 1.5683e-08 0 1.5738e-08 0 1.5741e-08 0.0007 1.5744e-08 0 1.5799e-08 0 1.5802e-08 0.0007 1.5805e-08 0 1.586e-08 0 1.5863e-08 0.0007 1.5866e-08 0 1.59211e-08 0 1.59241e-08 0.0007 1.59271e-08 0 1.5982e-08 0 1.5985e-08 0.0007 1.59881e-08 0 1.6043e-08 0 1.6046e-08 0.0007 1.6049e-08 0 1.6104e-08 0 1.6107e-08 0.0007 1.611e-08 0 1.6165e-08 0 1.6168e-08 0.0007 1.6171e-08 0 1.6226e-08 0 1.6229e-08 0.0007 1.6232e-08 0 1.6287e-08 0 1.629e-08 0.0007 1.6293e-08 0 1.6348e-08 0 1.6351e-08 0.0007 1.6354e-08 0 1.6409e-08 0 1.6412e-08 0.0007 1.6415e-08 0 1.647e-08 0 1.6473e-08 0.0007 1.6476e-08 0 1.65311e-08 0 1.65341e-08 0.0007 1.65371e-08 0 1.65921e-08 0 1.65951e-08 0.0007 1.65981e-08 0 1.6653e-08 0 1.6656e-08 0.0007 1.6659e-08 0 1.6714e-08 0 1.6717e-08 0.0007 1.672e-08 0 1.6775e-08 0 1.6778e-08 0.0007 1.6781e-08 0 1.6836e-08 0 1.6839e-08 0.0007 1.6842e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6958e-08 0 1.6961e-08 0.0007 1.6964e-08 0 1.7019e-08 0 1.7022e-08 0.0007 1.7025e-08 0 1.708e-08 0 1.7083e-08 0.0007 1.7086e-08 0 1.7141e-08 0 1.7144e-08 0.0007 1.7147e-08 0 1.72021e-08 0 1.72051e-08 0.0007 1.72081e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.72691e-08 0 1.7324e-08 0 1.7327e-08 0.0007 1.733e-08 0 1.7385e-08 0 1.7388e-08 0.0007 1.7391e-08 0 1.7446e-08 0 1.7449e-08 0.0007 1.7452e-08 0 1.7507e-08 0 1.751e-08 0.0007 1.7513e-08 0 1.7568e-08 0 1.7571e-08 0.0007 1.7574e-08 0 1.7629e-08 0 1.7632e-08 0.0007 1.7635e-08 0 1.769e-08 0 1.7693e-08 0.0007 1.7696e-08 0 1.7751e-08 0 1.7754e-08 0.0007 1.7757e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.78731e-08 0 1.78761e-08 0.0007 1.78791e-08 0 1.7934e-08 0 1.7937e-08 0.0007 1.794e-08 0 1.7995e-08 0 1.7998e-08 0.0007 1.8001e-08 0 1.8056e-08 0 1.8059e-08 0.0007 1.8062e-08 0 1.8117e-08 0 1.812e-08 0.0007 1.8123e-08 0 1.8178e-08 0 1.8181e-08 0.0007 1.8184e-08 0 1.8239e-08 0 1.8242e-08 0.0007 1.8245e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.8361e-08 0 1.8364e-08 0.0007 1.8367e-08 0 1.8422e-08 0 1.8425e-08 0.0007 1.8428e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8544e-08 0 1.8547e-08 0.0007 1.85501e-08 0 1.8605e-08 0 1.8608e-08 0.0007 1.8611e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8727e-08 0 1.873e-08 0.0007 1.8733e-08 0 1.8788e-08 0 1.8791e-08 0.0007 1.8794e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.891e-08 0 1.8913e-08 0.0007 1.8916e-08 0 1.8971e-08 0 1.8974e-08 0.0007 1.8977e-08 0 1.9032e-08 0 1.9035e-08 0.0007 1.9038e-08 0 1.9093e-08 0 1.9096e-08 0.0007 1.9099e-08 0 1.91541e-08 0 1.91571e-08 0.0007 1.91601e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9276e-08 0 1.9279e-08 0.0007 1.9282e-08 0 1.9337e-08 0 1.934e-08 0.0007 1.9343e-08 0 1.9398e-08 0 1.9401e-08 0.0007 1.9404e-08 0 1.9459e-08 0 1.9462e-08 0.0007 1.9465e-08 0 1.952e-08 0 1.9523e-08 0.0007 1.9526e-08 0 1.9581e-08 0 1.9584e-08 0.0007 1.9587e-08 0 1.9642e-08 0 1.9645e-08 0.0007 1.9648e-08 0 1.9703e-08 0 1.9706e-08 0.0007 1.9709e-08 0 1.9764e-08 0 1.9767e-08 0.0007 1.977e-08 0 1.9825e-08 0 1.9828e-08 0.0007 1.98311e-08 0 1.9886e-08 0 1.9889e-08 0.0007 1.9892e-08 0 1.9947e-08 0 1.995e-08 0.0007 1.9953e-08 0 2.0008e-08 0 2.0011e-08 0.0007 2.0014e-08 0 2.0069e-08 0 2.0072e-08 0.0007 2.0075e-08 0 2.013e-08 0 2.0133e-08 0.0007 2.0136e-08 0 2.0191e-08 0 2.0194e-08 0.0007 2.0197e-08 0 2.0252e-08 0 2.0255e-08 0.0007 2.0258e-08 0 2.0313e-08 0 2.0316e-08 0.0007 2.0319e-08 0 2.0374e-08 0 2.0377e-08 0.0007 2.038e-08 0 2.04351e-08 0 2.04381e-08 0.0007 2.04411e-08 0 2.0496e-08 0 2.0499e-08 0.0007 2.0502e-08 0 2.0557e-08 0 2.056e-08 0.0007 2.0563e-08 0 2.0618e-08 0 2.0621e-08 0.0007 2.0624e-08 0 2.0679e-08 0 2.0682e-08 0.0007 2.0685e-08 0 2.074e-08 0 2.0743e-08 0.0007 2.0746e-08 0 2.0801e-08 0 2.0804e-08 0.0007 2.0807e-08 0 2.0862e-08 0 2.0865e-08 0.0007 2.0868e-08 0 2.0923e-08 0 2.0926e-08 0.0007 2.0929e-08 0 2.0984e-08 0 2.0987e-08 0.0007 2.099e-08 0 2.1045e-08 0 2.1048e-08 0.0007 2.1051e-08 0 2.1106e-08 0 2.11091e-08 0.0007 2.11121e-08 0 2.1167e-08 0 2.117e-08 0.0007 2.1173e-08 0 2.1228e-08 0 2.1231e-08 0.0007 2.1234e-08 0 2.1289e-08 0 2.1292e-08 0.0007 2.1295e-08 0 2.135e-08 0 2.1353e-08 0.0007 2.1356e-08 0 2.1411e-08 0 2.1414e-08 0.0007 2.1417e-08 0 2.1472e-08 0 2.1475e-08 0.0007 2.1478e-08 0 2.1533e-08 0 2.1536e-08 0.0007 2.1539e-08 0 2.1594e-08 0 2.1597e-08 0.0007 2.16e-08 0 2.1655e-08 0 2.1658e-08 0.0007 2.1661e-08 0 2.1716e-08 0 2.1719e-08 0.0007 2.1722e-08 0 2.1777e-08 0 2.178e-08 0.0007 2.1783e-08 0 2.1838e-08 0 2.1841e-08 0.0007 2.1844e-08 0 2.1899e-08 0 2.1902e-08 0.0007 2.1905e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.2021e-08 0 2.2024e-08 0.0007 2.2027e-08 0 2.2082e-08 0 2.2085e-08 0.0007 2.2088e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2204e-08 0 2.2207e-08 0.0007 2.221e-08 0 2.2265e-08 0 2.2268e-08 0.0007 2.2271e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2448e-08 0 2.2451e-08 0.0007 2.2454e-08 0 2.2509e-08 0 2.2512e-08 0.0007 2.2515e-08 0 2.257e-08 0 2.2573e-08 0.0007 2.2576e-08 0 2.2631e-08 0 2.2634e-08 0.0007 2.2637e-08 0 2.2692e-08 0 2.2695e-08 0.0007 2.2698e-08 0 2.2753e-08 0 2.2756e-08 0.0007 2.2759e-08 0 2.2814e-08 0 2.2817e-08 0.0007 2.282e-08 0 2.2875e-08 0 2.2878e-08 0.0007 2.2881e-08 0 2.2936e-08 0 2.2939e-08 0.0007 2.2942e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3058e-08 0 2.3061e-08 0.0007 2.3064e-08 0 2.3119e-08 0 2.3122e-08 0.0007 2.3125e-08 0 2.318e-08 0 2.3183e-08 0.0007 2.3186e-08 0 2.3241e-08 0 2.3244e-08 0.0007 2.3247e-08 0 2.3302e-08 0 2.3305e-08 0.0007 2.3308e-08 0 2.3363e-08 0 2.3366e-08 0.0007 2.3369e-08 0 2.3424e-08 0 2.3427e-08 0.0007 2.343e-08 0 2.3485e-08 0 2.3488e-08 0.0007 2.3491e-08 0 2.3546e-08 0 2.3549e-08 0.0007 2.3552e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3668e-08 0 2.3671e-08 0.0007 2.3674e-08 0 2.3729e-08 0 2.3732e-08 0.0007 2.3735e-08 0 2.379e-08 0 2.3793e-08 0.0007 2.3796e-08 0 2.3851e-08 0 2.3854e-08 0.0007 2.3857e-08 0 2.3912e-08 0 2.3915e-08 0.0007 2.3918e-08 0 2.3973e-08 0 2.3976e-08 0.0007 2.3979e-08 0 2.4034e-08 0 2.4037e-08 0.0007 2.404e-08 0 2.4095e-08 0 2.4098e-08 0.0007 2.4101e-08 0 2.4156e-08 0 2.4159e-08 0.0007 2.4162e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4278e-08 0 2.4281e-08 0.0007 2.4284e-08 0)
L_S3|A1 G2_2_RX _S3|A1  2.067833848e-12
L_S3|A2 _S3|A1 _S3|A2  4.135667696e-12
L_S3|A3 _S3|A3 _S3|AB  8.271335392e-12
L_S3|B1 IP3_2_OUT_RX _S3|B1  2.067833848e-12
L_S3|B2 _S3|B1 _S3|B2  4.135667696e-12
L_S3|B3 _S3|B3 _S3|AB  8.271335392e-12
L_S3|T1 T15 _S3|T1  2.067833848e-12
L_S3|T2 _S3|T1 _S3|T2  4.135667696e-12
L_S3|Q2 _S3|ABTQ _S3|Q1  4.135667696e-12
L_S3|Q1 _S3|Q1 S3  2.067833848e-12
IT16|T 0 T16  PWL(0 0 5e-14 0 3.05e-12 0.0007 6.05e-12 0 6.105e-11 0 6.405e-11 0.0007 6.705e-11 0 1.2205e-10 0 1.2505e-10 0.0007 1.2805e-10 0 1.8305e-10 0 1.8605e-10 0.0007 1.8905e-10 0 2.4405e-10 0 2.4705e-10 0.0007 2.5005e-10 0 3.0505e-10 0 3.0805e-10 0.0007 3.1105e-10 0 3.6605e-10 0 3.6905e-10 0.0007 3.7205e-10 0 4.2705e-10 0 4.3005e-10 0.0007 4.3305e-10 0 4.8805e-10 0 4.9105e-10 0.0007 4.9405e-10 0 5.4905e-10 0 5.5205e-10 0.0007 5.5505e-10 0 6.1005e-10 0 6.1305e-10 0.0007 6.1605e-10 0 6.7105e-10 0 6.7405e-10 0.0007 6.7705e-10 0 7.3205e-10 0 7.3505e-10 0.0007 7.3805e-10 0 7.9305e-10 0 7.9605e-10 0.0007 7.9905e-10 0 8.5405e-10 0 8.5705e-10 0.0007 8.6005e-10 0 9.1505e-10 0 9.1805e-10 0.0007 9.2105e-10 0 9.7605e-10 0 9.7905e-10 0.0007 9.8205e-10 0 1.03705e-09 0 1.04005e-09 0.0007 1.04305e-09 0 1.09805e-09 0 1.10105e-09 0.0007 1.10405e-09 0 1.15905e-09 0 1.16205e-09 0.0007 1.16505e-09 0 1.22005e-09 0 1.22305e-09 0.0007 1.22605e-09 0 1.28105e-09 0 1.28405e-09 0.0007 1.28705e-09 0 1.34205e-09 0 1.34505e-09 0.0007 1.34805e-09 0 1.40305e-09 0 1.40605e-09 0.0007 1.40905e-09 0 1.46405e-09 0 1.46705e-09 0.0007 1.47005e-09 0 1.52505e-09 0 1.52805e-09 0.0007 1.53105e-09 0 1.58605e-09 0 1.58905e-09 0.0007 1.59205e-09 0 1.64705e-09 0 1.65005e-09 0.0007 1.65305e-09 0 1.70805e-09 0 1.71105e-09 0.0007 1.71405e-09 0 1.76905e-09 0 1.77205e-09 0.0007 1.77505e-09 0 1.83005e-09 0 1.83305e-09 0.0007 1.83605e-09 0 1.89105e-09 0 1.89405e-09 0.0007 1.89705e-09 0 1.95205e-09 0 1.95505e-09 0.0007 1.95805e-09 0 2.01305e-09 0 2.01605e-09 0.0007 2.01905e-09 0 2.07405e-09 0 2.07705e-09 0.0007 2.08005e-09 0 2.13505e-09 0 2.13805e-09 0.0007 2.14105e-09 0 2.19605e-09 0 2.19905e-09 0.0007 2.20205e-09 0 2.25705e-09 0 2.26005e-09 0.0007 2.26305e-09 0 2.31805e-09 0 2.32105e-09 0.0007 2.32405e-09 0 2.37905e-09 0 2.38205e-09 0.0007 2.38505e-09 0 2.44005e-09 0 2.44305e-09 0.0007 2.44605e-09 0 2.50105e-09 0 2.50405e-09 0.0007 2.50705e-09 0 2.56205e-09 0 2.56505e-09 0.0007 2.56805e-09 0 2.62305e-09 0 2.62605e-09 0.0007 2.62905e-09 0 2.68405e-09 0 2.68705e-09 0.0007 2.69005e-09 0 2.74505e-09 0 2.74805e-09 0.0007 2.75105e-09 0 2.80605e-09 0 2.80905e-09 0.0007 2.81205e-09 0 2.86705e-09 0 2.87005e-09 0.0007 2.87305e-09 0 2.92805e-09 0 2.93105e-09 0.0007 2.93405e-09 0 2.98905e-09 0 2.99205e-09 0.0007 2.99505e-09 0 3.05005e-09 0 3.05305e-09 0.0007 3.05605e-09 0 3.11105e-09 0 3.11405e-09 0.0007 3.11705e-09 0 3.17205e-09 0 3.17505e-09 0.0007 3.17805e-09 0 3.23305e-09 0 3.23605e-09 0.0007 3.23905e-09 0 3.29405e-09 0 3.29705e-09 0.0007 3.30005e-09 0 3.35505e-09 0 3.35805e-09 0.0007 3.36105e-09 0 3.41605e-09 0 3.41905e-09 0.0007 3.42205e-09 0 3.47705e-09 0 3.48005e-09 0.0007 3.48305e-09 0 3.53805e-09 0 3.54105e-09 0.0007 3.54405e-09 0 3.59905e-09 0 3.60205e-09 0.0007 3.60505e-09 0 3.66005e-09 0 3.66305e-09 0.0007 3.66605e-09 0 3.72105e-09 0 3.72405e-09 0.0007 3.72705e-09 0 3.78205e-09 0 3.78505e-09 0.0007 3.78805e-09 0 3.84305e-09 0 3.84605e-09 0.0007 3.84905e-09 0 3.90405e-09 0 3.90705e-09 0.0007 3.91005e-09 0 3.96505e-09 0 3.96805e-09 0.0007 3.97105e-09 0 4.02605e-09 0 4.02905e-09 0.0007 4.03205e-09 0 4.08705e-09 0 4.09005e-09 0.0007 4.09305e-09 0 4.14805e-09 0 4.15105e-09 0.0007 4.15405e-09 0 4.20905e-09 0 4.21205e-09 0.0007 4.21505e-09 0 4.27005e-09 0 4.27305e-09 0.0007 4.27605e-09 0 4.33105e-09 0 4.33405e-09 0.0007 4.33705e-09 0 4.39205e-09 0 4.39505e-09 0.0007 4.39805e-09 0 4.45305e-09 0 4.45605e-09 0.0007 4.45905e-09 0 4.51405e-09 0 4.51705e-09 0.0007 4.52005e-09 0 4.57505e-09 0 4.57805e-09 0.0007 4.58105e-09 0 4.63605e-09 0 4.63905e-09 0.0007 4.64205e-09 0 4.69705e-09 0 4.70005e-09 0.0007 4.70305e-09 0 4.75805e-09 0 4.76105e-09 0.0007 4.76405e-09 0 4.81905e-09 0 4.82205e-09 0.0007 4.82505e-09 0 4.88005e-09 0 4.88305e-09 0.0007 4.88605e-09 0 4.94105e-09 0 4.94405e-09 0.0007 4.94705e-09 0 5.00205e-09 0 5.00505e-09 0.0007 5.00805e-09 0 5.06305e-09 0 5.06605e-09 0.0007 5.06905e-09 0 5.12405e-09 0 5.12705e-09 0.0007 5.13005e-09 0 5.18505e-09 0 5.18805e-09 0.0007 5.19105e-09 0 5.24605e-09 0 5.24905e-09 0.0007 5.25205e-09 0 5.30705e-09 0 5.31005e-09 0.0007 5.31305e-09 0 5.36805e-09 0 5.37105e-09 0.0007 5.37405e-09 0 5.42905e-09 0 5.43205e-09 0.0007 5.43505e-09 0 5.49005e-09 0 5.49305e-09 0.0007 5.49605e-09 0 5.55105e-09 0 5.55405e-09 0.0007 5.55705e-09 0 5.61205e-09 0 5.61505e-09 0.0007 5.61805e-09 0 5.67305e-09 0 5.67605e-09 0.0007 5.67905e-09 0 5.73405e-09 0 5.73705e-09 0.0007 5.74005e-09 0 5.79505e-09 0 5.79805e-09 0.0007 5.80105e-09 0 5.85605e-09 0 5.85905e-09 0.0007 5.86205e-09 0 5.91705e-09 0 5.92005e-09 0.0007 5.92305e-09 0 5.97805e-09 0 5.98105e-09 0.0007 5.98405e-09 0 6.03905e-09 0 6.04205e-09 0.0007 6.04505e-09 0 6.10005e-09 0 6.10305e-09 0.0007 6.10605e-09 0 6.16105e-09 0 6.16405e-09 0.0007 6.16705e-09 0 6.22205e-09 0 6.22505e-09 0.0007 6.22805e-09 0 6.28305e-09 0 6.28605e-09 0.0007 6.28905e-09 0 6.34405e-09 0 6.34705e-09 0.0007 6.35005e-09 0 6.40505e-09 0 6.40805e-09 0.0007 6.41105e-09 0 6.46605e-09 0 6.46905e-09 0.0007 6.47205e-09 0 6.52705e-09 0 6.53005e-09 0.0007 6.53305e-09 0 6.58805e-09 0 6.59105e-09 0.0007 6.59405e-09 0 6.64905e-09 0 6.65205e-09 0.0007 6.65505e-09 0 6.71005e-09 0 6.71305e-09 0.0007 6.71605e-09 0 6.77105e-09 0 6.77405e-09 0.0007 6.77705e-09 0 6.83205e-09 0 6.83505e-09 0.0007 6.83805e-09 0 6.89305e-09 0 6.89605e-09 0.0007 6.89905e-09 0 6.95405e-09 0 6.95705e-09 0.0007 6.96005e-09 0 7.01505e-09 0 7.01805e-09 0.0007 7.02105e-09 0 7.07605e-09 0 7.07905e-09 0.0007 7.08205e-09 0 7.13705e-09 0 7.14005e-09 0.0007 7.14305e-09 0 7.19805e-09 0 7.20105e-09 0.0007 7.20405e-09 0 7.25905e-09 0 7.26205e-09 0.0007 7.26505e-09 0 7.32005e-09 0 7.32305e-09 0.0007 7.32605e-09 0 7.38105e-09 0 7.38405e-09 0.0007 7.38705e-09 0 7.44205e-09 0 7.44505e-09 0.0007 7.44805e-09 0 7.50305e-09 0 7.50605e-09 0.0007 7.50905e-09 0 7.56405e-09 0 7.56705e-09 0.0007 7.57005e-09 0 7.62505e-09 0 7.62805e-09 0.0007 7.63105e-09 0 7.68605e-09 0 7.68905e-09 0.0007 7.69205e-09 0 7.74705e-09 0 7.75005e-09 0.0007 7.75305e-09 0 7.80805e-09 0 7.81105e-09 0.0007 7.81405e-09 0 7.86905e-09 0 7.87205e-09 0.0007 7.87505e-09 0 7.93005e-09 0 7.93305e-09 0.0007 7.93605e-09 0 7.99105e-09 0 7.99405e-09 0.0007 7.99705e-09 0 8.05205e-09 0 8.05505e-09 0.0007 8.05805e-09 0 8.11305e-09 0 8.11605e-09 0.0007 8.11905e-09 0 8.17405e-09 0 8.17705e-09 0.0007 8.18005e-09 0 8.23505e-09 0 8.23805e-09 0.0007 8.24105e-09 0 8.29605e-09 0 8.29905e-09 0.0007 8.30205e-09 0 8.35705e-09 0 8.36005e-09 0.0007 8.36305e-09 0 8.41805e-09 0 8.42105e-09 0.0007 8.42405e-09 0 8.47905e-09 0 8.48205e-09 0.0007 8.48505e-09 0 8.54005e-09 0 8.54305e-09 0.0007 8.54605e-09 0 8.60105e-09 0 8.60405e-09 0.0007 8.60705e-09 0 8.66205e-09 0 8.66505e-09 0.0007 8.66805e-09 0 8.72305e-09 0 8.72605e-09 0.0007 8.72905e-09 0 8.78405e-09 0 8.78705e-09 0.0007 8.79005e-09 0 8.84505e-09 0 8.84805e-09 0.0007 8.85105e-09 0 8.90605e-09 0 8.90905e-09 0.0007 8.91205e-09 0 8.96705e-09 0 8.97005e-09 0.0007 8.97305e-09 0 9.02805e-09 0 9.03105e-09 0.0007 9.03405e-09 0 9.08905e-09 0 9.09205e-09 0.0007 9.09505e-09 0 9.15005e-09 0 9.15305e-09 0.0007 9.15605e-09 0 9.21105e-09 0 9.21405e-09 0.0007 9.21705e-09 0 9.27205e-09 0 9.27505e-09 0.0007 9.27805e-09 0 9.33305e-09 0 9.33605e-09 0.0007 9.33905e-09 0 9.39405e-09 0 9.39705e-09 0.0007 9.40005e-09 0 9.45505e-09 0 9.45805e-09 0.0007 9.46105e-09 0 9.51605e-09 0 9.51905e-09 0.0007 9.52205e-09 0 9.57705e-09 0 9.58005e-09 0.0007 9.58305e-09 0 9.63805e-09 0 9.64105e-09 0.0007 9.64405e-09 0 9.69905e-09 0 9.70205e-09 0.0007 9.70505e-09 0 9.76005e-09 0 9.76305e-09 0.0007 9.76605e-09 0 9.82105e-09 0 9.82405e-09 0.0007 9.82705e-09 0 9.88205e-09 0 9.88505e-09 0.0007 9.88805e-09 0 9.94305e-09 0 9.94605e-09 0.0007 9.94905e-09 0 1.0004e-08 0 1.0007e-08 0.0007 1.001e-08 0 1.0065e-08 0 1.0068e-08 0.0007 1.0071e-08 0 1.0126e-08 0 1.0129e-08 0.0007 1.0132e-08 0 1.0187e-08 0 1.019e-08 0.0007 1.01931e-08 0 1.0248e-08 0 1.0251e-08 0.0007 1.0254e-08 0 1.0309e-08 0 1.0312e-08 0.0007 1.0315e-08 0 1.037e-08 0 1.0373e-08 0.0007 1.0376e-08 0 1.0431e-08 0 1.0434e-08 0.0007 1.0437e-08 0 1.0492e-08 0 1.0495e-08 0.0007 1.0498e-08 0 1.0553e-08 0 1.0556e-08 0.0007 1.0559e-08 0 1.0614e-08 0 1.0617e-08 0.0007 1.062e-08 0 1.0675e-08 0 1.0678e-08 0.0007 1.0681e-08 0 1.0736e-08 0 1.0739e-08 0.0007 1.0742e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0858e-08 0 1.0861e-08 0.0007 1.0864e-08 0 1.0919e-08 0 1.0922e-08 0.0007 1.0925e-08 0 1.098e-08 0 1.0983e-08 0.0007 1.0986e-08 0 1.1041e-08 0 1.1044e-08 0.0007 1.1047e-08 0 1.1102e-08 0 1.1105e-08 0.0007 1.1108e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1224e-08 0 1.1227e-08 0.0007 1.123e-08 0 1.1285e-08 0 1.1288e-08 0.0007 1.1291e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1468e-08 0 1.1471e-08 0.0007 1.1474e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.159e-08 0 1.1593e-08 0.0007 1.1596e-08 0 1.1651e-08 0 1.1654e-08 0.0007 1.1657e-08 0 1.1712e-08 0 1.1715e-08 0.0007 1.1718e-08 0 1.1773e-08 0 1.1776e-08 0.0007 1.1779e-08 0 1.1834e-08 0 1.1837e-08 0.0007 1.184e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.1956e-08 0 1.1959e-08 0.0007 1.1962e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2078e-08 0 1.2081e-08 0.0007 1.2084e-08 0 1.2139e-08 0 1.2142e-08 0.0007 1.2145e-08 0 1.22e-08 0 1.2203e-08 0.0007 1.2206e-08 0 1.2261e-08 0 1.2264e-08 0.0007 1.2267e-08 0 1.2322e-08 0 1.2325e-08 0.0007 1.2328e-08 0 1.2383e-08 0 1.2386e-08 0.0007 1.2389e-08 0 1.2444e-08 0 1.2447e-08 0.0007 1.245e-08 0 1.2505e-08 0 1.2508e-08 0.0007 1.2511e-08 0 1.2566e-08 0 1.2569e-08 0.0007 1.2572e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2688e-08 0 1.2691e-08 0.0007 1.2694e-08 0 1.2749e-08 0 1.2752e-08 0.0007 1.2755e-08 0 1.281e-08 0 1.2813e-08 0.0007 1.2816e-08 0 1.2871e-08 0 1.2874e-08 0.0007 1.2877e-08 0 1.2932e-08 0 1.2935e-08 0.0007 1.2938e-08 0 1.2993e-08 0 1.2996e-08 0.0007 1.2999e-08 0 1.3054e-08 0 1.3057e-08 0.0007 1.306e-08 0 1.3115e-08 0 1.3118e-08 0.0007 1.3121e-08 0 1.3176e-08 0 1.3179e-08 0.0007 1.3182e-08 0 1.3237e-08 0 1.324e-08 0.0007 1.3243e-08 0 1.3298e-08 0 1.3301e-08 0.0007 1.3304e-08 0 1.3359e-08 0 1.3362e-08 0.0007 1.3365e-08 0 1.342e-08 0 1.3423e-08 0.0007 1.3426e-08 0 1.3481e-08 0 1.3484e-08 0.0007 1.3487e-08 0 1.3542e-08 0 1.3545e-08 0.0007 1.3548e-08 0 1.3603e-08 0 1.3606e-08 0.0007 1.3609e-08 0 1.3664e-08 0 1.3667e-08 0.0007 1.367e-08 0 1.3725e-08 0 1.3728e-08 0.0007 1.3731e-08 0 1.3786e-08 0 1.3789e-08 0.0007 1.3792e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.3908e-08 0 1.3911e-08 0.0007 1.3914e-08 0 1.3969e-08 0 1.3972e-08 0.0007 1.3975e-08 0 1.403e-08 0 1.4033e-08 0.0007 1.4036e-08 0 1.4091e-08 0 1.4094e-08 0.0007 1.4097e-08 0 1.4152e-08 0 1.4155e-08 0.0007 1.4158e-08 0 1.4213e-08 0 1.4216e-08 0.0007 1.4219e-08 0 1.4274e-08 0 1.4277e-08 0.0007 1.428e-08 0 1.4335e-08 0 1.4338e-08 0.0007 1.4341e-08 0 1.4396e-08 0 1.4399e-08 0.0007 1.4402e-08 0 1.4457e-08 0 1.446e-08 0.0007 1.4463e-08 0 1.4518e-08 0 1.4521e-08 0.0007 1.4524e-08 0 1.4579e-08 0 1.4582e-08 0.0007 1.4585e-08 0 1.464e-08 0 1.4643e-08 0.0007 1.4646e-08 0 1.4701e-08 0 1.4704e-08 0.0007 1.4707e-08 0 1.4762e-08 0 1.4765e-08 0.0007 1.4768e-08 0 1.4823e-08 0 1.4826e-08 0.0007 1.4829e-08 0 1.4884e-08 0 1.4887e-08 0.0007 1.489e-08 0 1.4945e-08 0 1.4948e-08 0.0007 1.4951e-08 0 1.5006e-08 0 1.5009e-08 0.0007 1.5012e-08 0 1.5067e-08 0 1.507e-08 0.0007 1.5073e-08 0 1.5128e-08 0 1.5131e-08 0.0007 1.5134e-08 0 1.5189e-08 0 1.5192e-08 0.0007 1.5195e-08 0 1.52501e-08 0 1.52531e-08 0.0007 1.52561e-08 0 1.5311e-08 0 1.53141e-08 0.0007 1.53171e-08 0 1.5372e-08 0 1.5375e-08 0.0007 1.5378e-08 0 1.5433e-08 0 1.5436e-08 0.0007 1.5439e-08 0 1.5494e-08 0 1.5497e-08 0.0007 1.55e-08 0 1.5555e-08 0 1.5558e-08 0.0007 1.5561e-08 0 1.5616e-08 0 1.5619e-08 0.0007 1.5622e-08 0 1.5677e-08 0 1.568e-08 0.0007 1.5683e-08 0 1.5738e-08 0 1.5741e-08 0.0007 1.5744e-08 0 1.5799e-08 0 1.5802e-08 0.0007 1.5805e-08 0 1.586e-08 0 1.5863e-08 0.0007 1.5866e-08 0 1.59211e-08 0 1.59241e-08 0.0007 1.59271e-08 0 1.5982e-08 0 1.5985e-08 0.0007 1.59881e-08 0 1.6043e-08 0 1.6046e-08 0.0007 1.6049e-08 0 1.6104e-08 0 1.6107e-08 0.0007 1.611e-08 0 1.6165e-08 0 1.6168e-08 0.0007 1.6171e-08 0 1.6226e-08 0 1.6229e-08 0.0007 1.6232e-08 0 1.6287e-08 0 1.629e-08 0.0007 1.6293e-08 0 1.6348e-08 0 1.6351e-08 0.0007 1.6354e-08 0 1.6409e-08 0 1.6412e-08 0.0007 1.6415e-08 0 1.647e-08 0 1.6473e-08 0.0007 1.6476e-08 0 1.65311e-08 0 1.65341e-08 0.0007 1.65371e-08 0 1.65921e-08 0 1.65951e-08 0.0007 1.65981e-08 0 1.6653e-08 0 1.6656e-08 0.0007 1.6659e-08 0 1.6714e-08 0 1.6717e-08 0.0007 1.672e-08 0 1.6775e-08 0 1.6778e-08 0.0007 1.6781e-08 0 1.6836e-08 0 1.6839e-08 0.0007 1.6842e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6958e-08 0 1.6961e-08 0.0007 1.6964e-08 0 1.7019e-08 0 1.7022e-08 0.0007 1.7025e-08 0 1.708e-08 0 1.7083e-08 0.0007 1.7086e-08 0 1.7141e-08 0 1.7144e-08 0.0007 1.7147e-08 0 1.72021e-08 0 1.72051e-08 0.0007 1.72081e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.72691e-08 0 1.7324e-08 0 1.7327e-08 0.0007 1.733e-08 0 1.7385e-08 0 1.7388e-08 0.0007 1.7391e-08 0 1.7446e-08 0 1.7449e-08 0.0007 1.7452e-08 0 1.7507e-08 0 1.751e-08 0.0007 1.7513e-08 0 1.7568e-08 0 1.7571e-08 0.0007 1.7574e-08 0 1.7629e-08 0 1.7632e-08 0.0007 1.7635e-08 0 1.769e-08 0 1.7693e-08 0.0007 1.7696e-08 0 1.7751e-08 0 1.7754e-08 0.0007 1.7757e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.78731e-08 0 1.78761e-08 0.0007 1.78791e-08 0 1.7934e-08 0 1.7937e-08 0.0007 1.794e-08 0 1.7995e-08 0 1.7998e-08 0.0007 1.8001e-08 0 1.8056e-08 0 1.8059e-08 0.0007 1.8062e-08 0 1.8117e-08 0 1.812e-08 0.0007 1.8123e-08 0 1.8178e-08 0 1.8181e-08 0.0007 1.8184e-08 0 1.8239e-08 0 1.8242e-08 0.0007 1.8245e-08 0 1.83e-08 0 1.8303e-08 0.0007 1.8306e-08 0 1.8361e-08 0 1.8364e-08 0.0007 1.8367e-08 0 1.8422e-08 0 1.8425e-08 0.0007 1.8428e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8544e-08 0 1.8547e-08 0.0007 1.85501e-08 0 1.8605e-08 0 1.8608e-08 0.0007 1.8611e-08 0 1.8666e-08 0 1.8669e-08 0.0007 1.8672e-08 0 1.8727e-08 0 1.873e-08 0.0007 1.8733e-08 0 1.8788e-08 0 1.8791e-08 0.0007 1.8794e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.891e-08 0 1.8913e-08 0.0007 1.8916e-08 0 1.8971e-08 0 1.8974e-08 0.0007 1.8977e-08 0 1.9032e-08 0 1.9035e-08 0.0007 1.9038e-08 0 1.9093e-08 0 1.9096e-08 0.0007 1.9099e-08 0 1.91541e-08 0 1.91571e-08 0.0007 1.91601e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9276e-08 0 1.9279e-08 0.0007 1.9282e-08 0 1.9337e-08 0 1.934e-08 0.0007 1.9343e-08 0 1.9398e-08 0 1.9401e-08 0.0007 1.9404e-08 0 1.9459e-08 0 1.9462e-08 0.0007 1.9465e-08 0 1.952e-08 0 1.9523e-08 0.0007 1.9526e-08 0 1.9581e-08 0 1.9584e-08 0.0007 1.9587e-08 0 1.9642e-08 0 1.9645e-08 0.0007 1.9648e-08 0 1.9703e-08 0 1.9706e-08 0.0007 1.9709e-08 0 1.9764e-08 0 1.9767e-08 0.0007 1.977e-08 0 1.9825e-08 0 1.9828e-08 0.0007 1.98311e-08 0 1.9886e-08 0 1.9889e-08 0.0007 1.9892e-08 0 1.9947e-08 0 1.995e-08 0.0007 1.9953e-08 0 2.0008e-08 0 2.0011e-08 0.0007 2.0014e-08 0 2.0069e-08 0 2.0072e-08 0.0007 2.0075e-08 0 2.013e-08 0 2.0133e-08 0.0007 2.0136e-08 0 2.0191e-08 0 2.0194e-08 0.0007 2.0197e-08 0 2.0252e-08 0 2.0255e-08 0.0007 2.0258e-08 0 2.0313e-08 0 2.0316e-08 0.0007 2.0319e-08 0 2.0374e-08 0 2.0377e-08 0.0007 2.038e-08 0 2.04351e-08 0 2.04381e-08 0.0007 2.04411e-08 0 2.0496e-08 0 2.0499e-08 0.0007 2.0502e-08 0 2.0557e-08 0 2.056e-08 0.0007 2.0563e-08 0 2.0618e-08 0 2.0621e-08 0.0007 2.0624e-08 0 2.0679e-08 0 2.0682e-08 0.0007 2.0685e-08 0 2.074e-08 0 2.0743e-08 0.0007 2.0746e-08 0 2.0801e-08 0 2.0804e-08 0.0007 2.0807e-08 0 2.0862e-08 0 2.0865e-08 0.0007 2.0868e-08 0 2.0923e-08 0 2.0926e-08 0.0007 2.0929e-08 0 2.0984e-08 0 2.0987e-08 0.0007 2.099e-08 0 2.1045e-08 0 2.1048e-08 0.0007 2.1051e-08 0 2.1106e-08 0 2.11091e-08 0.0007 2.11121e-08 0 2.1167e-08 0 2.117e-08 0.0007 2.1173e-08 0 2.1228e-08 0 2.1231e-08 0.0007 2.1234e-08 0 2.1289e-08 0 2.1292e-08 0.0007 2.1295e-08 0 2.135e-08 0 2.1353e-08 0.0007 2.1356e-08 0 2.1411e-08 0 2.1414e-08 0.0007 2.1417e-08 0 2.1472e-08 0 2.1475e-08 0.0007 2.1478e-08 0 2.1533e-08 0 2.1536e-08 0.0007 2.1539e-08 0 2.1594e-08 0 2.1597e-08 0.0007 2.16e-08 0 2.1655e-08 0 2.1658e-08 0.0007 2.1661e-08 0 2.1716e-08 0 2.1719e-08 0.0007 2.1722e-08 0 2.1777e-08 0 2.178e-08 0.0007 2.1783e-08 0 2.1838e-08 0 2.1841e-08 0.0007 2.1844e-08 0 2.1899e-08 0 2.1902e-08 0.0007 2.1905e-08 0 2.196e-08 0 2.1963e-08 0.0007 2.1966e-08 0 2.2021e-08 0 2.2024e-08 0.0007 2.2027e-08 0 2.2082e-08 0 2.2085e-08 0.0007 2.2088e-08 0 2.2143e-08 0 2.2146e-08 0.0007 2.2149e-08 0 2.2204e-08 0 2.2207e-08 0.0007 2.221e-08 0 2.2265e-08 0 2.2268e-08 0.0007 2.2271e-08 0 2.2326e-08 0 2.2329e-08 0.0007 2.2332e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2448e-08 0 2.2451e-08 0.0007 2.2454e-08 0 2.2509e-08 0 2.2512e-08 0.0007 2.2515e-08 0 2.257e-08 0 2.2573e-08 0.0007 2.2576e-08 0 2.2631e-08 0 2.2634e-08 0.0007 2.2637e-08 0 2.2692e-08 0 2.2695e-08 0.0007 2.2698e-08 0 2.2753e-08 0 2.2756e-08 0.0007 2.2759e-08 0 2.2814e-08 0 2.2817e-08 0.0007 2.282e-08 0 2.2875e-08 0 2.2878e-08 0.0007 2.2881e-08 0 2.2936e-08 0 2.2939e-08 0.0007 2.2942e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3058e-08 0 2.3061e-08 0.0007 2.3064e-08 0 2.3119e-08 0 2.3122e-08 0.0007 2.3125e-08 0 2.318e-08 0 2.3183e-08 0.0007 2.3186e-08 0 2.3241e-08 0 2.3244e-08 0.0007 2.3247e-08 0 2.3302e-08 0 2.3305e-08 0.0007 2.3308e-08 0 2.3363e-08 0 2.3366e-08 0.0007 2.3369e-08 0 2.3424e-08 0 2.3427e-08 0.0007 2.343e-08 0 2.3485e-08 0 2.3488e-08 0.0007 2.3491e-08 0 2.3546e-08 0 2.3549e-08 0.0007 2.3552e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3668e-08 0 2.3671e-08 0.0007 2.3674e-08 0 2.3729e-08 0 2.3732e-08 0.0007 2.3735e-08 0 2.379e-08 0 2.3793e-08 0.0007 2.3796e-08 0 2.3851e-08 0 2.3854e-08 0.0007 2.3857e-08 0 2.3912e-08 0 2.3915e-08 0.0007 2.3918e-08 0 2.3973e-08 0 2.3976e-08 0.0007 2.3979e-08 0 2.4034e-08 0 2.4037e-08 0.0007 2.404e-08 0 2.4095e-08 0 2.4098e-08 0.0007 2.4101e-08 0 2.4156e-08 0 2.4159e-08 0.0007 2.4162e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4278e-08 0 2.4281e-08 0.0007 2.4284e-08 0)
L_S4|1 G3_2_RX _S4|A1  2.067833848e-12
L_S4|2 _S4|A1 _S4|A2  4.135667696e-12
L_S4|3 _S4|A3 _S4|A4  8.271335392e-12
L_S4|T T16 _S4|T1  2.067833848e-12
L_S4|4 _S4|T1 _S4|T2  4.135667696e-12
L_S4|5 _S4|A4 _S4|Q1  4.135667696e-12
L_S4|6 _S4|Q1 S4  2.067833848e-12
B_PTL_A0|_TX|1 _PTL_A0|_TX|1 _PTL_A0|_TX|2 JJMIT AREA=2.5
B_PTL_A0|_TX|2 _PTL_A0|_TX|4 _PTL_A0|_TX|5 JJMIT AREA=2.5
I_PTL_A0|_TX|B1 0 _PTL_A0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A0|_TX|B2 0 _PTL_A0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|3  1.684e-12
L_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|6  3.596e-12
L_PTL_A0|_TX|1 A0 _PTL_A0|_TX|1  2.063e-12
L_PTL_A0|_TX|2 _PTL_A0|_TX|1 _PTL_A0|_TX|4  4.123e-12
L_PTL_A0|_TX|3 _PTL_A0|_TX|4 _PTL_A0|_TX|7  2.193e-12
R_PTL_A0|_TX|D _PTL_A0|_TX|7 _PTL_A0|A_PTL  1.36
L_PTL_A0|_TX|P1 _PTL_A0|_TX|2 0  5.254e-13
L_PTL_A0|_TX|P2 _PTL_A0|_TX|5 0  5.141e-13
R_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|101  2.7439617672
R_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|104  2.7439617672
L_PTL_A0|_TX|RB1 _PTL_A0|_TX|101 0  1.550338398468e-12
L_PTL_A0|_TX|RB2 _PTL_A0|_TX|104 0  1.550338398468e-12
B_PTL_A0|_RX|1 _PTL_A0|_RX|1 _PTL_A0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A0|_RX|2 _PTL_A0|_RX|4 _PTL_A0|_RX|5 JJMIT AREA=2.0
B_PTL_A0|_RX|3 _PTL_A0|_RX|7 _PTL_A0|_RX|8 JJMIT AREA=2.5
I_PTL_A0|_RX|B1 0 _PTL_A0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|3  2.777e-12
I_PTL_A0|_RX|B2 0 _PTL_A0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|6  2.685e-12
I_PTL_A0|_RX|B3 0 _PTL_A0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|9  2.764e-12
L_PTL_A0|_RX|1 _PTL_A0|A_PTL _PTL_A0|_RX|1  1.346e-12
L_PTL_A0|_RX|2 _PTL_A0|_RX|1 _PTL_A0|_RX|4  6.348e-12
L_PTL_A0|_RX|3 _PTL_A0|_RX|4 _PTL_A0|_RX|7  5.197e-12
L_PTL_A0|_RX|4 _PTL_A0|_RX|7 A0_RX  2.058e-12
L_PTL_A0|_RX|P1 _PTL_A0|_RX|2 0  4.795e-13
L_PTL_A0|_RX|P2 _PTL_A0|_RX|5 0  5.431e-13
L_PTL_A0|_RX|P3 _PTL_A0|_RX|8 0  5.339e-13
R_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|101  4.225701121488
R_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|104  3.429952209
R_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|107  2.7439617672
L_PTL_A0|_RX|RB1 _PTL_A0|_RX|101 0  2.38752113364072e-12
L_PTL_A0|_RX|RB2 _PTL_A0|_RX|104 0  1.937922998085e-12
L_PTL_A0|_RX|RB3 _PTL_A0|_RX|107 0  1.550338398468e-12
B_PTL_B0|_TX|1 _PTL_B0|_TX|1 _PTL_B0|_TX|2 JJMIT AREA=2.5
B_PTL_B0|_TX|2 _PTL_B0|_TX|4 _PTL_B0|_TX|5 JJMIT AREA=2.5
I_PTL_B0|_TX|B1 0 _PTL_B0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B0|_TX|B2 0 _PTL_B0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|3  1.684e-12
L_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|6  3.596e-12
L_PTL_B0|_TX|1 B0 _PTL_B0|_TX|1  2.063e-12
L_PTL_B0|_TX|2 _PTL_B0|_TX|1 _PTL_B0|_TX|4  4.123e-12
L_PTL_B0|_TX|3 _PTL_B0|_TX|4 _PTL_B0|_TX|7  2.193e-12
R_PTL_B0|_TX|D _PTL_B0|_TX|7 _PTL_B0|A_PTL  1.36
L_PTL_B0|_TX|P1 _PTL_B0|_TX|2 0  5.254e-13
L_PTL_B0|_TX|P2 _PTL_B0|_TX|5 0  5.141e-13
R_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|101  2.7439617672
R_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|104  2.7439617672
L_PTL_B0|_TX|RB1 _PTL_B0|_TX|101 0  1.550338398468e-12
L_PTL_B0|_TX|RB2 _PTL_B0|_TX|104 0  1.550338398468e-12
B_PTL_B0|_RX|1 _PTL_B0|_RX|1 _PTL_B0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B0|_RX|2 _PTL_B0|_RX|4 _PTL_B0|_RX|5 JJMIT AREA=2.0
B_PTL_B0|_RX|3 _PTL_B0|_RX|7 _PTL_B0|_RX|8 JJMIT AREA=2.5
I_PTL_B0|_RX|B1 0 _PTL_B0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|3  2.777e-12
I_PTL_B0|_RX|B2 0 _PTL_B0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|6  2.685e-12
I_PTL_B0|_RX|B3 0 _PTL_B0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|9  2.764e-12
L_PTL_B0|_RX|1 _PTL_B0|A_PTL _PTL_B0|_RX|1  1.346e-12
L_PTL_B0|_RX|2 _PTL_B0|_RX|1 _PTL_B0|_RX|4  6.348e-12
L_PTL_B0|_RX|3 _PTL_B0|_RX|4 _PTL_B0|_RX|7  5.197e-12
L_PTL_B0|_RX|4 _PTL_B0|_RX|7 B0_RX  2.058e-12
L_PTL_B0|_RX|P1 _PTL_B0|_RX|2 0  4.795e-13
L_PTL_B0|_RX|P2 _PTL_B0|_RX|5 0  5.431e-13
L_PTL_B0|_RX|P3 _PTL_B0|_RX|8 0  5.339e-13
R_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|101  4.225701121488
R_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|104  3.429952209
R_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|107  2.7439617672
L_PTL_B0|_RX|RB1 _PTL_B0|_RX|101 0  2.38752113364072e-12
L_PTL_B0|_RX|RB2 _PTL_B0|_RX|104 0  1.937922998085e-12
L_PTL_B0|_RX|RB3 _PTL_B0|_RX|107 0  1.550338398468e-12
B_PTL_A1|_TX|1 _PTL_A1|_TX|1 _PTL_A1|_TX|2 JJMIT AREA=2.5
B_PTL_A1|_TX|2 _PTL_A1|_TX|4 _PTL_A1|_TX|5 JJMIT AREA=2.5
I_PTL_A1|_TX|B1 0 _PTL_A1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A1|_TX|B2 0 _PTL_A1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|3  1.684e-12
L_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|6  3.596e-12
L_PTL_A1|_TX|1 A1 _PTL_A1|_TX|1  2.063e-12
L_PTL_A1|_TX|2 _PTL_A1|_TX|1 _PTL_A1|_TX|4  4.123e-12
L_PTL_A1|_TX|3 _PTL_A1|_TX|4 _PTL_A1|_TX|7  2.193e-12
R_PTL_A1|_TX|D _PTL_A1|_TX|7 _PTL_A1|A_PTL  1.36
L_PTL_A1|_TX|P1 _PTL_A1|_TX|2 0  5.254e-13
L_PTL_A1|_TX|P2 _PTL_A1|_TX|5 0  5.141e-13
R_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|101  2.7439617672
R_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|104  2.7439617672
L_PTL_A1|_TX|RB1 _PTL_A1|_TX|101 0  1.550338398468e-12
L_PTL_A1|_TX|RB2 _PTL_A1|_TX|104 0  1.550338398468e-12
B_PTL_A1|_RX|1 _PTL_A1|_RX|1 _PTL_A1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A1|_RX|2 _PTL_A1|_RX|4 _PTL_A1|_RX|5 JJMIT AREA=2.0
B_PTL_A1|_RX|3 _PTL_A1|_RX|7 _PTL_A1|_RX|8 JJMIT AREA=2.5
I_PTL_A1|_RX|B1 0 _PTL_A1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|3  2.777e-12
I_PTL_A1|_RX|B2 0 _PTL_A1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|6  2.685e-12
I_PTL_A1|_RX|B3 0 _PTL_A1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|9  2.764e-12
L_PTL_A1|_RX|1 _PTL_A1|A_PTL _PTL_A1|_RX|1  1.346e-12
L_PTL_A1|_RX|2 _PTL_A1|_RX|1 _PTL_A1|_RX|4  6.348e-12
L_PTL_A1|_RX|3 _PTL_A1|_RX|4 _PTL_A1|_RX|7  5.197e-12
L_PTL_A1|_RX|4 _PTL_A1|_RX|7 A1_RX  2.058e-12
L_PTL_A1|_RX|P1 _PTL_A1|_RX|2 0  4.795e-13
L_PTL_A1|_RX|P2 _PTL_A1|_RX|5 0  5.431e-13
L_PTL_A1|_RX|P3 _PTL_A1|_RX|8 0  5.339e-13
R_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|101  4.225701121488
R_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|104  3.429952209
R_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|107  2.7439617672
L_PTL_A1|_RX|RB1 _PTL_A1|_RX|101 0  2.38752113364072e-12
L_PTL_A1|_RX|RB2 _PTL_A1|_RX|104 0  1.937922998085e-12
L_PTL_A1|_RX|RB3 _PTL_A1|_RX|107 0  1.550338398468e-12
B_PTL_B1|_TX|1 _PTL_B1|_TX|1 _PTL_B1|_TX|2 JJMIT AREA=2.5
B_PTL_B1|_TX|2 _PTL_B1|_TX|4 _PTL_B1|_TX|5 JJMIT AREA=2.5
I_PTL_B1|_TX|B1 0 _PTL_B1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B1|_TX|B2 0 _PTL_B1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|3  1.684e-12
L_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|6  3.596e-12
L_PTL_B1|_TX|1 B1 _PTL_B1|_TX|1  2.063e-12
L_PTL_B1|_TX|2 _PTL_B1|_TX|1 _PTL_B1|_TX|4  4.123e-12
L_PTL_B1|_TX|3 _PTL_B1|_TX|4 _PTL_B1|_TX|7  2.193e-12
R_PTL_B1|_TX|D _PTL_B1|_TX|7 _PTL_B1|A_PTL  1.36
L_PTL_B1|_TX|P1 _PTL_B1|_TX|2 0  5.254e-13
L_PTL_B1|_TX|P2 _PTL_B1|_TX|5 0  5.141e-13
R_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|101  2.7439617672
R_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|104  2.7439617672
L_PTL_B1|_TX|RB1 _PTL_B1|_TX|101 0  1.550338398468e-12
L_PTL_B1|_TX|RB2 _PTL_B1|_TX|104 0  1.550338398468e-12
B_PTL_B1|_RX|1 _PTL_B1|_RX|1 _PTL_B1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B1|_RX|2 _PTL_B1|_RX|4 _PTL_B1|_RX|5 JJMIT AREA=2.0
B_PTL_B1|_RX|3 _PTL_B1|_RX|7 _PTL_B1|_RX|8 JJMIT AREA=2.5
I_PTL_B1|_RX|B1 0 _PTL_B1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|3  2.777e-12
I_PTL_B1|_RX|B2 0 _PTL_B1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|6  2.685e-12
I_PTL_B1|_RX|B3 0 _PTL_B1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|9  2.764e-12
L_PTL_B1|_RX|1 _PTL_B1|A_PTL _PTL_B1|_RX|1  1.346e-12
L_PTL_B1|_RX|2 _PTL_B1|_RX|1 _PTL_B1|_RX|4  6.348e-12
L_PTL_B1|_RX|3 _PTL_B1|_RX|4 _PTL_B1|_RX|7  5.197e-12
L_PTL_B1|_RX|4 _PTL_B1|_RX|7 B1_RX  2.058e-12
L_PTL_B1|_RX|P1 _PTL_B1|_RX|2 0  4.795e-13
L_PTL_B1|_RX|P2 _PTL_B1|_RX|5 0  5.431e-13
L_PTL_B1|_RX|P3 _PTL_B1|_RX|8 0  5.339e-13
R_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|101  4.225701121488
R_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|104  3.429952209
R_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|107  2.7439617672
L_PTL_B1|_RX|RB1 _PTL_B1|_RX|101 0  2.38752113364072e-12
L_PTL_B1|_RX|RB2 _PTL_B1|_RX|104 0  1.937922998085e-12
L_PTL_B1|_RX|RB3 _PTL_B1|_RX|107 0  1.550338398468e-12
B_PTL_A2|_TX|1 _PTL_A2|_TX|1 _PTL_A2|_TX|2 JJMIT AREA=2.5
B_PTL_A2|_TX|2 _PTL_A2|_TX|4 _PTL_A2|_TX|5 JJMIT AREA=2.5
I_PTL_A2|_TX|B1 0 _PTL_A2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A2|_TX|B2 0 _PTL_A2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|3  1.684e-12
L_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|6  3.596e-12
L_PTL_A2|_TX|1 A2 _PTL_A2|_TX|1  2.063e-12
L_PTL_A2|_TX|2 _PTL_A2|_TX|1 _PTL_A2|_TX|4  4.123e-12
L_PTL_A2|_TX|3 _PTL_A2|_TX|4 _PTL_A2|_TX|7  2.193e-12
R_PTL_A2|_TX|D _PTL_A2|_TX|7 _PTL_A2|A_PTL  1.36
L_PTL_A2|_TX|P1 _PTL_A2|_TX|2 0  5.254e-13
L_PTL_A2|_TX|P2 _PTL_A2|_TX|5 0  5.141e-13
R_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|101  2.7439617672
R_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|104  2.7439617672
L_PTL_A2|_TX|RB1 _PTL_A2|_TX|101 0  1.550338398468e-12
L_PTL_A2|_TX|RB2 _PTL_A2|_TX|104 0  1.550338398468e-12
B_PTL_A2|_RX|1 _PTL_A2|_RX|1 _PTL_A2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A2|_RX|2 _PTL_A2|_RX|4 _PTL_A2|_RX|5 JJMIT AREA=2.0
B_PTL_A2|_RX|3 _PTL_A2|_RX|7 _PTL_A2|_RX|8 JJMIT AREA=2.5
I_PTL_A2|_RX|B1 0 _PTL_A2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|3  2.777e-12
I_PTL_A2|_RX|B2 0 _PTL_A2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|6  2.685e-12
I_PTL_A2|_RX|B3 0 _PTL_A2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|9  2.764e-12
L_PTL_A2|_RX|1 _PTL_A2|A_PTL _PTL_A2|_RX|1  1.346e-12
L_PTL_A2|_RX|2 _PTL_A2|_RX|1 _PTL_A2|_RX|4  6.348e-12
L_PTL_A2|_RX|3 _PTL_A2|_RX|4 _PTL_A2|_RX|7  5.197e-12
L_PTL_A2|_RX|4 _PTL_A2|_RX|7 A2_RX  2.058e-12
L_PTL_A2|_RX|P1 _PTL_A2|_RX|2 0  4.795e-13
L_PTL_A2|_RX|P2 _PTL_A2|_RX|5 0  5.431e-13
L_PTL_A2|_RX|P3 _PTL_A2|_RX|8 0  5.339e-13
R_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|101  4.225701121488
R_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|104  3.429952209
R_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|107  2.7439617672
L_PTL_A2|_RX|RB1 _PTL_A2|_RX|101 0  2.38752113364072e-12
L_PTL_A2|_RX|RB2 _PTL_A2|_RX|104 0  1.937922998085e-12
L_PTL_A2|_RX|RB3 _PTL_A2|_RX|107 0  1.550338398468e-12
B_PTL_B2|_TX|1 _PTL_B2|_TX|1 _PTL_B2|_TX|2 JJMIT AREA=2.5
B_PTL_B2|_TX|2 _PTL_B2|_TX|4 _PTL_B2|_TX|5 JJMIT AREA=2.5
I_PTL_B2|_TX|B1 0 _PTL_B2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B2|_TX|B2 0 _PTL_B2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|3  1.684e-12
L_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|6  3.596e-12
L_PTL_B2|_TX|1 B2 _PTL_B2|_TX|1  2.063e-12
L_PTL_B2|_TX|2 _PTL_B2|_TX|1 _PTL_B2|_TX|4  4.123e-12
L_PTL_B2|_TX|3 _PTL_B2|_TX|4 _PTL_B2|_TX|7  2.193e-12
R_PTL_B2|_TX|D _PTL_B2|_TX|7 _PTL_B2|A_PTL  1.36
L_PTL_B2|_TX|P1 _PTL_B2|_TX|2 0  5.254e-13
L_PTL_B2|_TX|P2 _PTL_B2|_TX|5 0  5.141e-13
R_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|101  2.7439617672
R_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|104  2.7439617672
L_PTL_B2|_TX|RB1 _PTL_B2|_TX|101 0  1.550338398468e-12
L_PTL_B2|_TX|RB2 _PTL_B2|_TX|104 0  1.550338398468e-12
B_PTL_B2|_RX|1 _PTL_B2|_RX|1 _PTL_B2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B2|_RX|2 _PTL_B2|_RX|4 _PTL_B2|_RX|5 JJMIT AREA=2.0
B_PTL_B2|_RX|3 _PTL_B2|_RX|7 _PTL_B2|_RX|8 JJMIT AREA=2.5
I_PTL_B2|_RX|B1 0 _PTL_B2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|3  2.777e-12
I_PTL_B2|_RX|B2 0 _PTL_B2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|6  2.685e-12
I_PTL_B2|_RX|B3 0 _PTL_B2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|9  2.764e-12
L_PTL_B2|_RX|1 _PTL_B2|A_PTL _PTL_B2|_RX|1  1.346e-12
L_PTL_B2|_RX|2 _PTL_B2|_RX|1 _PTL_B2|_RX|4  6.348e-12
L_PTL_B2|_RX|3 _PTL_B2|_RX|4 _PTL_B2|_RX|7  5.197e-12
L_PTL_B2|_RX|4 _PTL_B2|_RX|7 B2_RX  2.058e-12
L_PTL_B2|_RX|P1 _PTL_B2|_RX|2 0  4.795e-13
L_PTL_B2|_RX|P2 _PTL_B2|_RX|5 0  5.431e-13
L_PTL_B2|_RX|P3 _PTL_B2|_RX|8 0  5.339e-13
R_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|101  4.225701121488
R_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|104  3.429952209
R_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|107  2.7439617672
L_PTL_B2|_RX|RB1 _PTL_B2|_RX|101 0  2.38752113364072e-12
L_PTL_B2|_RX|RB2 _PTL_B2|_RX|104 0  1.937922998085e-12
L_PTL_B2|_RX|RB3 _PTL_B2|_RX|107 0  1.550338398468e-12
B_PTL_A3|_TX|1 _PTL_A3|_TX|1 _PTL_A3|_TX|2 JJMIT AREA=2.5
B_PTL_A3|_TX|2 _PTL_A3|_TX|4 _PTL_A3|_TX|5 JJMIT AREA=2.5
I_PTL_A3|_TX|B1 0 _PTL_A3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A3|_TX|B2 0 _PTL_A3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|3  1.684e-12
L_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|6  3.596e-12
L_PTL_A3|_TX|1 A3 _PTL_A3|_TX|1  2.063e-12
L_PTL_A3|_TX|2 _PTL_A3|_TX|1 _PTL_A3|_TX|4  4.123e-12
L_PTL_A3|_TX|3 _PTL_A3|_TX|4 _PTL_A3|_TX|7  2.193e-12
R_PTL_A3|_TX|D _PTL_A3|_TX|7 _PTL_A3|A_PTL  1.36
L_PTL_A3|_TX|P1 _PTL_A3|_TX|2 0  5.254e-13
L_PTL_A3|_TX|P2 _PTL_A3|_TX|5 0  5.141e-13
R_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|101  2.7439617672
R_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|104  2.7439617672
L_PTL_A3|_TX|RB1 _PTL_A3|_TX|101 0  1.550338398468e-12
L_PTL_A3|_TX|RB2 _PTL_A3|_TX|104 0  1.550338398468e-12
B_PTL_A3|_RX|1 _PTL_A3|_RX|1 _PTL_A3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A3|_RX|2 _PTL_A3|_RX|4 _PTL_A3|_RX|5 JJMIT AREA=2.0
B_PTL_A3|_RX|3 _PTL_A3|_RX|7 _PTL_A3|_RX|8 JJMIT AREA=2.5
I_PTL_A3|_RX|B1 0 _PTL_A3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|3  2.777e-12
I_PTL_A3|_RX|B2 0 _PTL_A3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|6  2.685e-12
I_PTL_A3|_RX|B3 0 _PTL_A3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|9  2.764e-12
L_PTL_A3|_RX|1 _PTL_A3|A_PTL _PTL_A3|_RX|1  1.346e-12
L_PTL_A3|_RX|2 _PTL_A3|_RX|1 _PTL_A3|_RX|4  6.348e-12
L_PTL_A3|_RX|3 _PTL_A3|_RX|4 _PTL_A3|_RX|7  5.197e-12
L_PTL_A3|_RX|4 _PTL_A3|_RX|7 A3_RX  2.058e-12
L_PTL_A3|_RX|P1 _PTL_A3|_RX|2 0  4.795e-13
L_PTL_A3|_RX|P2 _PTL_A3|_RX|5 0  5.431e-13
L_PTL_A3|_RX|P3 _PTL_A3|_RX|8 0  5.339e-13
R_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|101  4.225701121488
R_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|104  3.429952209
R_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|107  2.7439617672
L_PTL_A3|_RX|RB1 _PTL_A3|_RX|101 0  2.38752113364072e-12
L_PTL_A3|_RX|RB2 _PTL_A3|_RX|104 0  1.937922998085e-12
L_PTL_A3|_RX|RB3 _PTL_A3|_RX|107 0  1.550338398468e-12
B_PTL_B3|_TX|1 _PTL_B3|_TX|1 _PTL_B3|_TX|2 JJMIT AREA=2.5
B_PTL_B3|_TX|2 _PTL_B3|_TX|4 _PTL_B3|_TX|5 JJMIT AREA=2.5
I_PTL_B3|_TX|B1 0 _PTL_B3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B3|_TX|B2 0 _PTL_B3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|3  1.684e-12
L_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|6  3.596e-12
L_PTL_B3|_TX|1 B3 _PTL_B3|_TX|1  2.063e-12
L_PTL_B3|_TX|2 _PTL_B3|_TX|1 _PTL_B3|_TX|4  4.123e-12
L_PTL_B3|_TX|3 _PTL_B3|_TX|4 _PTL_B3|_TX|7  2.193e-12
R_PTL_B3|_TX|D _PTL_B3|_TX|7 _PTL_B3|A_PTL  1.36
L_PTL_B3|_TX|P1 _PTL_B3|_TX|2 0  5.254e-13
L_PTL_B3|_TX|P2 _PTL_B3|_TX|5 0  5.141e-13
R_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|101  2.7439617672
R_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|104  2.7439617672
L_PTL_B3|_TX|RB1 _PTL_B3|_TX|101 0  1.550338398468e-12
L_PTL_B3|_TX|RB2 _PTL_B3|_TX|104 0  1.550338398468e-12
B_PTL_B3|_RX|1 _PTL_B3|_RX|1 _PTL_B3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B3|_RX|2 _PTL_B3|_RX|4 _PTL_B3|_RX|5 JJMIT AREA=2.0
B_PTL_B3|_RX|3 _PTL_B3|_RX|7 _PTL_B3|_RX|8 JJMIT AREA=2.5
I_PTL_B3|_RX|B1 0 _PTL_B3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|3  2.777e-12
I_PTL_B3|_RX|B2 0 _PTL_B3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|6  2.685e-12
I_PTL_B3|_RX|B3 0 _PTL_B3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|9  2.764e-12
L_PTL_B3|_RX|1 _PTL_B3|A_PTL _PTL_B3|_RX|1  1.346e-12
L_PTL_B3|_RX|2 _PTL_B3|_RX|1 _PTL_B3|_RX|4  6.348e-12
L_PTL_B3|_RX|3 _PTL_B3|_RX|4 _PTL_B3|_RX|7  5.197e-12
L_PTL_B3|_RX|4 _PTL_B3|_RX|7 B3_RX  2.058e-12
L_PTL_B3|_RX|P1 _PTL_B3|_RX|2 0  4.795e-13
L_PTL_B3|_RX|P2 _PTL_B3|_RX|5 0  5.431e-13
L_PTL_B3|_RX|P3 _PTL_B3|_RX|8 0  5.339e-13
R_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|101  4.225701121488
R_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|104  3.429952209
R_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|107  2.7439617672
L_PTL_B3|_RX|RB1 _PTL_B3|_RX|101 0  2.38752113364072e-12
L_PTL_B3|_RX|RB2 _PTL_B3|_RX|104 0  1.937922998085e-12
L_PTL_B3|_RX|RB3 _PTL_B3|_RX|107 0  1.550338398468e-12
LI0|_SPL_A|1 A0_RX I0|_SPL_A|D1  2e-12
LI0|_SPL_A|2 I0|_SPL_A|D1 I0|_SPL_A|D2  4.135667696e-12
LI0|_SPL_A|3 I0|_SPL_A|D2 I0|_SPL_A|JCT  9.84682784761905e-13
LI0|_SPL_A|4 I0|_SPL_A|JCT I0|_SPL_A|QA1  9.84682784761905e-13
LI0|_SPL_A|5 I0|_SPL_A|QA1 I0|A1  2e-12
LI0|_SPL_A|6 I0|_SPL_A|JCT I0|_SPL_A|QB1  9.84682784761905e-13
LI0|_SPL_A|7 I0|_SPL_A|QB1 I0|A2  2e-12
LI0|_SPL_B|1 B0_RX I0|_SPL_B|D1  2e-12
LI0|_SPL_B|2 I0|_SPL_B|D1 I0|_SPL_B|D2  4.135667696e-12
LI0|_SPL_B|3 I0|_SPL_B|D2 I0|_SPL_B|JCT  9.84682784761905e-13
LI0|_SPL_B|4 I0|_SPL_B|JCT I0|_SPL_B|QA1  9.84682784761905e-13
LI0|_SPL_B|5 I0|_SPL_B|QA1 I0|B1  2e-12
LI0|_SPL_B|6 I0|_SPL_B|JCT I0|_SPL_B|QB1  9.84682784761905e-13
LI0|_SPL_B|7 I0|_SPL_B|QB1 I0|B2  2e-12
LI0|_DFF_A|1 I0|A1 I0|_DFF_A|A1  2.067833848e-12
LI0|_DFF_A|2 I0|_DFF_A|A1 I0|_DFF_A|A2  4.135667696e-12
LI0|_DFF_A|3 I0|_DFF_A|A3 I0|_DFF_A|A4  8.271335392e-12
LI0|_DFF_A|T T00 I0|_DFF_A|T1  2.067833848e-12
LI0|_DFF_A|4 I0|_DFF_A|T1 I0|_DFF_A|T2  4.135667696e-12
LI0|_DFF_A|5 I0|_DFF_A|A4 I0|_DFF_A|Q1  4.135667696e-12
LI0|_DFF_A|6 I0|_DFF_A|Q1 I0|A1_SYNC  2.067833848e-12
LI0|_DFF_B|1 I0|B1 I0|_DFF_B|A1  2.067833848e-12
LI0|_DFF_B|2 I0|_DFF_B|A1 I0|_DFF_B|A2  4.135667696e-12
LI0|_DFF_B|3 I0|_DFF_B|A3 I0|_DFF_B|A4  8.271335392e-12
LI0|_DFF_B|T T00 I0|_DFF_B|T1  2.067833848e-12
LI0|_DFF_B|4 I0|_DFF_B|T1 I0|_DFF_B|T2  4.135667696e-12
LI0|_DFF_B|5 I0|_DFF_B|A4 I0|_DFF_B|Q1  4.135667696e-12
LI0|_DFF_B|6 I0|_DFF_B|Q1 I0|B1_SYNC  2.067833848e-12
LI0|_XOR|A1 I0|A2 I0|_XOR|A1  2.067833848e-12
LI0|_XOR|A2 I0|_XOR|A1 I0|_XOR|A2  4.135667696e-12
LI0|_XOR|A3 I0|_XOR|A3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|B1 I0|B2 I0|_XOR|B1  2.067833848e-12
LI0|_XOR|B2 I0|_XOR|B1 I0|_XOR|B2  4.135667696e-12
LI0|_XOR|B3 I0|_XOR|B3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|T1 T00 I0|_XOR|T1  2.067833848e-12
LI0|_XOR|T2 I0|_XOR|T1 I0|_XOR|T2  4.135667696e-12
LI0|_XOR|Q2 I0|_XOR|ABTQ I0|_XOR|Q1  4.135667696e-12
LI0|_XOR|Q1 I0|_XOR|Q1 IP0_0  2.067833848e-12
LI0|_AND|A1 I0|A1_SYNC I0|_AND|A1  2.067833848e-12
LI0|_AND|A2 I0|_AND|A1 I0|_AND|A2  4.135667696e-12
LI0|_AND|A3 I0|_AND|A3 I0|_AND|Q3  1.2e-12
LI0|_AND|B1 I0|B1_SYNC I0|_AND|B1  2.067833848e-12
LI0|_AND|B2 I0|_AND|B1 I0|_AND|B2  4.135667696e-12
LI0|_AND|B3 I0|_AND|B3 I0|_AND|Q3  1.2e-12
LI0|_AND|Q3 I0|_AND|Q3 I0|_AND|Q2  4.135667696e-12
LI0|_AND|Q2 I0|_AND|Q2 I0|_AND|Q1  4.135667696e-12
LI0|_AND|Q1 I0|_AND|Q1 IG0_0  2.067833848e-12
LI1|_SPL_A|1 A1_RX I1|_SPL_A|D1  2e-12
LI1|_SPL_A|2 I1|_SPL_A|D1 I1|_SPL_A|D2  4.135667696e-12
LI1|_SPL_A|3 I1|_SPL_A|D2 I1|_SPL_A|JCT  9.84682784761905e-13
LI1|_SPL_A|4 I1|_SPL_A|JCT I1|_SPL_A|QA1  9.84682784761905e-13
LI1|_SPL_A|5 I1|_SPL_A|QA1 I1|A1  2e-12
LI1|_SPL_A|6 I1|_SPL_A|JCT I1|_SPL_A|QB1  9.84682784761905e-13
LI1|_SPL_A|7 I1|_SPL_A|QB1 I1|A2  2e-12
LI1|_SPL_B|1 B1_RX I1|_SPL_B|D1  2e-12
LI1|_SPL_B|2 I1|_SPL_B|D1 I1|_SPL_B|D2  4.135667696e-12
LI1|_SPL_B|3 I1|_SPL_B|D2 I1|_SPL_B|JCT  9.84682784761905e-13
LI1|_SPL_B|4 I1|_SPL_B|JCT I1|_SPL_B|QA1  9.84682784761905e-13
LI1|_SPL_B|5 I1|_SPL_B|QA1 I1|B1  2e-12
LI1|_SPL_B|6 I1|_SPL_B|JCT I1|_SPL_B|QB1  9.84682784761905e-13
LI1|_SPL_B|7 I1|_SPL_B|QB1 I1|B2  2e-12
LI1|_DFF_A|1 I1|A1 I1|_DFF_A|A1  2.067833848e-12
LI1|_DFF_A|2 I1|_DFF_A|A1 I1|_DFF_A|A2  4.135667696e-12
LI1|_DFF_A|3 I1|_DFF_A|A3 I1|_DFF_A|A4  8.271335392e-12
LI1|_DFF_A|T T01 I1|_DFF_A|T1  2.067833848e-12
LI1|_DFF_A|4 I1|_DFF_A|T1 I1|_DFF_A|T2  4.135667696e-12
LI1|_DFF_A|5 I1|_DFF_A|A4 I1|_DFF_A|Q1  4.135667696e-12
LI1|_DFF_A|6 I1|_DFF_A|Q1 I1|A1_SYNC  2.067833848e-12
LI1|_DFF_B|1 I1|B1 I1|_DFF_B|A1  2.067833848e-12
LI1|_DFF_B|2 I1|_DFF_B|A1 I1|_DFF_B|A2  4.135667696e-12
LI1|_DFF_B|3 I1|_DFF_B|A3 I1|_DFF_B|A4  8.271335392e-12
LI1|_DFF_B|T T01 I1|_DFF_B|T1  2.067833848e-12
LI1|_DFF_B|4 I1|_DFF_B|T1 I1|_DFF_B|T2  4.135667696e-12
LI1|_DFF_B|5 I1|_DFF_B|A4 I1|_DFF_B|Q1  4.135667696e-12
LI1|_DFF_B|6 I1|_DFF_B|Q1 I1|B1_SYNC  2.067833848e-12
LI1|_XOR|A1 I1|A2 I1|_XOR|A1  2.067833848e-12
LI1|_XOR|A2 I1|_XOR|A1 I1|_XOR|A2  4.135667696e-12
LI1|_XOR|A3 I1|_XOR|A3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|B1 I1|B2 I1|_XOR|B1  2.067833848e-12
LI1|_XOR|B2 I1|_XOR|B1 I1|_XOR|B2  4.135667696e-12
LI1|_XOR|B3 I1|_XOR|B3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|T1 T01 I1|_XOR|T1  2.067833848e-12
LI1|_XOR|T2 I1|_XOR|T1 I1|_XOR|T2  4.135667696e-12
LI1|_XOR|Q2 I1|_XOR|ABTQ I1|_XOR|Q1  4.135667696e-12
LI1|_XOR|Q1 I1|_XOR|Q1 IP1_0  2.067833848e-12
LI1|_AND|A1 I1|A1_SYNC I1|_AND|A1  2.067833848e-12
LI1|_AND|A2 I1|_AND|A1 I1|_AND|A2  4.135667696e-12
LI1|_AND|A3 I1|_AND|A3 I1|_AND|Q3  1.2e-12
LI1|_AND|B1 I1|B1_SYNC I1|_AND|B1  2.067833848e-12
LI1|_AND|B2 I1|_AND|B1 I1|_AND|B2  4.135667696e-12
LI1|_AND|B3 I1|_AND|B3 I1|_AND|Q3  1.2e-12
LI1|_AND|Q3 I1|_AND|Q3 I1|_AND|Q2  4.135667696e-12
LI1|_AND|Q2 I1|_AND|Q2 I1|_AND|Q1  4.135667696e-12
LI1|_AND|Q1 I1|_AND|Q1 IG1_0  2.067833848e-12
LI2|_SPL_A|1 A2_RX I2|_SPL_A|D1  2e-12
LI2|_SPL_A|2 I2|_SPL_A|D1 I2|_SPL_A|D2  4.135667696e-12
LI2|_SPL_A|3 I2|_SPL_A|D2 I2|_SPL_A|JCT  9.84682784761905e-13
LI2|_SPL_A|4 I2|_SPL_A|JCT I2|_SPL_A|QA1  9.84682784761905e-13
LI2|_SPL_A|5 I2|_SPL_A|QA1 I2|A1  2e-12
LI2|_SPL_A|6 I2|_SPL_A|JCT I2|_SPL_A|QB1  9.84682784761905e-13
LI2|_SPL_A|7 I2|_SPL_A|QB1 I2|A2  2e-12
LI2|_SPL_B|1 B2_RX I2|_SPL_B|D1  2e-12
LI2|_SPL_B|2 I2|_SPL_B|D1 I2|_SPL_B|D2  4.135667696e-12
LI2|_SPL_B|3 I2|_SPL_B|D2 I2|_SPL_B|JCT  9.84682784761905e-13
LI2|_SPL_B|4 I2|_SPL_B|JCT I2|_SPL_B|QA1  9.84682784761905e-13
LI2|_SPL_B|5 I2|_SPL_B|QA1 I2|B1  2e-12
LI2|_SPL_B|6 I2|_SPL_B|JCT I2|_SPL_B|QB1  9.84682784761905e-13
LI2|_SPL_B|7 I2|_SPL_B|QB1 I2|B2  2e-12
LI2|_DFF_A|1 I2|A1 I2|_DFF_A|A1  2.067833848e-12
LI2|_DFF_A|2 I2|_DFF_A|A1 I2|_DFF_A|A2  4.135667696e-12
LI2|_DFF_A|3 I2|_DFF_A|A3 I2|_DFF_A|A4  8.271335392e-12
LI2|_DFF_A|T T02 I2|_DFF_A|T1  2.067833848e-12
LI2|_DFF_A|4 I2|_DFF_A|T1 I2|_DFF_A|T2  4.135667696e-12
LI2|_DFF_A|5 I2|_DFF_A|A4 I2|_DFF_A|Q1  4.135667696e-12
LI2|_DFF_A|6 I2|_DFF_A|Q1 I2|A1_SYNC  2.067833848e-12
LI2|_DFF_B|1 I2|B1 I2|_DFF_B|A1  2.067833848e-12
LI2|_DFF_B|2 I2|_DFF_B|A1 I2|_DFF_B|A2  4.135667696e-12
LI2|_DFF_B|3 I2|_DFF_B|A3 I2|_DFF_B|A4  8.271335392e-12
LI2|_DFF_B|T T02 I2|_DFF_B|T1  2.067833848e-12
LI2|_DFF_B|4 I2|_DFF_B|T1 I2|_DFF_B|T2  4.135667696e-12
LI2|_DFF_B|5 I2|_DFF_B|A4 I2|_DFF_B|Q1  4.135667696e-12
LI2|_DFF_B|6 I2|_DFF_B|Q1 I2|B1_SYNC  2.067833848e-12
LI2|_XOR|A1 I2|A2 I2|_XOR|A1  2.067833848e-12
LI2|_XOR|A2 I2|_XOR|A1 I2|_XOR|A2  4.135667696e-12
LI2|_XOR|A3 I2|_XOR|A3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|B1 I2|B2 I2|_XOR|B1  2.067833848e-12
LI2|_XOR|B2 I2|_XOR|B1 I2|_XOR|B2  4.135667696e-12
LI2|_XOR|B3 I2|_XOR|B3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|T1 T02 I2|_XOR|T1  2.067833848e-12
LI2|_XOR|T2 I2|_XOR|T1 I2|_XOR|T2  4.135667696e-12
LI2|_XOR|Q2 I2|_XOR|ABTQ I2|_XOR|Q1  4.135667696e-12
LI2|_XOR|Q1 I2|_XOR|Q1 IP2_0  2.067833848e-12
LI2|_AND|A1 I2|A1_SYNC I2|_AND|A1  2.067833848e-12
LI2|_AND|A2 I2|_AND|A1 I2|_AND|A2  4.135667696e-12
LI2|_AND|A3 I2|_AND|A3 I2|_AND|Q3  1.2e-12
LI2|_AND|B1 I2|B1_SYNC I2|_AND|B1  2.067833848e-12
LI2|_AND|B2 I2|_AND|B1 I2|_AND|B2  4.135667696e-12
LI2|_AND|B3 I2|_AND|B3 I2|_AND|Q3  1.2e-12
LI2|_AND|Q3 I2|_AND|Q3 I2|_AND|Q2  4.135667696e-12
LI2|_AND|Q2 I2|_AND|Q2 I2|_AND|Q1  4.135667696e-12
LI2|_AND|Q1 I2|_AND|Q1 IG2_0  2.067833848e-12
LI3|_SPL_A|1 A3_RX I3|_SPL_A|D1  2e-12
LI3|_SPL_A|2 I3|_SPL_A|D1 I3|_SPL_A|D2  4.135667696e-12
LI3|_SPL_A|3 I3|_SPL_A|D2 I3|_SPL_A|JCT  9.84682784761905e-13
LI3|_SPL_A|4 I3|_SPL_A|JCT I3|_SPL_A|QA1  9.84682784761905e-13
LI3|_SPL_A|5 I3|_SPL_A|QA1 I3|A1  2e-12
LI3|_SPL_A|6 I3|_SPL_A|JCT I3|_SPL_A|QB1  9.84682784761905e-13
LI3|_SPL_A|7 I3|_SPL_A|QB1 I3|A2  2e-12
LI3|_SPL_B|1 B3_RX I3|_SPL_B|D1  2e-12
LI3|_SPL_B|2 I3|_SPL_B|D1 I3|_SPL_B|D2  4.135667696e-12
LI3|_SPL_B|3 I3|_SPL_B|D2 I3|_SPL_B|JCT  9.84682784761905e-13
LI3|_SPL_B|4 I3|_SPL_B|JCT I3|_SPL_B|QA1  9.84682784761905e-13
LI3|_SPL_B|5 I3|_SPL_B|QA1 I3|B1  2e-12
LI3|_SPL_B|6 I3|_SPL_B|JCT I3|_SPL_B|QB1  9.84682784761905e-13
LI3|_SPL_B|7 I3|_SPL_B|QB1 I3|B2  2e-12
LI3|_DFF_A|1 I3|A1 I3|_DFF_A|A1  2.067833848e-12
LI3|_DFF_A|2 I3|_DFF_A|A1 I3|_DFF_A|A2  4.135667696e-12
LI3|_DFF_A|3 I3|_DFF_A|A3 I3|_DFF_A|A4  8.271335392e-12
LI3|_DFF_A|T T03 I3|_DFF_A|T1  2.067833848e-12
LI3|_DFF_A|4 I3|_DFF_A|T1 I3|_DFF_A|T2  4.135667696e-12
LI3|_DFF_A|5 I3|_DFF_A|A4 I3|_DFF_A|Q1  4.135667696e-12
LI3|_DFF_A|6 I3|_DFF_A|Q1 I3|A1_SYNC  2.067833848e-12
LI3|_DFF_B|1 I3|B1 I3|_DFF_B|A1  2.067833848e-12
LI3|_DFF_B|2 I3|_DFF_B|A1 I3|_DFF_B|A2  4.135667696e-12
LI3|_DFF_B|3 I3|_DFF_B|A3 I3|_DFF_B|A4  8.271335392e-12
LI3|_DFF_B|T T03 I3|_DFF_B|T1  2.067833848e-12
LI3|_DFF_B|4 I3|_DFF_B|T1 I3|_DFF_B|T2  4.135667696e-12
LI3|_DFF_B|5 I3|_DFF_B|A4 I3|_DFF_B|Q1  4.135667696e-12
LI3|_DFF_B|6 I3|_DFF_B|Q1 I3|B1_SYNC  2.067833848e-12
LI3|_XOR|A1 I3|A2 I3|_XOR|A1  2.067833848e-12
LI3|_XOR|A2 I3|_XOR|A1 I3|_XOR|A2  4.135667696e-12
LI3|_XOR|A3 I3|_XOR|A3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|B1 I3|B2 I3|_XOR|B1  2.067833848e-12
LI3|_XOR|B2 I3|_XOR|B1 I3|_XOR|B2  4.135667696e-12
LI3|_XOR|B3 I3|_XOR|B3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|T1 T03 I3|_XOR|T1  2.067833848e-12
LI3|_XOR|T2 I3|_XOR|T1 I3|_XOR|T2  4.135667696e-12
LI3|_XOR|Q2 I3|_XOR|ABTQ I3|_XOR|Q1  4.135667696e-12
LI3|_XOR|Q1 I3|_XOR|Q1 IP3_0  2.067833848e-12
LI3|_AND|A1 I3|A1_SYNC I3|_AND|A1  2.067833848e-12
LI3|_AND|A2 I3|_AND|A1 I3|_AND|A2  4.135667696e-12
LI3|_AND|A3 I3|_AND|A3 I3|_AND|Q3  1.2e-12
LI3|_AND|B1 I3|B1_SYNC I3|_AND|B1  2.067833848e-12
LI3|_AND|B2 I3|_AND|B1 I3|_AND|B2  4.135667696e-12
LI3|_AND|B3 I3|_AND|B3 I3|_AND|Q3  1.2e-12
LI3|_AND|Q3 I3|_AND|Q3 I3|_AND|Q2  4.135667696e-12
LI3|_AND|Q2 I3|_AND|Q2 I3|_AND|Q1  4.135667696e-12
LI3|_AND|Q1 I3|_AND|Q1 IG3_0  2.067833848e-12
B_PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP0_0|_TX|B1 0 _PTL_IP0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP0_0|_TX|B2 0 _PTL_IP0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|3  1.684e-12
L_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|6  3.596e-12
L_PTL_IP0_0|_TX|1 IP0_0 _PTL_IP0_0|_TX|1  2.063e-12
L_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|4  4.123e-12
L_PTL_IP0_0|_TX|3 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|7  2.193e-12
R_PTL_IP0_0|_TX|D _PTL_IP0_0|_TX|7 _PTL_IP0_0|A_PTL  1.36
L_PTL_IP0_0|_TX|P1 _PTL_IP0_0|_TX|2 0  5.254e-13
L_PTL_IP0_0|_TX|P2 _PTL_IP0_0|_TX|5 0  5.141e-13
R_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|101  2.7439617672
R_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|104  2.7439617672
L_PTL_IP0_0|_TX|RB1 _PTL_IP0_0|_TX|101 0  1.550338398468e-12
L_PTL_IP0_0|_TX|RB2 _PTL_IP0_0|_TX|104 0  1.550338398468e-12
B_PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP0_0|_RX|B1 0 _PTL_IP0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|3  2.777e-12
I_PTL_IP0_0|_RX|B2 0 _PTL_IP0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|6  2.685e-12
I_PTL_IP0_0|_RX|B3 0 _PTL_IP0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|9  2.764e-12
L_PTL_IP0_0|_RX|1 _PTL_IP0_0|A_PTL _PTL_IP0_0|_RX|1  1.346e-12
L_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|4  6.348e-12
L_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7  5.197e-12
L_PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7 IP0_0_RX  2.058e-12
L_PTL_IP0_0|_RX|P1 _PTL_IP0_0|_RX|2 0  4.795e-13
L_PTL_IP0_0|_RX|P2 _PTL_IP0_0|_RX|5 0  5.431e-13
L_PTL_IP0_0|_RX|P3 _PTL_IP0_0|_RX|8 0  5.339e-13
R_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|101  4.225701121488
R_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|104  3.429952209
R_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|107  2.7439617672
L_PTL_IP0_0|_RX|RB1 _PTL_IP0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP0_0|_RX|RB2 _PTL_IP0_0|_RX|104 0  1.937922998085e-12
L_PTL_IP0_0|_RX|RB3 _PTL_IP0_0|_RX|107 0  1.550338398468e-12
B_PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG0_0|_TX|B1 0 _PTL_IG0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG0_0|_TX|B2 0 _PTL_IG0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|3  1.684e-12
L_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|6  3.596e-12
L_PTL_IG0_0|_TX|1 IG0_0 _PTL_IG0_0|_TX|1  2.063e-12
L_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|4  4.123e-12
L_PTL_IG0_0|_TX|3 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|7  2.193e-12
R_PTL_IG0_0|_TX|D _PTL_IG0_0|_TX|7 _PTL_IG0_0|A_PTL  1.36
L_PTL_IG0_0|_TX|P1 _PTL_IG0_0|_TX|2 0  5.254e-13
L_PTL_IG0_0|_TX|P2 _PTL_IG0_0|_TX|5 0  5.141e-13
R_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|101  2.7439617672
R_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|104  2.7439617672
L_PTL_IG0_0|_TX|RB1 _PTL_IG0_0|_TX|101 0  1.550338398468e-12
L_PTL_IG0_0|_TX|RB2 _PTL_IG0_0|_TX|104 0  1.550338398468e-12
B_PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG0_0|_RX|B1 0 _PTL_IG0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|3  2.777e-12
I_PTL_IG0_0|_RX|B2 0 _PTL_IG0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|6  2.685e-12
I_PTL_IG0_0|_RX|B3 0 _PTL_IG0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|9  2.764e-12
L_PTL_IG0_0|_RX|1 _PTL_IG0_0|A_PTL _PTL_IG0_0|_RX|1  1.346e-12
L_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|4  6.348e-12
L_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7  5.197e-12
L_PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7 IG0_0_RX  2.058e-12
L_PTL_IG0_0|_RX|P1 _PTL_IG0_0|_RX|2 0  4.795e-13
L_PTL_IG0_0|_RX|P2 _PTL_IG0_0|_RX|5 0  5.431e-13
L_PTL_IG0_0|_RX|P3 _PTL_IG0_0|_RX|8 0  5.339e-13
R_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|101  4.225701121488
R_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|104  3.429952209
R_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|107  2.7439617672
L_PTL_IG0_0|_RX|RB1 _PTL_IG0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG0_0|_RX|RB2 _PTL_IG0_0|_RX|104 0  1.937922998085e-12
L_PTL_IG0_0|_RX|RB3 _PTL_IG0_0|_RX|107 0  1.550338398468e-12
B_PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_0|_TX|B1 0 _PTL_IP1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_0|_TX|B2 0 _PTL_IP1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|3  1.684e-12
L_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|6  3.596e-12
L_PTL_IP1_0|_TX|1 IP1_0 _PTL_IP1_0|_TX|1  2.063e-12
L_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|4  4.123e-12
L_PTL_IP1_0|_TX|3 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|7  2.193e-12
R_PTL_IP1_0|_TX|D _PTL_IP1_0|_TX|7 _PTL_IP1_0|A_PTL  1.36
L_PTL_IP1_0|_TX|P1 _PTL_IP1_0|_TX|2 0  5.254e-13
L_PTL_IP1_0|_TX|P2 _PTL_IP1_0|_TX|5 0  5.141e-13
R_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|101  2.7439617672
R_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|104  2.7439617672
L_PTL_IP1_0|_TX|RB1 _PTL_IP1_0|_TX|101 0  1.550338398468e-12
L_PTL_IP1_0|_TX|RB2 _PTL_IP1_0|_TX|104 0  1.550338398468e-12
B_PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_0|_RX|B1 0 _PTL_IP1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|3  2.777e-12
I_PTL_IP1_0|_RX|B2 0 _PTL_IP1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|6  2.685e-12
I_PTL_IP1_0|_RX|B3 0 _PTL_IP1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|9  2.764e-12
L_PTL_IP1_0|_RX|1 _PTL_IP1_0|A_PTL _PTL_IP1_0|_RX|1  1.346e-12
L_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|4  6.348e-12
L_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7  5.197e-12
L_PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7 IP1_0_RX  2.058e-12
L_PTL_IP1_0|_RX|P1 _PTL_IP1_0|_RX|2 0  4.795e-13
L_PTL_IP1_0|_RX|P2 _PTL_IP1_0|_RX|5 0  5.431e-13
L_PTL_IP1_0|_RX|P3 _PTL_IP1_0|_RX|8 0  5.339e-13
R_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|101  4.225701121488
R_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|104  3.429952209
R_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|107  2.7439617672
L_PTL_IP1_0|_RX|RB1 _PTL_IP1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_0|_RX|RB2 _PTL_IP1_0|_RX|104 0  1.937922998085e-12
L_PTL_IP1_0|_RX|RB3 _PTL_IP1_0|_RX|107 0  1.550338398468e-12
B_PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG1_0|_TX|B1 0 _PTL_IG1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG1_0|_TX|B2 0 _PTL_IG1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|3  1.684e-12
L_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|6  3.596e-12
L_PTL_IG1_0|_TX|1 IG1_0 _PTL_IG1_0|_TX|1  2.063e-12
L_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|4  4.123e-12
L_PTL_IG1_0|_TX|3 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|7  2.193e-12
R_PTL_IG1_0|_TX|D _PTL_IG1_0|_TX|7 _PTL_IG1_0|A_PTL  1.36
L_PTL_IG1_0|_TX|P1 _PTL_IG1_0|_TX|2 0  5.254e-13
L_PTL_IG1_0|_TX|P2 _PTL_IG1_0|_TX|5 0  5.141e-13
R_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|101  2.7439617672
R_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|104  2.7439617672
L_PTL_IG1_0|_TX|RB1 _PTL_IG1_0|_TX|101 0  1.550338398468e-12
L_PTL_IG1_0|_TX|RB2 _PTL_IG1_0|_TX|104 0  1.550338398468e-12
B_PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG1_0|_RX|B1 0 _PTL_IG1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|3  2.777e-12
I_PTL_IG1_0|_RX|B2 0 _PTL_IG1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|6  2.685e-12
I_PTL_IG1_0|_RX|B3 0 _PTL_IG1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|9  2.764e-12
L_PTL_IG1_0|_RX|1 _PTL_IG1_0|A_PTL _PTL_IG1_0|_RX|1  1.346e-12
L_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|4  6.348e-12
L_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7  5.197e-12
L_PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7 IG1_0_RX  2.058e-12
L_PTL_IG1_0|_RX|P1 _PTL_IG1_0|_RX|2 0  4.795e-13
L_PTL_IG1_0|_RX|P2 _PTL_IG1_0|_RX|5 0  5.431e-13
L_PTL_IG1_0|_RX|P3 _PTL_IG1_0|_RX|8 0  5.339e-13
R_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|101  4.225701121488
R_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|104  3.429952209
R_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|107  2.7439617672
L_PTL_IG1_0|_RX|RB1 _PTL_IG1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG1_0|_RX|RB2 _PTL_IG1_0|_RX|104 0  1.937922998085e-12
L_PTL_IG1_0|_RX|RB3 _PTL_IG1_0|_RX|107 0  1.550338398468e-12
B_PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_0|_TX|B1 0 _PTL_IP2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_0|_TX|B2 0 _PTL_IP2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|3  1.684e-12
L_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|6  3.596e-12
L_PTL_IP2_0|_TX|1 IP2_0 _PTL_IP2_0|_TX|1  2.063e-12
L_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|4  4.123e-12
L_PTL_IP2_0|_TX|3 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|7  2.193e-12
R_PTL_IP2_0|_TX|D _PTL_IP2_0|_TX|7 _PTL_IP2_0|A_PTL  1.36
L_PTL_IP2_0|_TX|P1 _PTL_IP2_0|_TX|2 0  5.254e-13
L_PTL_IP2_0|_TX|P2 _PTL_IP2_0|_TX|5 0  5.141e-13
R_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|101  2.7439617672
R_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|104  2.7439617672
L_PTL_IP2_0|_TX|RB1 _PTL_IP2_0|_TX|101 0  1.550338398468e-12
L_PTL_IP2_0|_TX|RB2 _PTL_IP2_0|_TX|104 0  1.550338398468e-12
B_PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_0|_RX|B1 0 _PTL_IP2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|3  2.777e-12
I_PTL_IP2_0|_RX|B2 0 _PTL_IP2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|6  2.685e-12
I_PTL_IP2_0|_RX|B3 0 _PTL_IP2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|9  2.764e-12
L_PTL_IP2_0|_RX|1 _PTL_IP2_0|A_PTL _PTL_IP2_0|_RX|1  1.346e-12
L_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|4  6.348e-12
L_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7  5.197e-12
L_PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7 IP2_0_RX  2.058e-12
L_PTL_IP2_0|_RX|P1 _PTL_IP2_0|_RX|2 0  4.795e-13
L_PTL_IP2_0|_RX|P2 _PTL_IP2_0|_RX|5 0  5.431e-13
L_PTL_IP2_0|_RX|P3 _PTL_IP2_0|_RX|8 0  5.339e-13
R_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|101  4.225701121488
R_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|104  3.429952209
R_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|107  2.7439617672
L_PTL_IP2_0|_RX|RB1 _PTL_IP2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_0|_RX|RB2 _PTL_IP2_0|_RX|104 0  1.937922998085e-12
L_PTL_IP2_0|_RX|RB3 _PTL_IP2_0|_RX|107 0  1.550338398468e-12
B_PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG2_0|_TX|B1 0 _PTL_IG2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG2_0|_TX|B2 0 _PTL_IG2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|3  1.684e-12
L_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|6  3.596e-12
L_PTL_IG2_0|_TX|1 IG2_0 _PTL_IG2_0|_TX|1  2.063e-12
L_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|4  4.123e-12
L_PTL_IG2_0|_TX|3 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|7  2.193e-12
R_PTL_IG2_0|_TX|D _PTL_IG2_0|_TX|7 _PTL_IG2_0|A_PTL  1.36
L_PTL_IG2_0|_TX|P1 _PTL_IG2_0|_TX|2 0  5.254e-13
L_PTL_IG2_0|_TX|P2 _PTL_IG2_0|_TX|5 0  5.141e-13
R_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|101  2.7439617672
R_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|104  2.7439617672
L_PTL_IG2_0|_TX|RB1 _PTL_IG2_0|_TX|101 0  1.550338398468e-12
L_PTL_IG2_0|_TX|RB2 _PTL_IG2_0|_TX|104 0  1.550338398468e-12
B_PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG2_0|_RX|B1 0 _PTL_IG2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|3  2.777e-12
I_PTL_IG2_0|_RX|B2 0 _PTL_IG2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|6  2.685e-12
I_PTL_IG2_0|_RX|B3 0 _PTL_IG2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|9  2.764e-12
L_PTL_IG2_0|_RX|1 _PTL_IG2_0|A_PTL _PTL_IG2_0|_RX|1  1.346e-12
L_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|4  6.348e-12
L_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7  5.197e-12
L_PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7 IG2_0_RX  2.058e-12
L_PTL_IG2_0|_RX|P1 _PTL_IG2_0|_RX|2 0  4.795e-13
L_PTL_IG2_0|_RX|P2 _PTL_IG2_0|_RX|5 0  5.431e-13
L_PTL_IG2_0|_RX|P3 _PTL_IG2_0|_RX|8 0  5.339e-13
R_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|101  4.225701121488
R_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|104  3.429952209
R_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|107  2.7439617672
L_PTL_IG2_0|_RX|RB1 _PTL_IG2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG2_0|_RX|RB2 _PTL_IG2_0|_RX|104 0  1.937922998085e-12
L_PTL_IG2_0|_RX|RB3 _PTL_IG2_0|_RX|107 0  1.550338398468e-12
B_PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_0|_TX|B1 0 _PTL_IP3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_0|_TX|B2 0 _PTL_IP3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|3  1.684e-12
L_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|6  3.596e-12
L_PTL_IP3_0|_TX|1 IP3_0 _PTL_IP3_0|_TX|1  2.063e-12
L_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|4  4.123e-12
L_PTL_IP3_0|_TX|3 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|7  2.193e-12
R_PTL_IP3_0|_TX|D _PTL_IP3_0|_TX|7 _PTL_IP3_0|A_PTL  1.36
L_PTL_IP3_0|_TX|P1 _PTL_IP3_0|_TX|2 0  5.254e-13
L_PTL_IP3_0|_TX|P2 _PTL_IP3_0|_TX|5 0  5.141e-13
R_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|101  2.7439617672
R_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|104  2.7439617672
L_PTL_IP3_0|_TX|RB1 _PTL_IP3_0|_TX|101 0  1.550338398468e-12
L_PTL_IP3_0|_TX|RB2 _PTL_IP3_0|_TX|104 0  1.550338398468e-12
B_PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_0|_RX|B1 0 _PTL_IP3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|3  2.777e-12
I_PTL_IP3_0|_RX|B2 0 _PTL_IP3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|6  2.685e-12
I_PTL_IP3_0|_RX|B3 0 _PTL_IP3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|9  2.764e-12
L_PTL_IP3_0|_RX|1 _PTL_IP3_0|A_PTL _PTL_IP3_0|_RX|1  1.346e-12
L_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|4  6.348e-12
L_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7  5.197e-12
L_PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7 IP3_0_RX  2.058e-12
L_PTL_IP3_0|_RX|P1 _PTL_IP3_0|_RX|2 0  4.795e-13
L_PTL_IP3_0|_RX|P2 _PTL_IP3_0|_RX|5 0  5.431e-13
L_PTL_IP3_0|_RX|P3 _PTL_IP3_0|_RX|8 0  5.339e-13
R_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|101  4.225701121488
R_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|104  3.429952209
R_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|107  2.7439617672
L_PTL_IP3_0|_RX|RB1 _PTL_IP3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_0|_RX|RB2 _PTL_IP3_0|_RX|104 0  1.937922998085e-12
L_PTL_IP3_0|_RX|RB3 _PTL_IP3_0|_RX|107 0  1.550338398468e-12
B_PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG3_0|_TX|B1 0 _PTL_IG3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG3_0|_TX|B2 0 _PTL_IG3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|3  1.684e-12
L_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|6  3.596e-12
L_PTL_IG3_0|_TX|1 IG3_0 _PTL_IG3_0|_TX|1  2.063e-12
L_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|4  4.123e-12
L_PTL_IG3_0|_TX|3 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|7  2.193e-12
R_PTL_IG3_0|_TX|D _PTL_IG3_0|_TX|7 _PTL_IG3_0|A_PTL  1.36
L_PTL_IG3_0|_TX|P1 _PTL_IG3_0|_TX|2 0  5.254e-13
L_PTL_IG3_0|_TX|P2 _PTL_IG3_0|_TX|5 0  5.141e-13
R_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|101  2.7439617672
R_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|104  2.7439617672
L_PTL_IG3_0|_TX|RB1 _PTL_IG3_0|_TX|101 0  1.550338398468e-12
L_PTL_IG3_0|_TX|RB2 _PTL_IG3_0|_TX|104 0  1.550338398468e-12
B_PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG3_0|_RX|B1 0 _PTL_IG3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|3  2.777e-12
I_PTL_IG3_0|_RX|B2 0 _PTL_IG3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|6  2.685e-12
I_PTL_IG3_0|_RX|B3 0 _PTL_IG3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|9  2.764e-12
L_PTL_IG3_0|_RX|1 _PTL_IG3_0|A_PTL _PTL_IG3_0|_RX|1  1.346e-12
L_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|4  6.348e-12
L_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7  5.197e-12
L_PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7 IG3_0_RX  2.058e-12
L_PTL_IG3_0|_RX|P1 _PTL_IG3_0|_RX|2 0  4.795e-13
L_PTL_IG3_0|_RX|P2 _PTL_IG3_0|_RX|5 0  5.431e-13
L_PTL_IG3_0|_RX|P3 _PTL_IG3_0|_RX|8 0  5.339e-13
R_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|101  4.225701121488
R_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|104  3.429952209
R_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|107  2.7439617672
L_PTL_IG3_0|_RX|RB1 _PTL_IG3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG3_0|_RX|RB2 _PTL_IG3_0|_RX|104 0  1.937922998085e-12
L_PTL_IG3_0|_RX|RB3 _PTL_IG3_0|_RX|107 0  1.550338398468e-12
LSPL_IG0_0|I_D1|B SPL_IG0_0|D1 SPL_IG0_0|I_D1|MID  2e-12
ISPL_IG0_0|I_D1|B 0 SPL_IG0_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_D2|B SPL_IG0_0|D2 SPL_IG0_0|I_D2|MID  2e-12
ISPL_IG0_0|I_D2|B 0 SPL_IG0_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG0_0|I_Q1|B SPL_IG0_0|QA1 SPL_IG0_0|I_Q1|MID  2e-12
ISPL_IG0_0|I_Q1|B 0 SPL_IG0_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_Q2|B SPL_IG0_0|QB1 SPL_IG0_0|I_Q2|MID  2e-12
ISPL_IG0_0|I_Q2|B 0 SPL_IG0_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG0_0|1|1 SPL_IG0_0|D1 SPL_IG0_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|1|P SPL_IG0_0|1|MID_SERIES 0  2e-13
RSPL_IG0_0|1|B SPL_IG0_0|D1 SPL_IG0_0|1|MID_SHUNT  2.7439617672
LSPL_IG0_0|1|RB SPL_IG0_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|2|1 SPL_IG0_0|D2 SPL_IG0_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|2|P SPL_IG0_0|2|MID_SERIES 0  2e-13
RSPL_IG0_0|2|B SPL_IG0_0|D2 SPL_IG0_0|2|MID_SHUNT  2.7439617672
LSPL_IG0_0|2|RB SPL_IG0_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|A|1 SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|A|P SPL_IG0_0|A|MID_SERIES 0  2e-13
RSPL_IG0_0|A|B SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SHUNT  2.7439617672
LSPL_IG0_0|A|RB SPL_IG0_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|B|1 SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|B|P SPL_IG0_0|B|MID_SERIES 0  2e-13
RSPL_IG0_0|B|B SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SHUNT  2.7439617672
LSPL_IG0_0|B|RB SPL_IG0_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP1_0|I_D1|B SPL_IP1_0|D1 SPL_IP1_0|I_D1|MID  2e-12
ISPL_IP1_0|I_D1|B 0 SPL_IP1_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_D2|B SPL_IP1_0|D2 SPL_IP1_0|I_D2|MID  2e-12
ISPL_IP1_0|I_D2|B 0 SPL_IP1_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP1_0|I_Q1|B SPL_IP1_0|QA1 SPL_IP1_0|I_Q1|MID  2e-12
ISPL_IP1_0|I_Q1|B 0 SPL_IP1_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_Q2|B SPL_IP1_0|QB1 SPL_IP1_0|I_Q2|MID  2e-12
ISPL_IP1_0|I_Q2|B 0 SPL_IP1_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP1_0|1|1 SPL_IP1_0|D1 SPL_IP1_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|1|P SPL_IP1_0|1|MID_SERIES 0  2e-13
RSPL_IP1_0|1|B SPL_IP1_0|D1 SPL_IP1_0|1|MID_SHUNT  2.7439617672
LSPL_IP1_0|1|RB SPL_IP1_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|2|1 SPL_IP1_0|D2 SPL_IP1_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|2|P SPL_IP1_0|2|MID_SERIES 0  2e-13
RSPL_IP1_0|2|B SPL_IP1_0|D2 SPL_IP1_0|2|MID_SHUNT  2.7439617672
LSPL_IP1_0|2|RB SPL_IP1_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|A|1 SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|A|P SPL_IP1_0|A|MID_SERIES 0  2e-13
RSPL_IP1_0|A|B SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SHUNT  2.7439617672
LSPL_IP1_0|A|RB SPL_IP1_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|B|1 SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|B|P SPL_IP1_0|B|MID_SERIES 0  2e-13
RSPL_IP1_0|B|B SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SHUNT  2.7439617672
LSPL_IP1_0|B|RB SPL_IP1_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|1 IP2_0_RX SPL_IP2_0|SPL1|D1  2e-12
LSPL_IP2_0|SPL1|2 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|D2  4.135667696e-12
LSPL_IP2_0|SPL1|3 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL1|4 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL1|5 SPL_IP2_0|SPL1|QA1 IP2_0_TO2  2e-12
LSPL_IP2_0|SPL1|6 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL1|7 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|QTMP  2e-12
LSPL_IP2_0|SPL2|1 SPL_IP2_0|QTMP SPL_IP2_0|SPL2|D1  2e-12
LSPL_IP2_0|SPL2|2 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|D2  4.135667696e-12
LSPL_IP2_0|SPL2|3 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL2|4 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL2|5 SPL_IP2_0|SPL2|QA1 IP2_0_TO3  2e-12
LSPL_IP2_0|SPL2|6 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL2|7 SPL_IP2_0|SPL2|QB1 IP2_0_OUT  2e-12
LSPL_IG2_0|I_D1|B SPL_IG2_0|D1 SPL_IG2_0|I_D1|MID  2e-12
ISPL_IG2_0|I_D1|B 0 SPL_IG2_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_D2|B SPL_IG2_0|D2 SPL_IG2_0|I_D2|MID  2e-12
ISPL_IG2_0|I_D2|B 0 SPL_IG2_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG2_0|I_Q1|B SPL_IG2_0|QA1 SPL_IG2_0|I_Q1|MID  2e-12
ISPL_IG2_0|I_Q1|B 0 SPL_IG2_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_Q2|B SPL_IG2_0|QB1 SPL_IG2_0|I_Q2|MID  2e-12
ISPL_IG2_0|I_Q2|B 0 SPL_IG2_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG2_0|1|1 SPL_IG2_0|D1 SPL_IG2_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|1|P SPL_IG2_0|1|MID_SERIES 0  2e-13
RSPL_IG2_0|1|B SPL_IG2_0|D1 SPL_IG2_0|1|MID_SHUNT  2.7439617672
LSPL_IG2_0|1|RB SPL_IG2_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|2|1 SPL_IG2_0|D2 SPL_IG2_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|2|P SPL_IG2_0|2|MID_SERIES 0  2e-13
RSPL_IG2_0|2|B SPL_IG2_0|D2 SPL_IG2_0|2|MID_SHUNT  2.7439617672
LSPL_IG2_0|2|RB SPL_IG2_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|A|1 SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|A|P SPL_IG2_0|A|MID_SERIES 0  2e-13
RSPL_IG2_0|A|B SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SHUNT  2.7439617672
LSPL_IG2_0|A|RB SPL_IG2_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|B|1 SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|B|P SPL_IG2_0|B|MID_SERIES 0  2e-13
RSPL_IG2_0|B|B SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SHUNT  2.7439617672
LSPL_IG2_0|B|RB SPL_IG2_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP3_0|I_D1|B SPL_IP3_0|D1 SPL_IP3_0|I_D1|MID  2e-12
ISPL_IP3_0|I_D1|B 0 SPL_IP3_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_D2|B SPL_IP3_0|D2 SPL_IP3_0|I_D2|MID  2e-12
ISPL_IP3_0|I_D2|B 0 SPL_IP3_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP3_0|I_Q1|B SPL_IP3_0|QA1 SPL_IP3_0|I_Q1|MID  2e-12
ISPL_IP3_0|I_Q1|B 0 SPL_IP3_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_Q2|B SPL_IP3_0|QB1 SPL_IP3_0|I_Q2|MID  2e-12
ISPL_IP3_0|I_Q2|B 0 SPL_IP3_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP3_0|1|1 SPL_IP3_0|D1 SPL_IP3_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|1|P SPL_IP3_0|1|MID_SERIES 0  2e-13
RSPL_IP3_0|1|B SPL_IP3_0|D1 SPL_IP3_0|1|MID_SHUNT  2.7439617672
LSPL_IP3_0|1|RB SPL_IP3_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|2|1 SPL_IP3_0|D2 SPL_IP3_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|2|P SPL_IP3_0|2|MID_SERIES 0  2e-13
RSPL_IP3_0|2|B SPL_IP3_0|D2 SPL_IP3_0|2|MID_SHUNT  2.7439617672
LSPL_IP3_0|2|RB SPL_IP3_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|A|1 SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|A|P SPL_IP3_0|A|MID_SERIES 0  2e-13
RSPL_IP3_0|A|B SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SHUNT  2.7439617672
LSPL_IP3_0|A|RB SPL_IP3_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|B|1 SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|B|P SPL_IP3_0|B|MID_SERIES 0  2e-13
RSPL_IP3_0|B|B SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SHUNT  2.7439617672
LSPL_IP3_0|B|RB SPL_IP3_0|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|1 IP0_0_RX _PG0_01|P|A1  2.067833848e-12
L_PG0_01|P|2 _PG0_01|P|A1 _PG0_01|P|A2  4.135667696e-12
L_PG0_01|P|3 _PG0_01|P|A3 _PG0_01|P|A4  8.271335392e-12
L_PG0_01|P|T T04 _PG0_01|P|T1  2.067833848e-12
L_PG0_01|P|4 _PG0_01|P|T1 _PG0_01|P|T2  4.135667696e-12
L_PG0_01|P|5 _PG0_01|P|A4 _PG0_01|P|Q1  4.135667696e-12
L_PG0_01|P|6 _PG0_01|P|Q1 P0_1  2.067833848e-12
L_PG0_01|G|1 IG0_0_TO0 _PG0_01|G|A1  2.067833848e-12
L_PG0_01|G|2 _PG0_01|G|A1 _PG0_01|G|A2  4.135667696e-12
L_PG0_01|G|3 _PG0_01|G|A3 _PG0_01|G|A4  8.271335392e-12
L_PG0_01|G|T T04 _PG0_01|G|T1  2.067833848e-12
L_PG0_01|G|4 _PG0_01|G|T1 _PG0_01|G|T2  4.135667696e-12
L_PG0_01|G|5 _PG0_01|G|A4 _PG0_01|G|Q1  4.135667696e-12
L_PG0_01|G|6 _PG0_01|G|Q1 G0_1  2.067833848e-12
L_PG1_01|_SPL_G1|1 IG1_0_RX _PG1_01|_SPL_G1|D1  2e-12
L_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|D2  4.135667696e-12
L_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG1_01|_SPL_G1|5 _PG1_01|_SPL_G1|QA1 _PG1_01|G1_COPY_1  2e-12
L_PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|QB1 _PG1_01|G1_COPY_2  2e-12
L_PG1_01|_PG|A1 IP1_0_TO1 _PG1_01|_PG|A1  2.067833848e-12
L_PG1_01|_PG|A2 _PG1_01|_PG|A1 _PG1_01|_PG|A2  4.135667696e-12
L_PG1_01|_PG|A3 _PG1_01|_PG|A3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|B1 _PG1_01|G1_COPY_1 _PG1_01|_PG|B1  2.067833848e-12
L_PG1_01|_PG|B2 _PG1_01|_PG|B1 _PG1_01|_PG|B2  4.135667696e-12
L_PG1_01|_PG|B3 _PG1_01|_PG|B3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|Q3 _PG1_01|_PG|Q3 _PG1_01|_PG|Q2  4.135667696e-12
L_PG1_01|_PG|Q2 _PG1_01|_PG|Q2 _PG1_01|_PG|Q1  4.135667696e-12
L_PG1_01|_PG|Q1 _PG1_01|_PG|Q1 _PG1_01|PG  2.067833848e-12
L_PG1_01|_GG|A1 IG0_0_TO1 _PG1_01|_GG|A1  2.067833848e-12
L_PG1_01|_GG|A2 _PG1_01|_GG|A1 _PG1_01|_GG|A2  4.135667696e-12
L_PG1_01|_GG|A3 _PG1_01|_GG|A3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|B1 _PG1_01|G1_COPY_2 _PG1_01|_GG|B1  2.067833848e-12
L_PG1_01|_GG|B2 _PG1_01|_GG|B1 _PG1_01|_GG|B2  4.135667696e-12
L_PG1_01|_GG|B3 _PG1_01|_GG|B3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|Q3 _PG1_01|_GG|Q3 _PG1_01|_GG|Q2  4.135667696e-12
L_PG1_01|_GG|Q2 _PG1_01|_GG|Q2 _PG1_01|_GG|Q1  4.135667696e-12
L_PG1_01|_GG|Q1 _PG1_01|_GG|Q1 _PG1_01|GG  2.067833848e-12
L_PG1_01|_DFF_PG|1 _PG1_01|PG _PG1_01|_DFF_PG|A1  2.067833848e-12
L_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|A2  4.135667696e-12
L_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|A4  8.271335392e-12
L_PG1_01|_DFF_PG|T T05 _PG1_01|_DFF_PG|T1  2.067833848e-12
L_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T2  4.135667696e-12
L_PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|Q1  4.135667696e-12
L_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|Q1 _PG1_01|PG_SYNC  2.067833848e-12
L_PG1_01|_DFF_GG|1 _PG1_01|GG _PG1_01|_DFF_GG|A1  2.067833848e-12
L_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|A2  4.135667696e-12
L_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|A4  8.271335392e-12
L_PG1_01|_DFF_GG|T T05 _PG1_01|_DFF_GG|T1  2.067833848e-12
L_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T2  4.135667696e-12
L_PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|Q1  4.135667696e-12
L_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|Q1 _PG1_01|GG_SYNC  2.067833848e-12
L_PG1_01|_AND_G|A1 _PG1_01|PG_SYNC _PG1_01|_AND_G|A1  2.067833848e-12
L_PG1_01|_AND_G|A2 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A2  4.135667696e-12
L_PG1_01|_AND_G|A3 _PG1_01|_AND_G|A3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|B1 _PG1_01|GG_SYNC _PG1_01|_AND_G|B1  2.067833848e-12
L_PG1_01|_AND_G|B2 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B2  4.135667696e-12
L_PG1_01|_AND_G|B3 _PG1_01|_AND_G|B3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q2  4.135667696e-12
L_PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q1  4.135667696e-12
L_PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1 G1_1  2.067833848e-12
L_PG2_01|P|1 IP2_0_TO2 _PG2_01|P|A1  2.067833848e-12
L_PG2_01|P|2 _PG2_01|P|A1 _PG2_01|P|A2  4.135667696e-12
L_PG2_01|P|3 _PG2_01|P|A3 _PG2_01|P|A4  8.271335392e-12
L_PG2_01|P|T T06 _PG2_01|P|T1  2.067833848e-12
L_PG2_01|P|4 _PG2_01|P|T1 _PG2_01|P|T2  4.135667696e-12
L_PG2_01|P|5 _PG2_01|P|A4 _PG2_01|P|Q1  4.135667696e-12
L_PG2_01|P|6 _PG2_01|P|Q1 P2_1  2.067833848e-12
L_PG2_01|G|1 IG2_0_TO2 _PG2_01|G|A1  2.067833848e-12
L_PG2_01|G|2 _PG2_01|G|A1 _PG2_01|G|A2  4.135667696e-12
L_PG2_01|G|3 _PG2_01|G|A3 _PG2_01|G|A4  8.271335392e-12
L_PG2_01|G|T T06 _PG2_01|G|T1  2.067833848e-12
L_PG2_01|G|4 _PG2_01|G|T1 _PG2_01|G|T2  4.135667696e-12
L_PG2_01|G|5 _PG2_01|G|A4 _PG2_01|G|Q1  4.135667696e-12
L_PG2_01|G|6 _PG2_01|G|Q1 G2_1  2.067833848e-12
L_PG3_01|_SPL_G1|1 IG3_0_RX _PG3_01|_SPL_G1|D1  2e-12
L_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|D2  4.135667696e-12
L_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_G1|5 _PG3_01|_SPL_G1|QA1 _PG3_01|G1_COPY_1  2e-12
L_PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|QB1 _PG3_01|G1_COPY_2  2e-12
L_PG3_01|_SPL_P1|1 IP3_0_TO1 _PG3_01|_SPL_P1|D1  2e-12
L_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|D2  4.135667696e-12
L_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_P1|5 _PG3_01|_SPL_P1|QA1 _PG3_01|P1_COPY_1  2e-12
L_PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|QB1 _PG3_01|P1_COPY_2  2e-12
L_PG3_01|_PG|A1 _PG3_01|P1_COPY_1 _PG3_01|_PG|A1  2.067833848e-12
L_PG3_01|_PG|A2 _PG3_01|_PG|A1 _PG3_01|_PG|A2  4.135667696e-12
L_PG3_01|_PG|A3 _PG3_01|_PG|A3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|B1 _PG3_01|G1_COPY_1 _PG3_01|_PG|B1  2.067833848e-12
L_PG3_01|_PG|B2 _PG3_01|_PG|B1 _PG3_01|_PG|B2  4.135667696e-12
L_PG3_01|_PG|B3 _PG3_01|_PG|B3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|Q3 _PG3_01|_PG|Q3 _PG3_01|_PG|Q2  4.135667696e-12
L_PG3_01|_PG|Q2 _PG3_01|_PG|Q2 _PG3_01|_PG|Q1  4.135667696e-12
L_PG3_01|_PG|Q1 _PG3_01|_PG|Q1 _PG3_01|PG  2.067833848e-12
L_PG3_01|_GG|A1 IG2_0_TO3 _PG3_01|_GG|A1  2.067833848e-12
L_PG3_01|_GG|A2 _PG3_01|_GG|A1 _PG3_01|_GG|A2  4.135667696e-12
L_PG3_01|_GG|A3 _PG3_01|_GG|A3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|B1 _PG3_01|G1_COPY_2 _PG3_01|_GG|B1  2.067833848e-12
L_PG3_01|_GG|B2 _PG3_01|_GG|B1 _PG3_01|_GG|B2  4.135667696e-12
L_PG3_01|_GG|B3 _PG3_01|_GG|B3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|Q3 _PG3_01|_GG|Q3 _PG3_01|_GG|Q2  4.135667696e-12
L_PG3_01|_GG|Q2 _PG3_01|_GG|Q2 _PG3_01|_GG|Q1  4.135667696e-12
L_PG3_01|_GG|Q1 _PG3_01|_GG|Q1 _PG3_01|GG  2.067833848e-12
L_PG3_01|_DFF_P0|1 IP2_0_TO3 _PG3_01|_DFF_P0|A1  2.067833848e-12
L_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|A2  4.135667696e-12
L_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|A4  8.271335392e-12
L_PG3_01|_DFF_P0|T T07 _PG3_01|_DFF_P0|T1  2.067833848e-12
L_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T2  4.135667696e-12
L_PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|Q1  4.135667696e-12
L_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|Q1 _PG3_01|P0_SYNC  2.067833848e-12
L_PG3_01|_DFF_P1|1 _PG3_01|P1_COPY_2 _PG3_01|_DFF_P1|A1  2.067833848e-12
L_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|A2  4.135667696e-12
L_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|A4  8.271335392e-12
L_PG3_01|_DFF_P1|T T07 _PG3_01|_DFF_P1|T1  2.067833848e-12
L_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T2  4.135667696e-12
L_PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|Q1  4.135667696e-12
L_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|Q1 _PG3_01|P1_SYNC  2.067833848e-12
L_PG3_01|_DFF_PG|1 _PG3_01|PG _PG3_01|_DFF_PG|A1  2.067833848e-12
L_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|A2  4.135667696e-12
L_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|A4  8.271335392e-12
L_PG3_01|_DFF_PG|T T07 _PG3_01|_DFF_PG|T1  2.067833848e-12
L_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T2  4.135667696e-12
L_PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|Q1  4.135667696e-12
L_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|Q1 _PG3_01|PG_SYNC  2.067833848e-12
L_PG3_01|_DFF_GG|1 _PG3_01|GG _PG3_01|_DFF_GG|A1  2.067833848e-12
L_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|A2  4.135667696e-12
L_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|A4  8.271335392e-12
L_PG3_01|_DFF_GG|T T07 _PG3_01|_DFF_GG|T1  2.067833848e-12
L_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T2  4.135667696e-12
L_PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|Q1  4.135667696e-12
L_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|Q1 _PG3_01|GG_SYNC  2.067833848e-12
L_PG3_01|_AND_G|A1 _PG3_01|PG_SYNC _PG3_01|_AND_G|A1  2.067833848e-12
L_PG3_01|_AND_G|A2 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A2  4.135667696e-12
L_PG3_01|_AND_G|A3 _PG3_01|_AND_G|A3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|B1 _PG3_01|GG_SYNC _PG3_01|_AND_G|B1  2.067833848e-12
L_PG3_01|_AND_G|B2 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B2  4.135667696e-12
L_PG3_01|_AND_G|B3 _PG3_01|_AND_G|B3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q2  4.135667696e-12
L_PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q1  4.135667696e-12
L_PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1 G3_1  2.067833848e-12
L_PG3_01|_AND_P|A1 _PG3_01|P0_SYNC _PG3_01|_AND_P|A1  2.067833848e-12
L_PG3_01|_AND_P|A2 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A2  4.135667696e-12
L_PG3_01|_AND_P|A3 _PG3_01|_AND_P|A3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|B1 _PG3_01|P1_SYNC _PG3_01|_AND_P|B1  2.067833848e-12
L_PG3_01|_AND_P|B2 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B2  4.135667696e-12
L_PG3_01|_AND_P|B3 _PG3_01|_AND_P|B3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q2  4.135667696e-12
L_PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q1  4.135667696e-12
L_PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1 P3_1  2.067833848e-12
L_DFF_IP1_01|I_1|B _DFF_IP1_01|A1 _DFF_IP1_01|I_1|MID  2e-12
I_DFF_IP1_01|I_1|B 0 _DFF_IP1_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_3|B _DFF_IP1_01|A3 _DFF_IP1_01|I_3|MID  2e-12
I_DFF_IP1_01|I_3|B 0 _DFF_IP1_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_01|I_T|B _DFF_IP1_01|T1 _DFF_IP1_01|I_T|MID  2e-12
I_DFF_IP1_01|I_T|B 0 _DFF_IP1_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_6|B _DFF_IP1_01|Q1 _DFF_IP1_01|I_6|MID  2e-12
I_DFF_IP1_01|I_6|B 0 _DFF_IP1_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_01|1|1 _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|1|P _DFF_IP1_01|1|MID_SERIES 0  2e-13
R_DFF_IP1_01|1|B _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SHUNT  2.7439617672
L_DFF_IP1_01|1|RB _DFF_IP1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|23|1 _DFF_IP1_01|A2 _DFF_IP1_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|23|B _DFF_IP1_01|A2 _DFF_IP1_01|23|MID_SHUNT  3.84154647408
L_DFF_IP1_01|23|RB _DFF_IP1_01|23|MID_SHUNT _DFF_IP1_01|A3  2.1704737578552e-12
B_DFF_IP1_01|3|1 _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|3|P _DFF_IP1_01|3|MID_SERIES 0  2e-13
R_DFF_IP1_01|3|B _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SHUNT  2.7439617672
L_DFF_IP1_01|3|RB _DFF_IP1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|4|1 _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|4|P _DFF_IP1_01|4|MID_SERIES 0  2e-13
R_DFF_IP1_01|4|B _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SHUNT  2.7439617672
L_DFF_IP1_01|4|RB _DFF_IP1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|T|1 _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|T|P _DFF_IP1_01|T|MID_SERIES 0  2e-13
R_DFF_IP1_01|T|B _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SHUNT  2.7439617672
L_DFF_IP1_01|T|RB _DFF_IP1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|45|1 _DFF_IP1_01|T2 _DFF_IP1_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|45|B _DFF_IP1_01|T2 _DFF_IP1_01|45|MID_SHUNT  3.84154647408
L_DFF_IP1_01|45|RB _DFF_IP1_01|45|MID_SHUNT _DFF_IP1_01|A4  2.1704737578552e-12
B_DFF_IP1_01|6|1 _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|6|P _DFF_IP1_01|6|MID_SERIES 0  2e-13
R_DFF_IP1_01|6|B _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SHUNT  2.7439617672
L_DFF_IP1_01|6|RB _DFF_IP1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_01|I_1|B _DFF_IP2_01|A1 _DFF_IP2_01|I_1|MID  2e-12
I_DFF_IP2_01|I_1|B 0 _DFF_IP2_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_3|B _DFF_IP2_01|A3 _DFF_IP2_01|I_3|MID  2e-12
I_DFF_IP2_01|I_3|B 0 _DFF_IP2_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_01|I_T|B _DFF_IP2_01|T1 _DFF_IP2_01|I_T|MID  2e-12
I_DFF_IP2_01|I_T|B 0 _DFF_IP2_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_6|B _DFF_IP2_01|Q1 _DFF_IP2_01|I_6|MID  2e-12
I_DFF_IP2_01|I_6|B 0 _DFF_IP2_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_01|1|1 _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|1|P _DFF_IP2_01|1|MID_SERIES 0  2e-13
R_DFF_IP2_01|1|B _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SHUNT  2.7439617672
L_DFF_IP2_01|1|RB _DFF_IP2_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|23|1 _DFF_IP2_01|A2 _DFF_IP2_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|23|B _DFF_IP2_01|A2 _DFF_IP2_01|23|MID_SHUNT  3.84154647408
L_DFF_IP2_01|23|RB _DFF_IP2_01|23|MID_SHUNT _DFF_IP2_01|A3  2.1704737578552e-12
B_DFF_IP2_01|3|1 _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|3|P _DFF_IP2_01|3|MID_SERIES 0  2e-13
R_DFF_IP2_01|3|B _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SHUNT  2.7439617672
L_DFF_IP2_01|3|RB _DFF_IP2_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|4|1 _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|4|P _DFF_IP2_01|4|MID_SERIES 0  2e-13
R_DFF_IP2_01|4|B _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SHUNT  2.7439617672
L_DFF_IP2_01|4|RB _DFF_IP2_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|T|1 _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|T|P _DFF_IP2_01|T|MID_SERIES 0  2e-13
R_DFF_IP2_01|T|B _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SHUNT  2.7439617672
L_DFF_IP2_01|T|RB _DFF_IP2_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|45|1 _DFF_IP2_01|T2 _DFF_IP2_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|45|B _DFF_IP2_01|T2 _DFF_IP2_01|45|MID_SHUNT  3.84154647408
L_DFF_IP2_01|45|RB _DFF_IP2_01|45|MID_SHUNT _DFF_IP2_01|A4  2.1704737578552e-12
B_DFF_IP2_01|6|1 _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|6|P _DFF_IP2_01|6|MID_SERIES 0  2e-13
R_DFF_IP2_01|6|B _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SHUNT  2.7439617672
L_DFF_IP2_01|6|RB _DFF_IP2_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_01|I_1|B _DFF_IP3_01|A1 _DFF_IP3_01|I_1|MID  2e-12
I_DFF_IP3_01|I_1|B 0 _DFF_IP3_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_3|B _DFF_IP3_01|A3 _DFF_IP3_01|I_3|MID  2e-12
I_DFF_IP3_01|I_3|B 0 _DFF_IP3_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_01|I_T|B _DFF_IP3_01|T1 _DFF_IP3_01|I_T|MID  2e-12
I_DFF_IP3_01|I_T|B 0 _DFF_IP3_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_6|B _DFF_IP3_01|Q1 _DFF_IP3_01|I_6|MID  2e-12
I_DFF_IP3_01|I_6|B 0 _DFF_IP3_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_01|1|1 _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|1|P _DFF_IP3_01|1|MID_SERIES 0  2e-13
R_DFF_IP3_01|1|B _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SHUNT  2.7439617672
L_DFF_IP3_01|1|RB _DFF_IP3_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|23|1 _DFF_IP3_01|A2 _DFF_IP3_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|23|B _DFF_IP3_01|A2 _DFF_IP3_01|23|MID_SHUNT  3.84154647408
L_DFF_IP3_01|23|RB _DFF_IP3_01|23|MID_SHUNT _DFF_IP3_01|A3  2.1704737578552e-12
B_DFF_IP3_01|3|1 _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|3|P _DFF_IP3_01|3|MID_SERIES 0  2e-13
R_DFF_IP3_01|3|B _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SHUNT  2.7439617672
L_DFF_IP3_01|3|RB _DFF_IP3_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|4|1 _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|4|P _DFF_IP3_01|4|MID_SERIES 0  2e-13
R_DFF_IP3_01|4|B _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SHUNT  2.7439617672
L_DFF_IP3_01|4|RB _DFF_IP3_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|T|1 _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|T|P _DFF_IP3_01|T|MID_SERIES 0  2e-13
R_DFF_IP3_01|T|B _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SHUNT  2.7439617672
L_DFF_IP3_01|T|RB _DFF_IP3_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|45|1 _DFF_IP3_01|T2 _DFF_IP3_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|45|B _DFF_IP3_01|T2 _DFF_IP3_01|45|MID_SHUNT  3.84154647408
L_DFF_IP3_01|45|RB _DFF_IP3_01|45|MID_SHUNT _DFF_IP3_01|A4  2.1704737578552e-12
B_DFF_IP3_01|6|1 _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|6|P _DFF_IP3_01|6|MID_SERIES 0  2e-13
R_DFF_IP3_01|6|B _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SHUNT  2.7439617672
L_DFF_IP3_01|6|RB _DFF_IP3_01|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_P0_1|_TX|1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|2 JJMIT AREA=2.5
B_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|5 JJMIT AREA=2.5
I_PTL_P0_1|_TX|B1 0 _PTL_P0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_1|_TX|B2 0 _PTL_P0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|3  1.684e-12
L_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|6  3.596e-12
L_PTL_P0_1|_TX|1 P0_1 _PTL_P0_1|_TX|1  2.063e-12
L_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|4  4.123e-12
L_PTL_P0_1|_TX|3 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|7  2.193e-12
R_PTL_P0_1|_TX|D _PTL_P0_1|_TX|7 _PTL_P0_1|A_PTL  1.36
L_PTL_P0_1|_TX|P1 _PTL_P0_1|_TX|2 0  5.254e-13
L_PTL_P0_1|_TX|P2 _PTL_P0_1|_TX|5 0  5.141e-13
R_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|101  2.7439617672
R_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|104  2.7439617672
L_PTL_P0_1|_TX|RB1 _PTL_P0_1|_TX|101 0  1.550338398468e-12
L_PTL_P0_1|_TX|RB2 _PTL_P0_1|_TX|104 0  1.550338398468e-12
B_PTL_P0_1|_RX|1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|5 JJMIT AREA=2.0
B_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|8 JJMIT AREA=2.5
I_PTL_P0_1|_RX|B1 0 _PTL_P0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|3  2.777e-12
I_PTL_P0_1|_RX|B2 0 _PTL_P0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|6  2.685e-12
I_PTL_P0_1|_RX|B3 0 _PTL_P0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|9  2.764e-12
L_PTL_P0_1|_RX|1 _PTL_P0_1|A_PTL _PTL_P0_1|_RX|1  1.346e-12
L_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|4  6.348e-12
L_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7  5.197e-12
L_PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7 P0_1_RX  2.058e-12
L_PTL_P0_1|_RX|P1 _PTL_P0_1|_RX|2 0  4.795e-13
L_PTL_P0_1|_RX|P2 _PTL_P0_1|_RX|5 0  5.431e-13
L_PTL_P0_1|_RX|P3 _PTL_P0_1|_RX|8 0  5.339e-13
R_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|101  4.225701121488
R_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|104  3.429952209
R_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|107  2.7439617672
L_PTL_P0_1|_RX|RB1 _PTL_P0_1|_RX|101 0  2.38752113364072e-12
L_PTL_P0_1|_RX|RB2 _PTL_P0_1|_RX|104 0  1.937922998085e-12
L_PTL_P0_1|_RX|RB3 _PTL_P0_1|_RX|107 0  1.550338398468e-12
B_PTL_G0_1|_TX|1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|2 JJMIT AREA=2.5
B_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|5 JJMIT AREA=2.5
I_PTL_G0_1|_TX|B1 0 _PTL_G0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_1|_TX|B2 0 _PTL_G0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|3  1.684e-12
L_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|6  3.596e-12
L_PTL_G0_1|_TX|1 G0_1 _PTL_G0_1|_TX|1  2.063e-12
L_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|4  4.123e-12
L_PTL_G0_1|_TX|3 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|7  2.193e-12
R_PTL_G0_1|_TX|D _PTL_G0_1|_TX|7 _PTL_G0_1|A_PTL  1.36
L_PTL_G0_1|_TX|P1 _PTL_G0_1|_TX|2 0  5.254e-13
L_PTL_G0_1|_TX|P2 _PTL_G0_1|_TX|5 0  5.141e-13
R_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|101  2.7439617672
R_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|104  2.7439617672
L_PTL_G0_1|_TX|RB1 _PTL_G0_1|_TX|101 0  1.550338398468e-12
L_PTL_G0_1|_TX|RB2 _PTL_G0_1|_TX|104 0  1.550338398468e-12
B_PTL_G0_1|_RX|1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|5 JJMIT AREA=2.0
B_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|8 JJMIT AREA=2.5
I_PTL_G0_1|_RX|B1 0 _PTL_G0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|3  2.777e-12
I_PTL_G0_1|_RX|B2 0 _PTL_G0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|6  2.685e-12
I_PTL_G0_1|_RX|B3 0 _PTL_G0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|9  2.764e-12
L_PTL_G0_1|_RX|1 _PTL_G0_1|A_PTL _PTL_G0_1|_RX|1  1.346e-12
L_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|4  6.348e-12
L_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7  5.197e-12
L_PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7 G0_1_RX  2.058e-12
L_PTL_G0_1|_RX|P1 _PTL_G0_1|_RX|2 0  4.795e-13
L_PTL_G0_1|_RX|P2 _PTL_G0_1|_RX|5 0  5.431e-13
L_PTL_G0_1|_RX|P3 _PTL_G0_1|_RX|8 0  5.339e-13
R_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|101  4.225701121488
R_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|104  3.429952209
R_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|107  2.7439617672
L_PTL_G0_1|_RX|RB1 _PTL_G0_1|_RX|101 0  2.38752113364072e-12
L_PTL_G0_1|_RX|RB2 _PTL_G0_1|_RX|104 0  1.937922998085e-12
L_PTL_G0_1|_RX|RB3 _PTL_G0_1|_RX|107 0  1.550338398468e-12
B_PTL_G1_1|_TX|1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|2 JJMIT AREA=2.5
B_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|5 JJMIT AREA=2.5
I_PTL_G1_1|_TX|B1 0 _PTL_G1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_1|_TX|B2 0 _PTL_G1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|3  1.684e-12
L_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|6  3.596e-12
L_PTL_G1_1|_TX|1 G1_1 _PTL_G1_1|_TX|1  2.063e-12
L_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|4  4.123e-12
L_PTL_G1_1|_TX|3 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|7  2.193e-12
R_PTL_G1_1|_TX|D _PTL_G1_1|_TX|7 _PTL_G1_1|A_PTL  1.36
L_PTL_G1_1|_TX|P1 _PTL_G1_1|_TX|2 0  5.254e-13
L_PTL_G1_1|_TX|P2 _PTL_G1_1|_TX|5 0  5.141e-13
R_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|101  2.7439617672
R_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|104  2.7439617672
L_PTL_G1_1|_TX|RB1 _PTL_G1_1|_TX|101 0  1.550338398468e-12
L_PTL_G1_1|_TX|RB2 _PTL_G1_1|_TX|104 0  1.550338398468e-12
B_PTL_G1_1|_RX|1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|5 JJMIT AREA=2.0
B_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|8 JJMIT AREA=2.5
I_PTL_G1_1|_RX|B1 0 _PTL_G1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|3  2.777e-12
I_PTL_G1_1|_RX|B2 0 _PTL_G1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|6  2.685e-12
I_PTL_G1_1|_RX|B3 0 _PTL_G1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|9  2.764e-12
L_PTL_G1_1|_RX|1 _PTL_G1_1|A_PTL _PTL_G1_1|_RX|1  1.346e-12
L_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|4  6.348e-12
L_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7  5.197e-12
L_PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7 G1_1_RX  2.058e-12
L_PTL_G1_1|_RX|P1 _PTL_G1_1|_RX|2 0  4.795e-13
L_PTL_G1_1|_RX|P2 _PTL_G1_1|_RX|5 0  5.431e-13
L_PTL_G1_1|_RX|P3 _PTL_G1_1|_RX|8 0  5.339e-13
R_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|101  4.225701121488
R_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|104  3.429952209
R_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|107  2.7439617672
L_PTL_G1_1|_RX|RB1 _PTL_G1_1|_RX|101 0  2.38752113364072e-12
L_PTL_G1_1|_RX|RB2 _PTL_G1_1|_RX|104 0  1.937922998085e-12
L_PTL_G1_1|_RX|RB3 _PTL_G1_1|_RX|107 0  1.550338398468e-12
B_PTL_P2_1|_TX|1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|2 JJMIT AREA=2.5
B_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|5 JJMIT AREA=2.5
I_PTL_P2_1|_TX|B1 0 _PTL_P2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P2_1|_TX|B2 0 _PTL_P2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|3  1.684e-12
L_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|6  3.596e-12
L_PTL_P2_1|_TX|1 P2_1 _PTL_P2_1|_TX|1  2.063e-12
L_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|4  4.123e-12
L_PTL_P2_1|_TX|3 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|7  2.193e-12
R_PTL_P2_1|_TX|D _PTL_P2_1|_TX|7 _PTL_P2_1|A_PTL  1.36
L_PTL_P2_1|_TX|P1 _PTL_P2_1|_TX|2 0  5.254e-13
L_PTL_P2_1|_TX|P2 _PTL_P2_1|_TX|5 0  5.141e-13
R_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|101  2.7439617672
R_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|104  2.7439617672
L_PTL_P2_1|_TX|RB1 _PTL_P2_1|_TX|101 0  1.550338398468e-12
L_PTL_P2_1|_TX|RB2 _PTL_P2_1|_TX|104 0  1.550338398468e-12
B_PTL_P2_1|_RX|1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|5 JJMIT AREA=2.0
B_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|8 JJMIT AREA=2.5
I_PTL_P2_1|_RX|B1 0 _PTL_P2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|3  2.777e-12
I_PTL_P2_1|_RX|B2 0 _PTL_P2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|6  2.685e-12
I_PTL_P2_1|_RX|B3 0 _PTL_P2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|9  2.764e-12
L_PTL_P2_1|_RX|1 _PTL_P2_1|A_PTL _PTL_P2_1|_RX|1  1.346e-12
L_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|4  6.348e-12
L_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7  5.197e-12
L_PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7 P2_1_RX  2.058e-12
L_PTL_P2_1|_RX|P1 _PTL_P2_1|_RX|2 0  4.795e-13
L_PTL_P2_1|_RX|P2 _PTL_P2_1|_RX|5 0  5.431e-13
L_PTL_P2_1|_RX|P3 _PTL_P2_1|_RX|8 0  5.339e-13
R_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|101  4.225701121488
R_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|104  3.429952209
R_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|107  2.7439617672
L_PTL_P2_1|_RX|RB1 _PTL_P2_1|_RX|101 0  2.38752113364072e-12
L_PTL_P2_1|_RX|RB2 _PTL_P2_1|_RX|104 0  1.937922998085e-12
L_PTL_P2_1|_RX|RB3 _PTL_P2_1|_RX|107 0  1.550338398468e-12
B_PTL_G2_1|_TX|1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|2 JJMIT AREA=2.5
B_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|5 JJMIT AREA=2.5
I_PTL_G2_1|_TX|B1 0 _PTL_G2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_1|_TX|B2 0 _PTL_G2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|3  1.684e-12
L_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|6  3.596e-12
L_PTL_G2_1|_TX|1 G2_1 _PTL_G2_1|_TX|1  2.063e-12
L_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|4  4.123e-12
L_PTL_G2_1|_TX|3 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|7  2.193e-12
R_PTL_G2_1|_TX|D _PTL_G2_1|_TX|7 _PTL_G2_1|A_PTL  1.36
L_PTL_G2_1|_TX|P1 _PTL_G2_1|_TX|2 0  5.254e-13
L_PTL_G2_1|_TX|P2 _PTL_G2_1|_TX|5 0  5.141e-13
R_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|101  2.7439617672
R_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|104  2.7439617672
L_PTL_G2_1|_TX|RB1 _PTL_G2_1|_TX|101 0  1.550338398468e-12
L_PTL_G2_1|_TX|RB2 _PTL_G2_1|_TX|104 0  1.550338398468e-12
B_PTL_G2_1|_RX|1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|5 JJMIT AREA=2.0
B_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|8 JJMIT AREA=2.5
I_PTL_G2_1|_RX|B1 0 _PTL_G2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|3  2.777e-12
I_PTL_G2_1|_RX|B2 0 _PTL_G2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|6  2.685e-12
I_PTL_G2_1|_RX|B3 0 _PTL_G2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|9  2.764e-12
L_PTL_G2_1|_RX|1 _PTL_G2_1|A_PTL _PTL_G2_1|_RX|1  1.346e-12
L_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|4  6.348e-12
L_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7  5.197e-12
L_PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7 G2_1_RX  2.058e-12
L_PTL_G2_1|_RX|P1 _PTL_G2_1|_RX|2 0  4.795e-13
L_PTL_G2_1|_RX|P2 _PTL_G2_1|_RX|5 0  5.431e-13
L_PTL_G2_1|_RX|P3 _PTL_G2_1|_RX|8 0  5.339e-13
R_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|101  4.225701121488
R_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|104  3.429952209
R_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|107  2.7439617672
L_PTL_G2_1|_RX|RB1 _PTL_G2_1|_RX|101 0  2.38752113364072e-12
L_PTL_G2_1|_RX|RB2 _PTL_G2_1|_RX|104 0  1.937922998085e-12
L_PTL_G2_1|_RX|RB3 _PTL_G2_1|_RX|107 0  1.550338398468e-12
B_PTL_P3_1|_TX|1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|2 JJMIT AREA=2.5
B_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|5 JJMIT AREA=2.5
I_PTL_P3_1|_TX|B1 0 _PTL_P3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P3_1|_TX|B2 0 _PTL_P3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|3  1.684e-12
L_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|6  3.596e-12
L_PTL_P3_1|_TX|1 P3_1 _PTL_P3_1|_TX|1  2.063e-12
L_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|4  4.123e-12
L_PTL_P3_1|_TX|3 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|7  2.193e-12
R_PTL_P3_1|_TX|D _PTL_P3_1|_TX|7 _PTL_P3_1|A_PTL  1.36
L_PTL_P3_1|_TX|P1 _PTL_P3_1|_TX|2 0  5.254e-13
L_PTL_P3_1|_TX|P2 _PTL_P3_1|_TX|5 0  5.141e-13
R_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|101  2.7439617672
R_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|104  2.7439617672
L_PTL_P3_1|_TX|RB1 _PTL_P3_1|_TX|101 0  1.550338398468e-12
L_PTL_P3_1|_TX|RB2 _PTL_P3_1|_TX|104 0  1.550338398468e-12
B_PTL_P3_1|_RX|1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|5 JJMIT AREA=2.0
B_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|8 JJMIT AREA=2.5
I_PTL_P3_1|_RX|B1 0 _PTL_P3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|3  2.777e-12
I_PTL_P3_1|_RX|B2 0 _PTL_P3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|6  2.685e-12
I_PTL_P3_1|_RX|B3 0 _PTL_P3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|9  2.764e-12
L_PTL_P3_1|_RX|1 _PTL_P3_1|A_PTL _PTL_P3_1|_RX|1  1.346e-12
L_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|4  6.348e-12
L_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7  5.197e-12
L_PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7 P3_1_RX  2.058e-12
L_PTL_P3_1|_RX|P1 _PTL_P3_1|_RX|2 0  4.795e-13
L_PTL_P3_1|_RX|P2 _PTL_P3_1|_RX|5 0  5.431e-13
L_PTL_P3_1|_RX|P3 _PTL_P3_1|_RX|8 0  5.339e-13
R_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|101  4.225701121488
R_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|104  3.429952209
R_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|107  2.7439617672
L_PTL_P3_1|_RX|RB1 _PTL_P3_1|_RX|101 0  2.38752113364072e-12
L_PTL_P3_1|_RX|RB2 _PTL_P3_1|_RX|104 0  1.937922998085e-12
L_PTL_P3_1|_RX|RB3 _PTL_P3_1|_RX|107 0  1.550338398468e-12
B_PTL_G3_1|_TX|1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|2 JJMIT AREA=2.5
B_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|5 JJMIT AREA=2.5
I_PTL_G3_1|_TX|B1 0 _PTL_G3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_1|_TX|B2 0 _PTL_G3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|3  1.684e-12
L_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|6  3.596e-12
L_PTL_G3_1|_TX|1 G3_1 _PTL_G3_1|_TX|1  2.063e-12
L_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|4  4.123e-12
L_PTL_G3_1|_TX|3 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|7  2.193e-12
R_PTL_G3_1|_TX|D _PTL_G3_1|_TX|7 _PTL_G3_1|A_PTL  1.36
L_PTL_G3_1|_TX|P1 _PTL_G3_1|_TX|2 0  5.254e-13
L_PTL_G3_1|_TX|P2 _PTL_G3_1|_TX|5 0  5.141e-13
R_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|101  2.7439617672
R_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|104  2.7439617672
L_PTL_G3_1|_TX|RB1 _PTL_G3_1|_TX|101 0  1.550338398468e-12
L_PTL_G3_1|_TX|RB2 _PTL_G3_1|_TX|104 0  1.550338398468e-12
B_PTL_G3_1|_RX|1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|5 JJMIT AREA=2.0
B_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|8 JJMIT AREA=2.5
I_PTL_G3_1|_RX|B1 0 _PTL_G3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|3  2.777e-12
I_PTL_G3_1|_RX|B2 0 _PTL_G3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|6  2.685e-12
I_PTL_G3_1|_RX|B3 0 _PTL_G3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|9  2.764e-12
L_PTL_G3_1|_RX|1 _PTL_G3_1|A_PTL _PTL_G3_1|_RX|1  1.346e-12
L_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|4  6.348e-12
L_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7  5.197e-12
L_PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7 G3_1_RX  2.058e-12
L_PTL_G3_1|_RX|P1 _PTL_G3_1|_RX|2 0  4.795e-13
L_PTL_G3_1|_RX|P2 _PTL_G3_1|_RX|5 0  5.431e-13
L_PTL_G3_1|_RX|P3 _PTL_G3_1|_RX|8 0  5.339e-13
R_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|101  4.225701121488
R_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|104  3.429952209
R_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|107  2.7439617672
L_PTL_G3_1|_RX|RB1 _PTL_G3_1|_RX|101 0  2.38752113364072e-12
L_PTL_G3_1|_RX|RB2 _PTL_G3_1|_RX|104 0  1.937922998085e-12
L_PTL_G3_1|_RX|RB3 _PTL_G3_1|_RX|107 0  1.550338398468e-12
B_PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_1|_TX|B1 0 _PTL_IP1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_1|_TX|B2 0 _PTL_IP1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|3  1.684e-12
L_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|6  3.596e-12
L_PTL_IP1_1|_TX|1 IP1_1_OUT _PTL_IP1_1|_TX|1  2.063e-12
L_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|4  4.123e-12
L_PTL_IP1_1|_TX|3 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|7  2.193e-12
R_PTL_IP1_1|_TX|D _PTL_IP1_1|_TX|7 _PTL_IP1_1|A_PTL  1.36
L_PTL_IP1_1|_TX|P1 _PTL_IP1_1|_TX|2 0  5.254e-13
L_PTL_IP1_1|_TX|P2 _PTL_IP1_1|_TX|5 0  5.141e-13
R_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|101  2.7439617672
R_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|104  2.7439617672
L_PTL_IP1_1|_TX|RB1 _PTL_IP1_1|_TX|101 0  1.550338398468e-12
L_PTL_IP1_1|_TX|RB2 _PTL_IP1_1|_TX|104 0  1.550338398468e-12
B_PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_1|_RX|B1 0 _PTL_IP1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|3  2.777e-12
I_PTL_IP1_1|_RX|B2 0 _PTL_IP1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|6  2.685e-12
I_PTL_IP1_1|_RX|B3 0 _PTL_IP1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|9  2.764e-12
L_PTL_IP1_1|_RX|1 _PTL_IP1_1|A_PTL _PTL_IP1_1|_RX|1  1.346e-12
L_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|4  6.348e-12
L_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7  5.197e-12
L_PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7 IP1_1_OUT_RX  2.058e-12
L_PTL_IP1_1|_RX|P1 _PTL_IP1_1|_RX|2 0  4.795e-13
L_PTL_IP1_1|_RX|P2 _PTL_IP1_1|_RX|5 0  5.431e-13
L_PTL_IP1_1|_RX|P3 _PTL_IP1_1|_RX|8 0  5.339e-13
R_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|101  4.225701121488
R_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|104  3.429952209
R_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|107  2.7439617672
L_PTL_IP1_1|_RX|RB1 _PTL_IP1_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_1|_RX|RB2 _PTL_IP1_1|_RX|104 0  1.937922998085e-12
L_PTL_IP1_1|_RX|RB3 _PTL_IP1_1|_RX|107 0  1.550338398468e-12
B_PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_1|_TX|B1 0 _PTL_IP2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_1|_TX|B2 0 _PTL_IP2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|3  1.684e-12
L_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|6  3.596e-12
L_PTL_IP2_1|_TX|1 IP2_1_OUT _PTL_IP2_1|_TX|1  2.063e-12
L_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|4  4.123e-12
L_PTL_IP2_1|_TX|3 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|7  2.193e-12
R_PTL_IP2_1|_TX|D _PTL_IP2_1|_TX|7 _PTL_IP2_1|A_PTL  1.36
L_PTL_IP2_1|_TX|P1 _PTL_IP2_1|_TX|2 0  5.254e-13
L_PTL_IP2_1|_TX|P2 _PTL_IP2_1|_TX|5 0  5.141e-13
R_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|101  2.7439617672
R_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|104  2.7439617672
L_PTL_IP2_1|_TX|RB1 _PTL_IP2_1|_TX|101 0  1.550338398468e-12
L_PTL_IP2_1|_TX|RB2 _PTL_IP2_1|_TX|104 0  1.550338398468e-12
B_PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_1|_RX|B1 0 _PTL_IP2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|3  2.777e-12
I_PTL_IP2_1|_RX|B2 0 _PTL_IP2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|6  2.685e-12
I_PTL_IP2_1|_RX|B3 0 _PTL_IP2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|9  2.764e-12
L_PTL_IP2_1|_RX|1 _PTL_IP2_1|A_PTL _PTL_IP2_1|_RX|1  1.346e-12
L_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|4  6.348e-12
L_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7  5.197e-12
L_PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7 IP2_1_OUT_RX  2.058e-12
L_PTL_IP2_1|_RX|P1 _PTL_IP2_1|_RX|2 0  4.795e-13
L_PTL_IP2_1|_RX|P2 _PTL_IP2_1|_RX|5 0  5.431e-13
L_PTL_IP2_1|_RX|P3 _PTL_IP2_1|_RX|8 0  5.339e-13
R_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|101  4.225701121488
R_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|104  3.429952209
R_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|107  2.7439617672
L_PTL_IP2_1|_RX|RB1 _PTL_IP2_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_1|_RX|RB2 _PTL_IP2_1|_RX|104 0  1.937922998085e-12
L_PTL_IP2_1|_RX|RB3 _PTL_IP2_1|_RX|107 0  1.550338398468e-12
B_PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_1|_TX|B1 0 _PTL_IP3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_1|_TX|B2 0 _PTL_IP3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|3  1.684e-12
L_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|6  3.596e-12
L_PTL_IP3_1|_TX|1 IP3_1_OUT _PTL_IP3_1|_TX|1  2.063e-12
L_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|4  4.123e-12
L_PTL_IP3_1|_TX|3 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|7  2.193e-12
R_PTL_IP3_1|_TX|D _PTL_IP3_1|_TX|7 _PTL_IP3_1|A_PTL  1.36
L_PTL_IP3_1|_TX|P1 _PTL_IP3_1|_TX|2 0  5.254e-13
L_PTL_IP3_1|_TX|P2 _PTL_IP3_1|_TX|5 0  5.141e-13
R_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|101  2.7439617672
R_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|104  2.7439617672
L_PTL_IP3_1|_TX|RB1 _PTL_IP3_1|_TX|101 0  1.550338398468e-12
L_PTL_IP3_1|_TX|RB2 _PTL_IP3_1|_TX|104 0  1.550338398468e-12
B_PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_1|_RX|B1 0 _PTL_IP3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|3  2.777e-12
I_PTL_IP3_1|_RX|B2 0 _PTL_IP3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|6  2.685e-12
I_PTL_IP3_1|_RX|B3 0 _PTL_IP3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|9  2.764e-12
L_PTL_IP3_1|_RX|1 _PTL_IP3_1|A_PTL _PTL_IP3_1|_RX|1  1.346e-12
L_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|4  6.348e-12
L_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7  5.197e-12
L_PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7 IP3_1_OUT_RX  2.058e-12
L_PTL_IP3_1|_RX|P1 _PTL_IP3_1|_RX|2 0  4.795e-13
L_PTL_IP3_1|_RX|P2 _PTL_IP3_1|_RX|5 0  5.431e-13
L_PTL_IP3_1|_RX|P3 _PTL_IP3_1|_RX|8 0  5.339e-13
R_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|101  4.225701121488
R_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|104  3.429952209
R_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|107  2.7439617672
L_PTL_IP3_1|_RX|RB1 _PTL_IP3_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_1|_RX|RB2 _PTL_IP3_1|_RX|104 0  1.937922998085e-12
L_PTL_IP3_1|_RX|RB3 _PTL_IP3_1|_RX|107 0  1.550338398468e-12
LSPL_G1_1|SPL1|1 G1_1_RX SPL_G1_1|SPL1|D1  2e-12
LSPL_G1_1|SPL1|2 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|D2  4.135667696e-12
LSPL_G1_1|SPL1|3 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|JCT  9.84682784761905e-13
LSPL_G1_1|SPL1|4 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QA1  9.84682784761905e-13
LSPL_G1_1|SPL1|5 SPL_G1_1|SPL1|QA1 G1_1_TO1  2e-12
LSPL_G1_1|SPL1|6 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QB1  9.84682784761905e-13
LSPL_G1_1|SPL1|7 SPL_G1_1|SPL1|QB1 SPL_G1_1|QTMP  2e-12
LSPL_G1_1|SPL2|1 SPL_G1_1|QTMP SPL_G1_1|SPL2|D1  2e-12
LSPL_G1_1|SPL2|2 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|D2  4.135667696e-12
LSPL_G1_1|SPL2|3 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|JCT  9.84682784761905e-13
LSPL_G1_1|SPL2|4 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QA1  9.84682784761905e-13
LSPL_G1_1|SPL2|5 SPL_G1_1|SPL2|QA1 G1_1_TO2  2e-12
LSPL_G1_1|SPL2|6 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QB1  9.84682784761905e-13
LSPL_G1_1|SPL2|7 SPL_G1_1|SPL2|QB1 G1_1_TO3  2e-12
L_PG0_12|P|1 P0_1_RX _PG0_12|P|A1  2.067833848e-12
L_PG0_12|P|2 _PG0_12|P|A1 _PG0_12|P|A2  4.135667696e-12
L_PG0_12|P|3 _PG0_12|P|A3 _PG0_12|P|A4  8.271335392e-12
L_PG0_12|P|T T08 _PG0_12|P|T1  2.067833848e-12
L_PG0_12|P|4 _PG0_12|P|T1 _PG0_12|P|T2  4.135667696e-12
L_PG0_12|P|5 _PG0_12|P|A4 _PG0_12|P|Q1  4.135667696e-12
L_PG0_12|P|6 _PG0_12|P|Q1 P0_2  2.067833848e-12
L_PG0_12|G|1 G0_1_RX _PG0_12|G|A1  2.067833848e-12
L_PG0_12|G|2 _PG0_12|G|A1 _PG0_12|G|A2  4.135667696e-12
L_PG0_12|G|3 _PG0_12|G|A3 _PG0_12|G|A4  8.271335392e-12
L_PG0_12|G|T T08 _PG0_12|G|T1  2.067833848e-12
L_PG0_12|G|4 _PG0_12|G|T1 _PG0_12|G|T2  4.135667696e-12
L_PG0_12|G|5 _PG0_12|G|A4 _PG0_12|G|Q1  4.135667696e-12
L_PG0_12|G|6 _PG0_12|G|Q1 G0_2  2.067833848e-12
L_PG1_12|I_1|B _PG1_12|A1 _PG1_12|I_1|MID  2e-12
I_PG1_12|I_1|B 0 _PG1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_3|B _PG1_12|A3 _PG1_12|I_3|MID  2e-12
I_PG1_12|I_3|B 0 _PG1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_12|I_T|B _PG1_12|T1 _PG1_12|I_T|MID  2e-12
I_PG1_12|I_T|B 0 _PG1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_6|B _PG1_12|Q1 _PG1_12|I_6|MID  2e-12
I_PG1_12|I_6|B 0 _PG1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_12|1|1 _PG1_12|A1 _PG1_12|1|MID_SERIES JJMIT AREA=2.5
L_PG1_12|1|P _PG1_12|1|MID_SERIES 0  2e-13
R_PG1_12|1|B _PG1_12|A1 _PG1_12|1|MID_SHUNT  2.7439617672
L_PG1_12|1|RB _PG1_12|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|23|1 _PG1_12|A2 _PG1_12|A3 JJMIT AREA=1.7857142857142858
R_PG1_12|23|B _PG1_12|A2 _PG1_12|23|MID_SHUNT  3.84154647408
L_PG1_12|23|RB _PG1_12|23|MID_SHUNT _PG1_12|A3  2.1704737578552e-12
B_PG1_12|3|1 _PG1_12|A3 _PG1_12|3|MID_SERIES JJMIT AREA=2.5
L_PG1_12|3|P _PG1_12|3|MID_SERIES 0  2e-13
R_PG1_12|3|B _PG1_12|A3 _PG1_12|3|MID_SHUNT  2.7439617672
L_PG1_12|3|RB _PG1_12|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|4|1 _PG1_12|A4 _PG1_12|4|MID_SERIES JJMIT AREA=2.5
L_PG1_12|4|P _PG1_12|4|MID_SERIES 0  2e-13
R_PG1_12|4|B _PG1_12|A4 _PG1_12|4|MID_SHUNT  2.7439617672
L_PG1_12|4|RB _PG1_12|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|T|1 _PG1_12|T1 _PG1_12|T|MID_SERIES JJMIT AREA=2.5
L_PG1_12|T|P _PG1_12|T|MID_SERIES 0  2e-13
R_PG1_12|T|B _PG1_12|T1 _PG1_12|T|MID_SHUNT  2.7439617672
L_PG1_12|T|RB _PG1_12|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|45|1 _PG1_12|T2 _PG1_12|A4 JJMIT AREA=1.7857142857142858
R_PG1_12|45|B _PG1_12|T2 _PG1_12|45|MID_SHUNT  3.84154647408
L_PG1_12|45|RB _PG1_12|45|MID_SHUNT _PG1_12|A4  2.1704737578552e-12
B_PG1_12|6|1 _PG1_12|Q1 _PG1_12|6|MID_SERIES JJMIT AREA=2.5
L_PG1_12|6|P _PG1_12|6|MID_SERIES 0  2e-13
R_PG1_12|6|B _PG1_12|Q1 _PG1_12|6|MID_SHUNT  2.7439617672
L_PG1_12|6|RB _PG1_12|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|1 G2_1_RX _PG2_12|_SPL_G1|D1  2e-12
L_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|D2  4.135667696e-12
L_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG2_12|_SPL_G1|5 _PG2_12|_SPL_G1|QA1 _PG2_12|G1_COPY_1  2e-12
L_PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|QB1 _PG2_12|G1_COPY_2  2e-12
L_PG2_12|_PG|A1 P2_1_RX _PG2_12|_PG|A1  2.067833848e-12
L_PG2_12|_PG|A2 _PG2_12|_PG|A1 _PG2_12|_PG|A2  4.135667696e-12
L_PG2_12|_PG|A3 _PG2_12|_PG|A3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|B1 _PG2_12|G1_COPY_1 _PG2_12|_PG|B1  2.067833848e-12
L_PG2_12|_PG|B2 _PG2_12|_PG|B1 _PG2_12|_PG|B2  4.135667696e-12
L_PG2_12|_PG|B3 _PG2_12|_PG|B3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|Q3 _PG2_12|_PG|Q3 _PG2_12|_PG|Q2  4.135667696e-12
L_PG2_12|_PG|Q2 _PG2_12|_PG|Q2 _PG2_12|_PG|Q1  4.135667696e-12
L_PG2_12|_PG|Q1 _PG2_12|_PG|Q1 _PG2_12|PG  2.067833848e-12
L_PG2_12|_GG|A1 G1_1_TO2 _PG2_12|_GG|A1  2.067833848e-12
L_PG2_12|_GG|A2 _PG2_12|_GG|A1 _PG2_12|_GG|A2  4.135667696e-12
L_PG2_12|_GG|A3 _PG2_12|_GG|A3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|B1 _PG2_12|G1_COPY_2 _PG2_12|_GG|B1  2.067833848e-12
L_PG2_12|_GG|B2 _PG2_12|_GG|B1 _PG2_12|_GG|B2  4.135667696e-12
L_PG2_12|_GG|B3 _PG2_12|_GG|B3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|Q3 _PG2_12|_GG|Q3 _PG2_12|_GG|Q2  4.135667696e-12
L_PG2_12|_GG|Q2 _PG2_12|_GG|Q2 _PG2_12|_GG|Q1  4.135667696e-12
L_PG2_12|_GG|Q1 _PG2_12|_GG|Q1 _PG2_12|GG  2.067833848e-12
L_PG2_12|_DFF_PG|1 _PG2_12|PG _PG2_12|_DFF_PG|A1  2.067833848e-12
L_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|A2  4.135667696e-12
L_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|A4  8.271335392e-12
L_PG2_12|_DFF_PG|T T10 _PG2_12|_DFF_PG|T1  2.067833848e-12
L_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T2  4.135667696e-12
L_PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|Q1  4.135667696e-12
L_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|Q1 _PG2_12|PG_SYNC  2.067833848e-12
L_PG2_12|_DFF_GG|1 _PG2_12|GG _PG2_12|_DFF_GG|A1  2.067833848e-12
L_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|A2  4.135667696e-12
L_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|A4  8.271335392e-12
L_PG2_12|_DFF_GG|T T10 _PG2_12|_DFF_GG|T1  2.067833848e-12
L_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T2  4.135667696e-12
L_PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|Q1  4.135667696e-12
L_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|Q1 _PG2_12|GG_SYNC  2.067833848e-12
L_PG2_12|_AND_G|A1 _PG2_12|PG_SYNC _PG2_12|_AND_G|A1  2.067833848e-12
L_PG2_12|_AND_G|A2 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A2  4.135667696e-12
L_PG2_12|_AND_G|A3 _PG2_12|_AND_G|A3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|B1 _PG2_12|GG_SYNC _PG2_12|_AND_G|B1  2.067833848e-12
L_PG2_12|_AND_G|B2 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B2  4.135667696e-12
L_PG2_12|_AND_G|B3 _PG2_12|_AND_G|B3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q2  4.135667696e-12
L_PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q1  4.135667696e-12
L_PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1 G2_2  2.067833848e-12
L_PG3_12|_SPL_G1|1 G3_1_RX _PG3_12|_SPL_G1|D1  2e-12
L_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|D2  4.135667696e-12
L_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_12|_SPL_G1|5 _PG3_12|_SPL_G1|QA1 _PG3_12|G1_COPY_1  2e-12
L_PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|QB1 _PG3_12|G1_COPY_2  2e-12
L_PG3_12|_PG|A1 P3_1_RX _PG3_12|_PG|A1  2.067833848e-12
L_PG3_12|_PG|A2 _PG3_12|_PG|A1 _PG3_12|_PG|A2  4.135667696e-12
L_PG3_12|_PG|A3 _PG3_12|_PG|A3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|B1 _PG3_12|G1_COPY_1 _PG3_12|_PG|B1  2.067833848e-12
L_PG3_12|_PG|B2 _PG3_12|_PG|B1 _PG3_12|_PG|B2  4.135667696e-12
L_PG3_12|_PG|B3 _PG3_12|_PG|B3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|Q3 _PG3_12|_PG|Q3 _PG3_12|_PG|Q2  4.135667696e-12
L_PG3_12|_PG|Q2 _PG3_12|_PG|Q2 _PG3_12|_PG|Q1  4.135667696e-12
L_PG3_12|_PG|Q1 _PG3_12|_PG|Q1 _PG3_12|PG  2.067833848e-12
L_PG3_12|_GG|A1 G1_1_TO3 _PG3_12|_GG|A1  2.067833848e-12
L_PG3_12|_GG|A2 _PG3_12|_GG|A1 _PG3_12|_GG|A2  4.135667696e-12
L_PG3_12|_GG|A3 _PG3_12|_GG|A3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|B1 _PG3_12|G1_COPY_2 _PG3_12|_GG|B1  2.067833848e-12
L_PG3_12|_GG|B2 _PG3_12|_GG|B1 _PG3_12|_GG|B2  4.135667696e-12
L_PG3_12|_GG|B3 _PG3_12|_GG|B3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|Q3 _PG3_12|_GG|Q3 _PG3_12|_GG|Q2  4.135667696e-12
L_PG3_12|_GG|Q2 _PG3_12|_GG|Q2 _PG3_12|_GG|Q1  4.135667696e-12
L_PG3_12|_GG|Q1 _PG3_12|_GG|Q1 _PG3_12|GG  2.067833848e-12
L_PG3_12|_DFF_PG|1 _PG3_12|PG _PG3_12|_DFF_PG|A1  2.067833848e-12
L_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|A2  4.135667696e-12
L_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|A4  8.271335392e-12
L_PG3_12|_DFF_PG|T T11 _PG3_12|_DFF_PG|T1  2.067833848e-12
L_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T2  4.135667696e-12
L_PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|Q1  4.135667696e-12
L_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|Q1 _PG3_12|PG_SYNC  2.067833848e-12
L_PG3_12|_DFF_GG|1 _PG3_12|GG _PG3_12|_DFF_GG|A1  2.067833848e-12
L_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|A2  4.135667696e-12
L_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|A4  8.271335392e-12
L_PG3_12|_DFF_GG|T T11 _PG3_12|_DFF_GG|T1  2.067833848e-12
L_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T2  4.135667696e-12
L_PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|Q1  4.135667696e-12
L_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|Q1 _PG3_12|GG_SYNC  2.067833848e-12
L_PG3_12|_AND_G|A1 _PG3_12|PG_SYNC _PG3_12|_AND_G|A1  2.067833848e-12
L_PG3_12|_AND_G|A2 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A2  4.135667696e-12
L_PG3_12|_AND_G|A3 _PG3_12|_AND_G|A3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|B1 _PG3_12|GG_SYNC _PG3_12|_AND_G|B1  2.067833848e-12
L_PG3_12|_AND_G|B2 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B2  4.135667696e-12
L_PG3_12|_AND_G|B3 _PG3_12|_AND_G|B3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q2  4.135667696e-12
L_PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q1  4.135667696e-12
L_PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1 G3_2  2.067833848e-12
L_DFF_IP1_12|I_1|B _DFF_IP1_12|A1 _DFF_IP1_12|I_1|MID  2e-12
I_DFF_IP1_12|I_1|B 0 _DFF_IP1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_3|B _DFF_IP1_12|A3 _DFF_IP1_12|I_3|MID  2e-12
I_DFF_IP1_12|I_3|B 0 _DFF_IP1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_12|I_T|B _DFF_IP1_12|T1 _DFF_IP1_12|I_T|MID  2e-12
I_DFF_IP1_12|I_T|B 0 _DFF_IP1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_6|B _DFF_IP1_12|Q1 _DFF_IP1_12|I_6|MID  2e-12
I_DFF_IP1_12|I_6|B 0 _DFF_IP1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_12|1|1 _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|1|P _DFF_IP1_12|1|MID_SERIES 0  2e-13
R_DFF_IP1_12|1|B _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SHUNT  2.7439617672
L_DFF_IP1_12|1|RB _DFF_IP1_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|23|1 _DFF_IP1_12|A2 _DFF_IP1_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|23|B _DFF_IP1_12|A2 _DFF_IP1_12|23|MID_SHUNT  3.84154647408
L_DFF_IP1_12|23|RB _DFF_IP1_12|23|MID_SHUNT _DFF_IP1_12|A3  2.1704737578552e-12
B_DFF_IP1_12|3|1 _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|3|P _DFF_IP1_12|3|MID_SERIES 0  2e-13
R_DFF_IP1_12|3|B _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SHUNT  2.7439617672
L_DFF_IP1_12|3|RB _DFF_IP1_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|4|1 _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|4|P _DFF_IP1_12|4|MID_SERIES 0  2e-13
R_DFF_IP1_12|4|B _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SHUNT  2.7439617672
L_DFF_IP1_12|4|RB _DFF_IP1_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|T|1 _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|T|P _DFF_IP1_12|T|MID_SERIES 0  2e-13
R_DFF_IP1_12|T|B _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SHUNT  2.7439617672
L_DFF_IP1_12|T|RB _DFF_IP1_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|45|1 _DFF_IP1_12|T2 _DFF_IP1_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|45|B _DFF_IP1_12|T2 _DFF_IP1_12|45|MID_SHUNT  3.84154647408
L_DFF_IP1_12|45|RB _DFF_IP1_12|45|MID_SHUNT _DFF_IP1_12|A4  2.1704737578552e-12
B_DFF_IP1_12|6|1 _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|6|P _DFF_IP1_12|6|MID_SERIES 0  2e-13
R_DFF_IP1_12|6|B _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SHUNT  2.7439617672
L_DFF_IP1_12|6|RB _DFF_IP1_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_12|I_1|B _DFF_IP2_12|A1 _DFF_IP2_12|I_1|MID  2e-12
I_DFF_IP2_12|I_1|B 0 _DFF_IP2_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_3|B _DFF_IP2_12|A3 _DFF_IP2_12|I_3|MID  2e-12
I_DFF_IP2_12|I_3|B 0 _DFF_IP2_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_12|I_T|B _DFF_IP2_12|T1 _DFF_IP2_12|I_T|MID  2e-12
I_DFF_IP2_12|I_T|B 0 _DFF_IP2_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_6|B _DFF_IP2_12|Q1 _DFF_IP2_12|I_6|MID  2e-12
I_DFF_IP2_12|I_6|B 0 _DFF_IP2_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_12|1|1 _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|1|P _DFF_IP2_12|1|MID_SERIES 0  2e-13
R_DFF_IP2_12|1|B _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SHUNT  2.7439617672
L_DFF_IP2_12|1|RB _DFF_IP2_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|23|1 _DFF_IP2_12|A2 _DFF_IP2_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|23|B _DFF_IP2_12|A2 _DFF_IP2_12|23|MID_SHUNT  3.84154647408
L_DFF_IP2_12|23|RB _DFF_IP2_12|23|MID_SHUNT _DFF_IP2_12|A3  2.1704737578552e-12
B_DFF_IP2_12|3|1 _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|3|P _DFF_IP2_12|3|MID_SERIES 0  2e-13
R_DFF_IP2_12|3|B _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SHUNT  2.7439617672
L_DFF_IP2_12|3|RB _DFF_IP2_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|4|1 _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|4|P _DFF_IP2_12|4|MID_SERIES 0  2e-13
R_DFF_IP2_12|4|B _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SHUNT  2.7439617672
L_DFF_IP2_12|4|RB _DFF_IP2_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|T|1 _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|T|P _DFF_IP2_12|T|MID_SERIES 0  2e-13
R_DFF_IP2_12|T|B _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SHUNT  2.7439617672
L_DFF_IP2_12|T|RB _DFF_IP2_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|45|1 _DFF_IP2_12|T2 _DFF_IP2_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|45|B _DFF_IP2_12|T2 _DFF_IP2_12|45|MID_SHUNT  3.84154647408
L_DFF_IP2_12|45|RB _DFF_IP2_12|45|MID_SHUNT _DFF_IP2_12|A4  2.1704737578552e-12
B_DFF_IP2_12|6|1 _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|6|P _DFF_IP2_12|6|MID_SERIES 0  2e-13
R_DFF_IP2_12|6|B _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SHUNT  2.7439617672
L_DFF_IP2_12|6|RB _DFF_IP2_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_12|I_1|B _DFF_IP3_12|A1 _DFF_IP3_12|I_1|MID  2e-12
I_DFF_IP3_12|I_1|B 0 _DFF_IP3_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_3|B _DFF_IP3_12|A3 _DFF_IP3_12|I_3|MID  2e-12
I_DFF_IP3_12|I_3|B 0 _DFF_IP3_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_12|I_T|B _DFF_IP3_12|T1 _DFF_IP3_12|I_T|MID  2e-12
I_DFF_IP3_12|I_T|B 0 _DFF_IP3_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_6|B _DFF_IP3_12|Q1 _DFF_IP3_12|I_6|MID  2e-12
I_DFF_IP3_12|I_6|B 0 _DFF_IP3_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_12|1|1 _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|1|P _DFF_IP3_12|1|MID_SERIES 0  2e-13
R_DFF_IP3_12|1|B _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SHUNT  2.7439617672
L_DFF_IP3_12|1|RB _DFF_IP3_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|23|1 _DFF_IP3_12|A2 _DFF_IP3_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|23|B _DFF_IP3_12|A2 _DFF_IP3_12|23|MID_SHUNT  3.84154647408
L_DFF_IP3_12|23|RB _DFF_IP3_12|23|MID_SHUNT _DFF_IP3_12|A3  2.1704737578552e-12
B_DFF_IP3_12|3|1 _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|3|P _DFF_IP3_12|3|MID_SERIES 0  2e-13
R_DFF_IP3_12|3|B _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SHUNT  2.7439617672
L_DFF_IP3_12|3|RB _DFF_IP3_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|4|1 _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|4|P _DFF_IP3_12|4|MID_SERIES 0  2e-13
R_DFF_IP3_12|4|B _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SHUNT  2.7439617672
L_DFF_IP3_12|4|RB _DFF_IP3_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|T|1 _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|T|P _DFF_IP3_12|T|MID_SERIES 0  2e-13
R_DFF_IP3_12|T|B _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SHUNT  2.7439617672
L_DFF_IP3_12|T|RB _DFF_IP3_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|45|1 _DFF_IP3_12|T2 _DFF_IP3_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|45|B _DFF_IP3_12|T2 _DFF_IP3_12|45|MID_SHUNT  3.84154647408
L_DFF_IP3_12|45|RB _DFF_IP3_12|45|MID_SHUNT _DFF_IP3_12|A4  2.1704737578552e-12
B_DFF_IP3_12|6|1 _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|6|P _DFF_IP3_12|6|MID_SERIES 0  2e-13
R_DFF_IP3_12|6|B _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SHUNT  2.7439617672
L_DFF_IP3_12|6|RB _DFF_IP3_12|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_P0_2|_TX|1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|2 JJMIT AREA=2.5
B_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|5 JJMIT AREA=2.5
I_PTL_P0_2|_TX|B1 0 _PTL_P0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_2|_TX|B2 0 _PTL_P0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|3  1.684e-12
L_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|6  3.596e-12
L_PTL_P0_2|_TX|1 P0_2 _PTL_P0_2|_TX|1  2.063e-12
L_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|4  4.123e-12
L_PTL_P0_2|_TX|3 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|7  2.193e-12
R_PTL_P0_2|_TX|D _PTL_P0_2|_TX|7 _PTL_P0_2|A_PTL  1.36
L_PTL_P0_2|_TX|P1 _PTL_P0_2|_TX|2 0  5.254e-13
L_PTL_P0_2|_TX|P2 _PTL_P0_2|_TX|5 0  5.141e-13
R_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|101  2.7439617672
R_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|104  2.7439617672
L_PTL_P0_2|_TX|RB1 _PTL_P0_2|_TX|101 0  1.550338398468e-12
L_PTL_P0_2|_TX|RB2 _PTL_P0_2|_TX|104 0  1.550338398468e-12
B_PTL_P0_2|_RX|1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|5 JJMIT AREA=2.0
B_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|8 JJMIT AREA=2.5
I_PTL_P0_2|_RX|B1 0 _PTL_P0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|3  2.777e-12
I_PTL_P0_2|_RX|B2 0 _PTL_P0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|6  2.685e-12
I_PTL_P0_2|_RX|B3 0 _PTL_P0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|9  2.764e-12
L_PTL_P0_2|_RX|1 _PTL_P0_2|A_PTL _PTL_P0_2|_RX|1  1.346e-12
L_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|4  6.348e-12
L_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7  5.197e-12
L_PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7 _PTL_P0_2|A_PTL_RX  2.058e-12
L_PTL_P0_2|_RX|P1 _PTL_P0_2|_RX|2 0  4.795e-13
L_PTL_P0_2|_RX|P2 _PTL_P0_2|_RX|5 0  5.431e-13
L_PTL_P0_2|_RX|P3 _PTL_P0_2|_RX|8 0  5.339e-13
R_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|101  4.225701121488
R_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|104  3.429952209
R_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|107  2.7439617672
L_PTL_P0_2|_RX|RB1 _PTL_P0_2|_RX|101 0  2.38752113364072e-12
L_PTL_P0_2|_RX|RB2 _PTL_P0_2|_RX|104 0  1.937922998085e-12
L_PTL_P0_2|_RX|RB3 _PTL_P0_2|_RX|107 0  1.550338398468e-12
B_PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|2 JJMIT AREA=2.5
B_PTL_P0_2|_JTL|2 _PTL_P0_2|_JTL|6 _PTL_P0_2|_JTL|7 JJMIT AREA=2.5
I_PTL_P0_2|_JTL|B1 0 _PTL_P0_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_P0_2|_JTL|1 _PTL_P0_2|A_PTL_RX _PTL_P0_2|_JTL|1  2.067833848e-12
L_PTL_P0_2|_JTL|2 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|4  2.067833848e-12
L_PTL_P0_2|_JTL|3 _PTL_P0_2|_JTL|4 _PTL_P0_2|_JTL|6  2.067833848e-12
L_PTL_P0_2|_JTL|4 _PTL_P0_2|_JTL|6 P0_2_RX  2.067833848e-12
L_PTL_P0_2|_JTL|P1 _PTL_P0_2|_JTL|2 0  2e-13
L_PTL_P0_2|_JTL|P2 _PTL_P0_2|_JTL|7 0  2e-13
L_PTL_P0_2|_JTL|B1 _PTL_P0_2|_JTL|5 _PTL_P0_2|_JTL|4  2e-12
R_PTL_P0_2|_JTL|B1 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|3  2.7439617672
R_PTL_P0_2|_JTL|B2 _PTL_P0_2|_JTL|6 _PTL_P0_2|_JTL|8  2.7439617672
L_PTL_P0_2|_JTL|RB1 _PTL_P0_2|_JTL|3 0  1.750338398468e-12
L_PTL_P0_2|_JTL|RB2 _PTL_P0_2|_JTL|8 0  1.750338398468e-12
B_PTL_G0_2|_TX|1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|2 JJMIT AREA=2.5
B_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|5 JJMIT AREA=2.5
I_PTL_G0_2|_TX|B1 0 _PTL_G0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_2|_TX|B2 0 _PTL_G0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|3  1.684e-12
L_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|6  3.596e-12
L_PTL_G0_2|_TX|1 G0_2 _PTL_G0_2|_TX|1  2.063e-12
L_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|4  4.123e-12
L_PTL_G0_2|_TX|3 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|7  2.193e-12
R_PTL_G0_2|_TX|D _PTL_G0_2|_TX|7 _PTL_G0_2|A_PTL  1.36
L_PTL_G0_2|_TX|P1 _PTL_G0_2|_TX|2 0  5.254e-13
L_PTL_G0_2|_TX|P2 _PTL_G0_2|_TX|5 0  5.141e-13
R_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|101  2.7439617672
R_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|104  2.7439617672
L_PTL_G0_2|_TX|RB1 _PTL_G0_2|_TX|101 0  1.550338398468e-12
L_PTL_G0_2|_TX|RB2 _PTL_G0_2|_TX|104 0  1.550338398468e-12
B_PTL_G0_2|_RX|1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|5 JJMIT AREA=2.0
B_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|8 JJMIT AREA=2.5
I_PTL_G0_2|_RX|B1 0 _PTL_G0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|3  2.777e-12
I_PTL_G0_2|_RX|B2 0 _PTL_G0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|6  2.685e-12
I_PTL_G0_2|_RX|B3 0 _PTL_G0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|9  2.764e-12
L_PTL_G0_2|_RX|1 _PTL_G0_2|A_PTL _PTL_G0_2|_RX|1  1.346e-12
L_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|4  6.348e-12
L_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7  5.197e-12
L_PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7 _PTL_G0_2|A_PTL_RX  2.058e-12
L_PTL_G0_2|_RX|P1 _PTL_G0_2|_RX|2 0  4.795e-13
L_PTL_G0_2|_RX|P2 _PTL_G0_2|_RX|5 0  5.431e-13
L_PTL_G0_2|_RX|P3 _PTL_G0_2|_RX|8 0  5.339e-13
R_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|101  4.225701121488
R_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|104  3.429952209
R_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|107  2.7439617672
L_PTL_G0_2|_RX|RB1 _PTL_G0_2|_RX|101 0  2.38752113364072e-12
L_PTL_G0_2|_RX|RB2 _PTL_G0_2|_RX|104 0  1.937922998085e-12
L_PTL_G0_2|_RX|RB3 _PTL_G0_2|_RX|107 0  1.550338398468e-12
B_PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G0_2|_JTL|2 _PTL_G0_2|_JTL|6 _PTL_G0_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G0_2|_JTL|B1 0 _PTL_G0_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G0_2|_JTL|1 _PTL_G0_2|A_PTL_RX _PTL_G0_2|_JTL|1  2.067833848e-12
L_PTL_G0_2|_JTL|2 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|4  2.067833848e-12
L_PTL_G0_2|_JTL|3 _PTL_G0_2|_JTL|4 _PTL_G0_2|_JTL|6  2.067833848e-12
L_PTL_G0_2|_JTL|4 _PTL_G0_2|_JTL|6 G0_2_RX  2.067833848e-12
L_PTL_G0_2|_JTL|P1 _PTL_G0_2|_JTL|2 0  2e-13
L_PTL_G0_2|_JTL|P2 _PTL_G0_2|_JTL|7 0  2e-13
L_PTL_G0_2|_JTL|B1 _PTL_G0_2|_JTL|5 _PTL_G0_2|_JTL|4  2e-12
R_PTL_G0_2|_JTL|B1 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|3  2.7439617672
R_PTL_G0_2|_JTL|B2 _PTL_G0_2|_JTL|6 _PTL_G0_2|_JTL|8  2.7439617672
L_PTL_G0_2|_JTL|RB1 _PTL_G0_2|_JTL|3 0  1.750338398468e-12
L_PTL_G0_2|_JTL|RB2 _PTL_G0_2|_JTL|8 0  1.750338398468e-12
B_PTL_G1_2|_TX|1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|2 JJMIT AREA=2.5
B_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|5 JJMIT AREA=2.5
I_PTL_G1_2|_TX|B1 0 _PTL_G1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_2|_TX|B2 0 _PTL_G1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|3  1.684e-12
L_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|6  3.596e-12
L_PTL_G1_2|_TX|1 G1_2 _PTL_G1_2|_TX|1  2.063e-12
L_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|4  4.123e-12
L_PTL_G1_2|_TX|3 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|7  2.193e-12
R_PTL_G1_2|_TX|D _PTL_G1_2|_TX|7 _PTL_G1_2|A_PTL  1.36
L_PTL_G1_2|_TX|P1 _PTL_G1_2|_TX|2 0  5.254e-13
L_PTL_G1_2|_TX|P2 _PTL_G1_2|_TX|5 0  5.141e-13
R_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|101  2.7439617672
R_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|104  2.7439617672
L_PTL_G1_2|_TX|RB1 _PTL_G1_2|_TX|101 0  1.550338398468e-12
L_PTL_G1_2|_TX|RB2 _PTL_G1_2|_TX|104 0  1.550338398468e-12
B_PTL_G1_2|_RX|1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|5 JJMIT AREA=2.0
B_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|8 JJMIT AREA=2.5
I_PTL_G1_2|_RX|B1 0 _PTL_G1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|3  2.777e-12
I_PTL_G1_2|_RX|B2 0 _PTL_G1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|6  2.685e-12
I_PTL_G1_2|_RX|B3 0 _PTL_G1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|9  2.764e-12
L_PTL_G1_2|_RX|1 _PTL_G1_2|A_PTL _PTL_G1_2|_RX|1  1.346e-12
L_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|4  6.348e-12
L_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7  5.197e-12
L_PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7 _PTL_G1_2|A_PTL_RX  2.058e-12
L_PTL_G1_2|_RX|P1 _PTL_G1_2|_RX|2 0  4.795e-13
L_PTL_G1_2|_RX|P2 _PTL_G1_2|_RX|5 0  5.431e-13
L_PTL_G1_2|_RX|P3 _PTL_G1_2|_RX|8 0  5.339e-13
R_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|101  4.225701121488
R_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|104  3.429952209
R_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|107  2.7439617672
L_PTL_G1_2|_RX|RB1 _PTL_G1_2|_RX|101 0  2.38752113364072e-12
L_PTL_G1_2|_RX|RB2 _PTL_G1_2|_RX|104 0  1.937922998085e-12
L_PTL_G1_2|_RX|RB3 _PTL_G1_2|_RX|107 0  1.550338398468e-12
B_PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G1_2|_JTL|2 _PTL_G1_2|_JTL|6 _PTL_G1_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G1_2|_JTL|B1 0 _PTL_G1_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G1_2|_JTL|1 _PTL_G1_2|A_PTL_RX _PTL_G1_2|_JTL|1  2.067833848e-12
L_PTL_G1_2|_JTL|2 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|4  2.067833848e-12
L_PTL_G1_2|_JTL|3 _PTL_G1_2|_JTL|4 _PTL_G1_2|_JTL|6  2.067833848e-12
L_PTL_G1_2|_JTL|4 _PTL_G1_2|_JTL|6 G1_2_RX  2.067833848e-12
L_PTL_G1_2|_JTL|P1 _PTL_G1_2|_JTL|2 0  2e-13
L_PTL_G1_2|_JTL|P2 _PTL_G1_2|_JTL|7 0  2e-13
L_PTL_G1_2|_JTL|B1 _PTL_G1_2|_JTL|5 _PTL_G1_2|_JTL|4  2e-12
R_PTL_G1_2|_JTL|B1 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|3  2.7439617672
R_PTL_G1_2|_JTL|B2 _PTL_G1_2|_JTL|6 _PTL_G1_2|_JTL|8  2.7439617672
L_PTL_G1_2|_JTL|RB1 _PTL_G1_2|_JTL|3 0  1.750338398468e-12
L_PTL_G1_2|_JTL|RB2 _PTL_G1_2|_JTL|8 0  1.750338398468e-12
B_PTL_G2_2|_TX|1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|2 JJMIT AREA=2.5
B_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|5 JJMIT AREA=2.5
I_PTL_G2_2|_TX|B1 0 _PTL_G2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_2|_TX|B2 0 _PTL_G2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|3  1.684e-12
L_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|6  3.596e-12
L_PTL_G2_2|_TX|1 G2_2 _PTL_G2_2|_TX|1  2.063e-12
L_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|4  4.123e-12
L_PTL_G2_2|_TX|3 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|7  2.193e-12
R_PTL_G2_2|_TX|D _PTL_G2_2|_TX|7 _PTL_G2_2|A_PTL  1.36
L_PTL_G2_2|_TX|P1 _PTL_G2_2|_TX|2 0  5.254e-13
L_PTL_G2_2|_TX|P2 _PTL_G2_2|_TX|5 0  5.141e-13
R_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|101  2.7439617672
R_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|104  2.7439617672
L_PTL_G2_2|_TX|RB1 _PTL_G2_2|_TX|101 0  1.550338398468e-12
L_PTL_G2_2|_TX|RB2 _PTL_G2_2|_TX|104 0  1.550338398468e-12
B_PTL_G2_2|_RX|1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|5 JJMIT AREA=2.0
B_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|8 JJMIT AREA=2.5
I_PTL_G2_2|_RX|B1 0 _PTL_G2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|3  2.777e-12
I_PTL_G2_2|_RX|B2 0 _PTL_G2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|6  2.685e-12
I_PTL_G2_2|_RX|B3 0 _PTL_G2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|9  2.764e-12
L_PTL_G2_2|_RX|1 _PTL_G2_2|A_PTL _PTL_G2_2|_RX|1  1.346e-12
L_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|4  6.348e-12
L_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7  5.197e-12
L_PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7 _PTL_G2_2|A_PTL_RX  2.058e-12
L_PTL_G2_2|_RX|P1 _PTL_G2_2|_RX|2 0  4.795e-13
L_PTL_G2_2|_RX|P2 _PTL_G2_2|_RX|5 0  5.431e-13
L_PTL_G2_2|_RX|P3 _PTL_G2_2|_RX|8 0  5.339e-13
R_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|101  4.225701121488
R_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|104  3.429952209
R_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|107  2.7439617672
L_PTL_G2_2|_RX|RB1 _PTL_G2_2|_RX|101 0  2.38752113364072e-12
L_PTL_G2_2|_RX|RB2 _PTL_G2_2|_RX|104 0  1.937922998085e-12
L_PTL_G2_2|_RX|RB3 _PTL_G2_2|_RX|107 0  1.550338398468e-12
B_PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G2_2|_JTL|2 _PTL_G2_2|_JTL|6 _PTL_G2_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G2_2|_JTL|B1 0 _PTL_G2_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G2_2|_JTL|1 _PTL_G2_2|A_PTL_RX _PTL_G2_2|_JTL|1  2.067833848e-12
L_PTL_G2_2|_JTL|2 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|4  2.067833848e-12
L_PTL_G2_2|_JTL|3 _PTL_G2_2|_JTL|4 _PTL_G2_2|_JTL|6  2.067833848e-12
L_PTL_G2_2|_JTL|4 _PTL_G2_2|_JTL|6 G2_2_RX  2.067833848e-12
L_PTL_G2_2|_JTL|P1 _PTL_G2_2|_JTL|2 0  2e-13
L_PTL_G2_2|_JTL|P2 _PTL_G2_2|_JTL|7 0  2e-13
L_PTL_G2_2|_JTL|B1 _PTL_G2_2|_JTL|5 _PTL_G2_2|_JTL|4  2e-12
R_PTL_G2_2|_JTL|B1 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|3  2.7439617672
R_PTL_G2_2|_JTL|B2 _PTL_G2_2|_JTL|6 _PTL_G2_2|_JTL|8  2.7439617672
L_PTL_G2_2|_JTL|RB1 _PTL_G2_2|_JTL|3 0  1.750338398468e-12
L_PTL_G2_2|_JTL|RB2 _PTL_G2_2|_JTL|8 0  1.750338398468e-12
B_PTL_G3_2|_TX|1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|2 JJMIT AREA=2.5
B_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|5 JJMIT AREA=2.5
I_PTL_G3_2|_TX|B1 0 _PTL_G3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_2|_TX|B2 0 _PTL_G3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|3  1.684e-12
L_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|6  3.596e-12
L_PTL_G3_2|_TX|1 G3_2 _PTL_G3_2|_TX|1  2.063e-12
L_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|4  4.123e-12
L_PTL_G3_2|_TX|3 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|7  2.193e-12
R_PTL_G3_2|_TX|D _PTL_G3_2|_TX|7 _PTL_G3_2|A_PTL  1.36
L_PTL_G3_2|_TX|P1 _PTL_G3_2|_TX|2 0  5.254e-13
L_PTL_G3_2|_TX|P2 _PTL_G3_2|_TX|5 0  5.141e-13
R_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|101  2.7439617672
R_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|104  2.7439617672
L_PTL_G3_2|_TX|RB1 _PTL_G3_2|_TX|101 0  1.550338398468e-12
L_PTL_G3_2|_TX|RB2 _PTL_G3_2|_TX|104 0  1.550338398468e-12
B_PTL_G3_2|_RX|1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|5 JJMIT AREA=2.0
B_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|8 JJMIT AREA=2.5
I_PTL_G3_2|_RX|B1 0 _PTL_G3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|3  2.777e-12
I_PTL_G3_2|_RX|B2 0 _PTL_G3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|6  2.685e-12
I_PTL_G3_2|_RX|B3 0 _PTL_G3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|9  2.764e-12
L_PTL_G3_2|_RX|1 _PTL_G3_2|A_PTL _PTL_G3_2|_RX|1  1.346e-12
L_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|4  6.348e-12
L_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7  5.197e-12
L_PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7 _PTL_G3_2|A_PTL_RX  2.058e-12
L_PTL_G3_2|_RX|P1 _PTL_G3_2|_RX|2 0  4.795e-13
L_PTL_G3_2|_RX|P2 _PTL_G3_2|_RX|5 0  5.431e-13
L_PTL_G3_2|_RX|P3 _PTL_G3_2|_RX|8 0  5.339e-13
R_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|101  4.225701121488
R_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|104  3.429952209
R_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|107  2.7439617672
L_PTL_G3_2|_RX|RB1 _PTL_G3_2|_RX|101 0  2.38752113364072e-12
L_PTL_G3_2|_RX|RB2 _PTL_G3_2|_RX|104 0  1.937922998085e-12
L_PTL_G3_2|_RX|RB3 _PTL_G3_2|_RX|107 0  1.550338398468e-12
B_PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G3_2|_JTL|2 _PTL_G3_2|_JTL|6 _PTL_G3_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G3_2|_JTL|B1 0 _PTL_G3_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G3_2|_JTL|1 _PTL_G3_2|A_PTL_RX _PTL_G3_2|_JTL|1  2.067833848e-12
L_PTL_G3_2|_JTL|2 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|4  2.067833848e-12
L_PTL_G3_2|_JTL|3 _PTL_G3_2|_JTL|4 _PTL_G3_2|_JTL|6  2.067833848e-12
L_PTL_G3_2|_JTL|4 _PTL_G3_2|_JTL|6 G3_2_RX  2.067833848e-12
L_PTL_G3_2|_JTL|P1 _PTL_G3_2|_JTL|2 0  2e-13
L_PTL_G3_2|_JTL|P2 _PTL_G3_2|_JTL|7 0  2e-13
L_PTL_G3_2|_JTL|B1 _PTL_G3_2|_JTL|5 _PTL_G3_2|_JTL|4  2e-12
R_PTL_G3_2|_JTL|B1 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|3  2.7439617672
R_PTL_G3_2|_JTL|B2 _PTL_G3_2|_JTL|6 _PTL_G3_2|_JTL|8  2.7439617672
L_PTL_G3_2|_JTL|RB1 _PTL_G3_2|_JTL|3 0  1.750338398468e-12
L_PTL_G3_2|_JTL|RB2 _PTL_G3_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_2|_TX|B1 0 _PTL_IP1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_2|_TX|B2 0 _PTL_IP1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|3  1.684e-12
L_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|6  3.596e-12
L_PTL_IP1_2|_TX|1 IP1_2_OUT _PTL_IP1_2|_TX|1  2.063e-12
L_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|4  4.123e-12
L_PTL_IP1_2|_TX|3 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|7  2.193e-12
R_PTL_IP1_2|_TX|D _PTL_IP1_2|_TX|7 _PTL_IP1_2|A_PTL  1.36
L_PTL_IP1_2|_TX|P1 _PTL_IP1_2|_TX|2 0  5.254e-13
L_PTL_IP1_2|_TX|P2 _PTL_IP1_2|_TX|5 0  5.141e-13
R_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|101  2.7439617672
R_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|104  2.7439617672
L_PTL_IP1_2|_TX|RB1 _PTL_IP1_2|_TX|101 0  1.550338398468e-12
L_PTL_IP1_2|_TX|RB2 _PTL_IP1_2|_TX|104 0  1.550338398468e-12
B_PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_2|_RX|B1 0 _PTL_IP1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|3  2.777e-12
I_PTL_IP1_2|_RX|B2 0 _PTL_IP1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|6  2.685e-12
I_PTL_IP1_2|_RX|B3 0 _PTL_IP1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|9  2.764e-12
L_PTL_IP1_2|_RX|1 _PTL_IP1_2|A_PTL _PTL_IP1_2|_RX|1  1.346e-12
L_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|4  6.348e-12
L_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7  5.197e-12
L_PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7 _PTL_IP1_2|A_PTL_RX  2.058e-12
L_PTL_IP1_2|_RX|P1 _PTL_IP1_2|_RX|2 0  4.795e-13
L_PTL_IP1_2|_RX|P2 _PTL_IP1_2|_RX|5 0  5.431e-13
L_PTL_IP1_2|_RX|P3 _PTL_IP1_2|_RX|8 0  5.339e-13
R_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|101  4.225701121488
R_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|104  3.429952209
R_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|107  2.7439617672
L_PTL_IP1_2|_RX|RB1 _PTL_IP1_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_2|_RX|RB2 _PTL_IP1_2|_RX|104 0  1.937922998085e-12
L_PTL_IP1_2|_RX|RB3 _PTL_IP1_2|_RX|107 0  1.550338398468e-12
B_PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP1_2|_JTL|2 _PTL_IP1_2|_JTL|6 _PTL_IP1_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP1_2|_JTL|B1 0 _PTL_IP1_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP1_2|_JTL|1 _PTL_IP1_2|A_PTL_RX _PTL_IP1_2|_JTL|1  2.067833848e-12
L_PTL_IP1_2|_JTL|2 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|4  2.067833848e-12
L_PTL_IP1_2|_JTL|3 _PTL_IP1_2|_JTL|4 _PTL_IP1_2|_JTL|6  2.067833848e-12
L_PTL_IP1_2|_JTL|4 _PTL_IP1_2|_JTL|6 IP1_2_OUT_RX  2.067833848e-12
L_PTL_IP1_2|_JTL|P1 _PTL_IP1_2|_JTL|2 0  2e-13
L_PTL_IP1_2|_JTL|P2 _PTL_IP1_2|_JTL|7 0  2e-13
L_PTL_IP1_2|_JTL|B1 _PTL_IP1_2|_JTL|5 _PTL_IP1_2|_JTL|4  2e-12
R_PTL_IP1_2|_JTL|B1 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|3  2.7439617672
R_PTL_IP1_2|_JTL|B2 _PTL_IP1_2|_JTL|6 _PTL_IP1_2|_JTL|8  2.7439617672
L_PTL_IP1_2|_JTL|RB1 _PTL_IP1_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP1_2|_JTL|RB2 _PTL_IP1_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_2|_TX|B1 0 _PTL_IP2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_2|_TX|B2 0 _PTL_IP2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|3  1.684e-12
L_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|6  3.596e-12
L_PTL_IP2_2|_TX|1 IP2_2_OUT _PTL_IP2_2|_TX|1  2.063e-12
L_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|4  4.123e-12
L_PTL_IP2_2|_TX|3 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|7  2.193e-12
R_PTL_IP2_2|_TX|D _PTL_IP2_2|_TX|7 _PTL_IP2_2|A_PTL  1.36
L_PTL_IP2_2|_TX|P1 _PTL_IP2_2|_TX|2 0  5.254e-13
L_PTL_IP2_2|_TX|P2 _PTL_IP2_2|_TX|5 0  5.141e-13
R_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|101  2.7439617672
R_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|104  2.7439617672
L_PTL_IP2_2|_TX|RB1 _PTL_IP2_2|_TX|101 0  1.550338398468e-12
L_PTL_IP2_2|_TX|RB2 _PTL_IP2_2|_TX|104 0  1.550338398468e-12
B_PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_2|_RX|B1 0 _PTL_IP2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|3  2.777e-12
I_PTL_IP2_2|_RX|B2 0 _PTL_IP2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|6  2.685e-12
I_PTL_IP2_2|_RX|B3 0 _PTL_IP2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|9  2.764e-12
L_PTL_IP2_2|_RX|1 _PTL_IP2_2|A_PTL _PTL_IP2_2|_RX|1  1.346e-12
L_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|4  6.348e-12
L_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7  5.197e-12
L_PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7 _PTL_IP2_2|A_PTL_RX  2.058e-12
L_PTL_IP2_2|_RX|P1 _PTL_IP2_2|_RX|2 0  4.795e-13
L_PTL_IP2_2|_RX|P2 _PTL_IP2_2|_RX|5 0  5.431e-13
L_PTL_IP2_2|_RX|P3 _PTL_IP2_2|_RX|8 0  5.339e-13
R_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|101  4.225701121488
R_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|104  3.429952209
R_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|107  2.7439617672
L_PTL_IP2_2|_RX|RB1 _PTL_IP2_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_2|_RX|RB2 _PTL_IP2_2|_RX|104 0  1.937922998085e-12
L_PTL_IP2_2|_RX|RB3 _PTL_IP2_2|_RX|107 0  1.550338398468e-12
B_PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP2_2|_JTL|2 _PTL_IP2_2|_JTL|6 _PTL_IP2_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP2_2|_JTL|B1 0 _PTL_IP2_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP2_2|_JTL|1 _PTL_IP2_2|A_PTL_RX _PTL_IP2_2|_JTL|1  2.067833848e-12
L_PTL_IP2_2|_JTL|2 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|4  2.067833848e-12
L_PTL_IP2_2|_JTL|3 _PTL_IP2_2|_JTL|4 _PTL_IP2_2|_JTL|6  2.067833848e-12
L_PTL_IP2_2|_JTL|4 _PTL_IP2_2|_JTL|6 IP2_2_OUT_RX  2.067833848e-12
L_PTL_IP2_2|_JTL|P1 _PTL_IP2_2|_JTL|2 0  2e-13
L_PTL_IP2_2|_JTL|P2 _PTL_IP2_2|_JTL|7 0  2e-13
L_PTL_IP2_2|_JTL|B1 _PTL_IP2_2|_JTL|5 _PTL_IP2_2|_JTL|4  2e-12
R_PTL_IP2_2|_JTL|B1 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|3  2.7439617672
R_PTL_IP2_2|_JTL|B2 _PTL_IP2_2|_JTL|6 _PTL_IP2_2|_JTL|8  2.7439617672
L_PTL_IP2_2|_JTL|RB1 _PTL_IP2_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP2_2|_JTL|RB2 _PTL_IP2_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_2|_TX|B1 0 _PTL_IP3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_2|_TX|B2 0 _PTL_IP3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|3  1.684e-12
L_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|6  3.596e-12
L_PTL_IP3_2|_TX|1 IP3_2_OUT _PTL_IP3_2|_TX|1  2.063e-12
L_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|4  4.123e-12
L_PTL_IP3_2|_TX|3 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|7  2.193e-12
R_PTL_IP3_2|_TX|D _PTL_IP3_2|_TX|7 _PTL_IP3_2|A_PTL  1.36
L_PTL_IP3_2|_TX|P1 _PTL_IP3_2|_TX|2 0  5.254e-13
L_PTL_IP3_2|_TX|P2 _PTL_IP3_2|_TX|5 0  5.141e-13
R_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|101  2.7439617672
R_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|104  2.7439617672
L_PTL_IP3_2|_TX|RB1 _PTL_IP3_2|_TX|101 0  1.550338398468e-12
L_PTL_IP3_2|_TX|RB2 _PTL_IP3_2|_TX|104 0  1.550338398468e-12
B_PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_2|_RX|B1 0 _PTL_IP3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|3  2.777e-12
I_PTL_IP3_2|_RX|B2 0 _PTL_IP3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|6  2.685e-12
I_PTL_IP3_2|_RX|B3 0 _PTL_IP3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|9  2.764e-12
L_PTL_IP3_2|_RX|1 _PTL_IP3_2|A_PTL _PTL_IP3_2|_RX|1  1.346e-12
L_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|4  6.348e-12
L_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7  5.197e-12
L_PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7 _PTL_IP3_2|A_PTL_RX  2.058e-12
L_PTL_IP3_2|_RX|P1 _PTL_IP3_2|_RX|2 0  4.795e-13
L_PTL_IP3_2|_RX|P2 _PTL_IP3_2|_RX|5 0  5.431e-13
L_PTL_IP3_2|_RX|P3 _PTL_IP3_2|_RX|8 0  5.339e-13
R_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|101  4.225701121488
R_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|104  3.429952209
R_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|107  2.7439617672
L_PTL_IP3_2|_RX|RB1 _PTL_IP3_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_2|_RX|RB2 _PTL_IP3_2|_RX|104 0  1.937922998085e-12
L_PTL_IP3_2|_RX|RB3 _PTL_IP3_2|_RX|107 0  1.550338398468e-12
B_PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP3_2|_JTL|2 _PTL_IP3_2|_JTL|6 _PTL_IP3_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP3_2|_JTL|B1 0 _PTL_IP3_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP3_2|_JTL|1 _PTL_IP3_2|A_PTL_RX _PTL_IP3_2|_JTL|1  2.067833848e-12
L_PTL_IP3_2|_JTL|2 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|4  2.067833848e-12
L_PTL_IP3_2|_JTL|3 _PTL_IP3_2|_JTL|4 _PTL_IP3_2|_JTL|6  2.067833848e-12
L_PTL_IP3_2|_JTL|4 _PTL_IP3_2|_JTL|6 IP3_2_OUT_RX  2.067833848e-12
L_PTL_IP3_2|_JTL|P1 _PTL_IP3_2|_JTL|2 0  2e-13
L_PTL_IP3_2|_JTL|P2 _PTL_IP3_2|_JTL|7 0  2e-13
L_PTL_IP3_2|_JTL|B1 _PTL_IP3_2|_JTL|5 _PTL_IP3_2|_JTL|4  2e-12
R_PTL_IP3_2|_JTL|B1 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|3  2.7439617672
R_PTL_IP3_2|_JTL|B2 _PTL_IP3_2|_JTL|6 _PTL_IP3_2|_JTL|8  2.7439617672
L_PTL_IP3_2|_JTL|RB1 _PTL_IP3_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP3_2|_JTL|RB2 _PTL_IP3_2|_JTL|8 0  1.750338398468e-12
L_S0|I_1|B _S0|A1 _S0|I_1|MID  2e-12
I_S0|I_1|B 0 _S0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_3|B _S0|A3 _S0|I_3|MID  2e-12
I_S0|I_3|B 0 _S0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0|I_T|B _S0|T1 _S0|I_T|MID  2e-12
I_S0|I_T|B 0 _S0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_6|B _S0|Q1 _S0|I_6|MID  2e-12
I_S0|I_6|B 0 _S0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0|1|1 _S0|A1 _S0|1|MID_SERIES JJMIT AREA=2.5
L_S0|1|P _S0|1|MID_SERIES 0  2e-13
R_S0|1|B _S0|A1 _S0|1|MID_SHUNT  2.7439617672
L_S0|1|RB _S0|1|MID_SHUNT 0  1.550338398468e-12
B_S0|23|1 _S0|A2 _S0|A3 JJMIT AREA=1.7857142857142858
R_S0|23|B _S0|A2 _S0|23|MID_SHUNT  3.84154647408
L_S0|23|RB _S0|23|MID_SHUNT _S0|A3  2.1704737578552e-12
B_S0|3|1 _S0|A3 _S0|3|MID_SERIES JJMIT AREA=2.5
L_S0|3|P _S0|3|MID_SERIES 0  2e-13
R_S0|3|B _S0|A3 _S0|3|MID_SHUNT  2.7439617672
L_S0|3|RB _S0|3|MID_SHUNT 0  1.550338398468e-12
B_S0|4|1 _S0|A4 _S0|4|MID_SERIES JJMIT AREA=2.5
L_S0|4|P _S0|4|MID_SERIES 0  2e-13
R_S0|4|B _S0|A4 _S0|4|MID_SHUNT  2.7439617672
L_S0|4|RB _S0|4|MID_SHUNT 0  1.550338398468e-12
B_S0|T|1 _S0|T1 _S0|T|MID_SERIES JJMIT AREA=2.5
L_S0|T|P _S0|T|MID_SERIES 0  2e-13
R_S0|T|B _S0|T1 _S0|T|MID_SHUNT  2.7439617672
L_S0|T|RB _S0|T|MID_SHUNT 0  1.550338398468e-12
B_S0|45|1 _S0|T2 _S0|A4 JJMIT AREA=1.7857142857142858
R_S0|45|B _S0|T2 _S0|45|MID_SHUNT  3.84154647408
L_S0|45|RB _S0|45|MID_SHUNT _S0|A4  2.1704737578552e-12
B_S0|6|1 _S0|Q1 _S0|6|MID_SERIES JJMIT AREA=2.5
L_S0|6|P _S0|6|MID_SERIES 0  2e-13
R_S0|6|B _S0|Q1 _S0|6|MID_SHUNT  2.7439617672
L_S0|6|RB _S0|6|MID_SHUNT 0  1.550338398468e-12
L_S1|I_A1|B _S1|A1 _S1|I_A1|MID  2e-12
I_S1|I_A1|B 0 _S1|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_A3|B _S1|A3 _S1|I_A3|MID  2e-12
I_S1|I_A3|B 0 _S1|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B1|B _S1|B1 _S1|I_B1|MID  2e-12
I_S1|I_B1|B 0 _S1|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B3|B _S1|B3 _S1|I_B3|MID  2e-12
I_S1|I_B3|B 0 _S1|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_Q1|B _S1|Q1 _S1|I_Q1|MID  2e-12
I_S1|I_Q1|B 0 _S1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S1|A1|1 _S1|A1 _S1|A1|MID_SERIES JJMIT AREA=2.5
L_S1|A1|P _S1|A1|MID_SERIES 0  5e-13
R_S1|A1|B _S1|A1 _S1|A1|MID_SHUNT  2.7439617672
L_S1|A1|RB _S1|A1|MID_SHUNT 0  2.050338398468e-12
B_S1|A2|1 _S1|A2 _S1|A2|MID_SERIES JJMIT AREA=2.5
L_S1|A2|P _S1|A2|MID_SERIES 0  5e-13
R_S1|A2|B _S1|A2 _S1|A2|MID_SHUNT  2.7439617672
L_S1|A2|RB _S1|A2|MID_SHUNT 0  2.050338398468e-12
B_S1|A3|1 _S1|A2 _S1|A3|MID_SERIES JJMIT AREA=2.5
L_S1|A3|P _S1|A3|MID_SERIES _S1|A3  1.2e-12
R_S1|A3|B _S1|A2 _S1|A3|MID_SHUNT  2.7439617672
L_S1|A3|RB _S1|A3|MID_SHUNT _S1|A3  2.050338398468e-12
B_S1|B1|1 _S1|B1 _S1|B1|MID_SERIES JJMIT AREA=2.5
L_S1|B1|P _S1|B1|MID_SERIES 0  5e-13
R_S1|B1|B _S1|B1 _S1|B1|MID_SHUNT  2.7439617672
L_S1|B1|RB _S1|B1|MID_SHUNT 0  2.050338398468e-12
B_S1|B2|1 _S1|B2 _S1|B2|MID_SERIES JJMIT AREA=2.5
L_S1|B2|P _S1|B2|MID_SERIES 0  5e-13
R_S1|B2|B _S1|B2 _S1|B2|MID_SHUNT  2.7439617672
L_S1|B2|RB _S1|B2|MID_SHUNT 0  2.050338398468e-12
B_S1|B3|1 _S1|B2 _S1|B3|MID_SERIES JJMIT AREA=2.5
L_S1|B3|P _S1|B3|MID_SERIES _S1|B3  1.2e-12
R_S1|B3|B _S1|B2 _S1|B3|MID_SHUNT  2.7439617672
L_S1|B3|RB _S1|B3|MID_SHUNT _S1|B3  2.050338398468e-12
B_S1|T1|1 _S1|T1 _S1|T1|MID_SERIES JJMIT AREA=2.5
L_S1|T1|P _S1|T1|MID_SERIES 0  5e-13
R_S1|T1|B _S1|T1 _S1|T1|MID_SHUNT  2.7439617672
L_S1|T1|RB _S1|T1|MID_SHUNT 0  2.050338398468e-12
B_S1|T2|1 _S1|T2 _S1|ABTQ JJMIT AREA=2.0
R_S1|T2|B _S1|T2 _S1|T2|MID_SHUNT  3.429952209
L_S1|T2|RB _S1|T2|MID_SHUNT _S1|ABTQ  2.437922998085e-12
B_S1|AB|1 _S1|AB _S1|AB|MID_SERIES JJMIT AREA=1.5
L_S1|AB|P _S1|AB|MID_SERIES _S1|ABTQ  1.2e-12
R_S1|AB|B _S1|AB _S1|AB|MID_SHUNT  4.573269612
L_S1|AB|RB _S1|AB|MID_SHUNT _S1|ABTQ  3.08389733078e-12
B_S1|ABTQ|1 _S1|ABTQ _S1|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S1|ABTQ|P _S1|ABTQ|MID_SERIES 0  5e-13
R_S1|ABTQ|B _S1|ABTQ _S1|ABTQ|MID_SHUNT  3.6586156896
L_S1|ABTQ|RB _S1|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S1|Q1|1 _S1|Q1 _S1|Q1|MID_SERIES JJMIT AREA=2.5
L_S1|Q1|P _S1|Q1|MID_SERIES 0  5e-13
R_S1|Q1|B _S1|Q1 _S1|Q1|MID_SHUNT  2.7439617672
L_S1|Q1|RB _S1|Q1|MID_SHUNT 0  2.050338398468e-12
L_S2|I_A1|B _S2|A1 _S2|I_A1|MID  2e-12
I_S2|I_A1|B 0 _S2|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_A3|B _S2|A3 _S2|I_A3|MID  2e-12
I_S2|I_A3|B 0 _S2|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B1|B _S2|B1 _S2|I_B1|MID  2e-12
I_S2|I_B1|B 0 _S2|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B3|B _S2|B3 _S2|I_B3|MID  2e-12
I_S2|I_B3|B 0 _S2|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_Q1|B _S2|Q1 _S2|I_Q1|MID  2e-12
I_S2|I_Q1|B 0 _S2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S2|A1|1 _S2|A1 _S2|A1|MID_SERIES JJMIT AREA=2.5
L_S2|A1|P _S2|A1|MID_SERIES 0  5e-13
R_S2|A1|B _S2|A1 _S2|A1|MID_SHUNT  2.7439617672
L_S2|A1|RB _S2|A1|MID_SHUNT 0  2.050338398468e-12
B_S2|A2|1 _S2|A2 _S2|A2|MID_SERIES JJMIT AREA=2.5
L_S2|A2|P _S2|A2|MID_SERIES 0  5e-13
R_S2|A2|B _S2|A2 _S2|A2|MID_SHUNT  2.7439617672
L_S2|A2|RB _S2|A2|MID_SHUNT 0  2.050338398468e-12
B_S2|A3|1 _S2|A2 _S2|A3|MID_SERIES JJMIT AREA=2.5
L_S2|A3|P _S2|A3|MID_SERIES _S2|A3  1.2e-12
R_S2|A3|B _S2|A2 _S2|A3|MID_SHUNT  2.7439617672
L_S2|A3|RB _S2|A3|MID_SHUNT _S2|A3  2.050338398468e-12
B_S2|B1|1 _S2|B1 _S2|B1|MID_SERIES JJMIT AREA=2.5
L_S2|B1|P _S2|B1|MID_SERIES 0  5e-13
R_S2|B1|B _S2|B1 _S2|B1|MID_SHUNT  2.7439617672
L_S2|B1|RB _S2|B1|MID_SHUNT 0  2.050338398468e-12
B_S2|B2|1 _S2|B2 _S2|B2|MID_SERIES JJMIT AREA=2.5
L_S2|B2|P _S2|B2|MID_SERIES 0  5e-13
R_S2|B2|B _S2|B2 _S2|B2|MID_SHUNT  2.7439617672
L_S2|B2|RB _S2|B2|MID_SHUNT 0  2.050338398468e-12
B_S2|B3|1 _S2|B2 _S2|B3|MID_SERIES JJMIT AREA=2.5
L_S2|B3|P _S2|B3|MID_SERIES _S2|B3  1.2e-12
R_S2|B3|B _S2|B2 _S2|B3|MID_SHUNT  2.7439617672
L_S2|B3|RB _S2|B3|MID_SHUNT _S2|B3  2.050338398468e-12
B_S2|T1|1 _S2|T1 _S2|T1|MID_SERIES JJMIT AREA=2.5
L_S2|T1|P _S2|T1|MID_SERIES 0  5e-13
R_S2|T1|B _S2|T1 _S2|T1|MID_SHUNT  2.7439617672
L_S2|T1|RB _S2|T1|MID_SHUNT 0  2.050338398468e-12
B_S2|T2|1 _S2|T2 _S2|ABTQ JJMIT AREA=2.0
R_S2|T2|B _S2|T2 _S2|T2|MID_SHUNT  3.429952209
L_S2|T2|RB _S2|T2|MID_SHUNT _S2|ABTQ  2.437922998085e-12
B_S2|AB|1 _S2|AB _S2|AB|MID_SERIES JJMIT AREA=1.5
L_S2|AB|P _S2|AB|MID_SERIES _S2|ABTQ  1.2e-12
R_S2|AB|B _S2|AB _S2|AB|MID_SHUNT  4.573269612
L_S2|AB|RB _S2|AB|MID_SHUNT _S2|ABTQ  3.08389733078e-12
B_S2|ABTQ|1 _S2|ABTQ _S2|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S2|ABTQ|P _S2|ABTQ|MID_SERIES 0  5e-13
R_S2|ABTQ|B _S2|ABTQ _S2|ABTQ|MID_SHUNT  3.6586156896
L_S2|ABTQ|RB _S2|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S2|Q1|1 _S2|Q1 _S2|Q1|MID_SERIES JJMIT AREA=2.5
L_S2|Q1|P _S2|Q1|MID_SERIES 0  5e-13
R_S2|Q1|B _S2|Q1 _S2|Q1|MID_SHUNT  2.7439617672
L_S2|Q1|RB _S2|Q1|MID_SHUNT 0  2.050338398468e-12
L_S3|I_A1|B _S3|A1 _S3|I_A1|MID  2e-12
I_S3|I_A1|B 0 _S3|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_A3|B _S3|A3 _S3|I_A3|MID  2e-12
I_S3|I_A3|B 0 _S3|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B1|B _S3|B1 _S3|I_B1|MID  2e-12
I_S3|I_B1|B 0 _S3|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B3|B _S3|B3 _S3|I_B3|MID  2e-12
I_S3|I_B3|B 0 _S3|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_Q1|B _S3|Q1 _S3|I_Q1|MID  2e-12
I_S3|I_Q1|B 0 _S3|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S3|A1|1 _S3|A1 _S3|A1|MID_SERIES JJMIT AREA=2.5
L_S3|A1|P _S3|A1|MID_SERIES 0  5e-13
R_S3|A1|B _S3|A1 _S3|A1|MID_SHUNT  2.7439617672
L_S3|A1|RB _S3|A1|MID_SHUNT 0  2.050338398468e-12
B_S3|A2|1 _S3|A2 _S3|A2|MID_SERIES JJMIT AREA=2.5
L_S3|A2|P _S3|A2|MID_SERIES 0  5e-13
R_S3|A2|B _S3|A2 _S3|A2|MID_SHUNT  2.7439617672
L_S3|A2|RB _S3|A2|MID_SHUNT 0  2.050338398468e-12
B_S3|A3|1 _S3|A2 _S3|A3|MID_SERIES JJMIT AREA=2.5
L_S3|A3|P _S3|A3|MID_SERIES _S3|A3  1.2e-12
R_S3|A3|B _S3|A2 _S3|A3|MID_SHUNT  2.7439617672
L_S3|A3|RB _S3|A3|MID_SHUNT _S3|A3  2.050338398468e-12
B_S3|B1|1 _S3|B1 _S3|B1|MID_SERIES JJMIT AREA=2.5
L_S3|B1|P _S3|B1|MID_SERIES 0  5e-13
R_S3|B1|B _S3|B1 _S3|B1|MID_SHUNT  2.7439617672
L_S3|B1|RB _S3|B1|MID_SHUNT 0  2.050338398468e-12
B_S3|B2|1 _S3|B2 _S3|B2|MID_SERIES JJMIT AREA=2.5
L_S3|B2|P _S3|B2|MID_SERIES 0  5e-13
R_S3|B2|B _S3|B2 _S3|B2|MID_SHUNT  2.7439617672
L_S3|B2|RB _S3|B2|MID_SHUNT 0  2.050338398468e-12
B_S3|B3|1 _S3|B2 _S3|B3|MID_SERIES JJMIT AREA=2.5
L_S3|B3|P _S3|B3|MID_SERIES _S3|B3  1.2e-12
R_S3|B3|B _S3|B2 _S3|B3|MID_SHUNT  2.7439617672
L_S3|B3|RB _S3|B3|MID_SHUNT _S3|B3  2.050338398468e-12
B_S3|T1|1 _S3|T1 _S3|T1|MID_SERIES JJMIT AREA=2.5
L_S3|T1|P _S3|T1|MID_SERIES 0  5e-13
R_S3|T1|B _S3|T1 _S3|T1|MID_SHUNT  2.7439617672
L_S3|T1|RB _S3|T1|MID_SHUNT 0  2.050338398468e-12
B_S3|T2|1 _S3|T2 _S3|ABTQ JJMIT AREA=2.0
R_S3|T2|B _S3|T2 _S3|T2|MID_SHUNT  3.429952209
L_S3|T2|RB _S3|T2|MID_SHUNT _S3|ABTQ  2.437922998085e-12
B_S3|AB|1 _S3|AB _S3|AB|MID_SERIES JJMIT AREA=1.5
L_S3|AB|P _S3|AB|MID_SERIES _S3|ABTQ  1.2e-12
R_S3|AB|B _S3|AB _S3|AB|MID_SHUNT  4.573269612
L_S3|AB|RB _S3|AB|MID_SHUNT _S3|ABTQ  3.08389733078e-12
B_S3|ABTQ|1 _S3|ABTQ _S3|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S3|ABTQ|P _S3|ABTQ|MID_SERIES 0  5e-13
R_S3|ABTQ|B _S3|ABTQ _S3|ABTQ|MID_SHUNT  3.6586156896
L_S3|ABTQ|RB _S3|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S3|Q1|1 _S3|Q1 _S3|Q1|MID_SERIES JJMIT AREA=2.5
L_S3|Q1|P _S3|Q1|MID_SERIES 0  5e-13
R_S3|Q1|B _S3|Q1 _S3|Q1|MID_SHUNT  2.7439617672
L_S3|Q1|RB _S3|Q1|MID_SHUNT 0  2.050338398468e-12
L_S4|I_1|B _S4|A1 _S4|I_1|MID  2e-12
I_S4|I_1|B 0 _S4|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_3|B _S4|A3 _S4|I_3|MID  2e-12
I_S4|I_3|B 0 _S4|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S4|I_T|B _S4|T1 _S4|I_T|MID  2e-12
I_S4|I_T|B 0 _S4|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_6|B _S4|Q1 _S4|I_6|MID  2e-12
I_S4|I_6|B 0 _S4|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S4|1|1 _S4|A1 _S4|1|MID_SERIES JJMIT AREA=2.5
L_S4|1|P _S4|1|MID_SERIES 0  2e-13
R_S4|1|B _S4|A1 _S4|1|MID_SHUNT  2.7439617672
L_S4|1|RB _S4|1|MID_SHUNT 0  1.550338398468e-12
B_S4|23|1 _S4|A2 _S4|A3 JJMIT AREA=1.7857142857142858
R_S4|23|B _S4|A2 _S4|23|MID_SHUNT  3.84154647408
L_S4|23|RB _S4|23|MID_SHUNT _S4|A3  2.1704737578552e-12
B_S4|3|1 _S4|A3 _S4|3|MID_SERIES JJMIT AREA=2.5
L_S4|3|P _S4|3|MID_SERIES 0  2e-13
R_S4|3|B _S4|A3 _S4|3|MID_SHUNT  2.7439617672
L_S4|3|RB _S4|3|MID_SHUNT 0  1.550338398468e-12
B_S4|4|1 _S4|A4 _S4|4|MID_SERIES JJMIT AREA=2.5
L_S4|4|P _S4|4|MID_SERIES 0  2e-13
R_S4|4|B _S4|A4 _S4|4|MID_SHUNT  2.7439617672
L_S4|4|RB _S4|4|MID_SHUNT 0  1.550338398468e-12
B_S4|T|1 _S4|T1 _S4|T|MID_SERIES JJMIT AREA=2.5
L_S4|T|P _S4|T|MID_SERIES 0  2e-13
R_S4|T|B _S4|T1 _S4|T|MID_SHUNT  2.7439617672
L_S4|T|RB _S4|T|MID_SHUNT 0  1.550338398468e-12
B_S4|45|1 _S4|T2 _S4|A4 JJMIT AREA=1.7857142857142858
R_S4|45|B _S4|T2 _S4|45|MID_SHUNT  3.84154647408
L_S4|45|RB _S4|45|MID_SHUNT _S4|A4  2.1704737578552e-12
B_S4|6|1 _S4|Q1 _S4|6|MID_SERIES JJMIT AREA=2.5
L_S4|6|P _S4|6|MID_SERIES 0  2e-13
R_S4|6|B _S4|Q1 _S4|6|MID_SHUNT  2.7439617672
L_S4|6|RB _S4|6|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_A|I_D1|B I0|_SPL_A|D1 I0|_SPL_A|I_D1|MID  2e-12
II0|_SPL_A|I_D1|B 0 I0|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_D2|B I0|_SPL_A|D2 I0|_SPL_A|I_D2|MID  2e-12
II0|_SPL_A|I_D2|B 0 I0|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_A|I_Q1|B I0|_SPL_A|QA1 I0|_SPL_A|I_Q1|MID  2e-12
II0|_SPL_A|I_Q1|B 0 I0|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_Q2|B I0|_SPL_A|QB1 I0|_SPL_A|I_Q2|MID  2e-12
II0|_SPL_A|I_Q2|B 0 I0|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_A|1|1 I0|_SPL_A|D1 I0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|1|P I0|_SPL_A|1|MID_SERIES 0  2e-13
RI0|_SPL_A|1|B I0|_SPL_A|D1 I0|_SPL_A|1|MID_SHUNT  2.7439617672
LI0|_SPL_A|1|RB I0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|2|1 I0|_SPL_A|D2 I0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|2|P I0|_SPL_A|2|MID_SERIES 0  2e-13
RI0|_SPL_A|2|B I0|_SPL_A|D2 I0|_SPL_A|2|MID_SHUNT  2.7439617672
LI0|_SPL_A|2|RB I0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|A|1 I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|A|P I0|_SPL_A|A|MID_SERIES 0  2e-13
RI0|_SPL_A|A|B I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SHUNT  2.7439617672
LI0|_SPL_A|A|RB I0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|B|1 I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|B|P I0|_SPL_A|B|MID_SERIES 0  2e-13
RI0|_SPL_A|B|B I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SHUNT  2.7439617672
LI0|_SPL_A|B|RB I0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_B|I_D1|B I0|_SPL_B|D1 I0|_SPL_B|I_D1|MID  2e-12
II0|_SPL_B|I_D1|B 0 I0|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_D2|B I0|_SPL_B|D2 I0|_SPL_B|I_D2|MID  2e-12
II0|_SPL_B|I_D2|B 0 I0|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_B|I_Q1|B I0|_SPL_B|QA1 I0|_SPL_B|I_Q1|MID  2e-12
II0|_SPL_B|I_Q1|B 0 I0|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_Q2|B I0|_SPL_B|QB1 I0|_SPL_B|I_Q2|MID  2e-12
II0|_SPL_B|I_Q2|B 0 I0|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_B|1|1 I0|_SPL_B|D1 I0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|1|P I0|_SPL_B|1|MID_SERIES 0  2e-13
RI0|_SPL_B|1|B I0|_SPL_B|D1 I0|_SPL_B|1|MID_SHUNT  2.7439617672
LI0|_SPL_B|1|RB I0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|2|1 I0|_SPL_B|D2 I0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|2|P I0|_SPL_B|2|MID_SERIES 0  2e-13
RI0|_SPL_B|2|B I0|_SPL_B|D2 I0|_SPL_B|2|MID_SHUNT  2.7439617672
LI0|_SPL_B|2|RB I0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|A|1 I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|A|P I0|_SPL_B|A|MID_SERIES 0  2e-13
RI0|_SPL_B|A|B I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SHUNT  2.7439617672
LI0|_SPL_B|A|RB I0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|B|1 I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|B|P I0|_SPL_B|B|MID_SERIES 0  2e-13
RI0|_SPL_B|B|B I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SHUNT  2.7439617672
LI0|_SPL_B|B|RB I0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_A|I_1|B I0|_DFF_A|A1 I0|_DFF_A|I_1|MID  2e-12
II0|_DFF_A|I_1|B 0 I0|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_3|B I0|_DFF_A|A3 I0|_DFF_A|I_3|MID  2e-12
II0|_DFF_A|I_3|B 0 I0|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_A|I_T|B I0|_DFF_A|T1 I0|_DFF_A|I_T|MID  2e-12
II0|_DFF_A|I_T|B 0 I0|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_6|B I0|_DFF_A|Q1 I0|_DFF_A|I_6|MID  2e-12
II0|_DFF_A|I_6|B 0 I0|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_A|1|1 I0|_DFF_A|A1 I0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|1|P I0|_DFF_A|1|MID_SERIES 0  2e-13
RI0|_DFF_A|1|B I0|_DFF_A|A1 I0|_DFF_A|1|MID_SHUNT  2.7439617672
LI0|_DFF_A|1|RB I0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|23|1 I0|_DFF_A|A2 I0|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|23|B I0|_DFF_A|A2 I0|_DFF_A|23|MID_SHUNT  3.84154647408
LI0|_DFF_A|23|RB I0|_DFF_A|23|MID_SHUNT I0|_DFF_A|A3  2.1704737578552e-12
BI0|_DFF_A|3|1 I0|_DFF_A|A3 I0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|3|P I0|_DFF_A|3|MID_SERIES 0  2e-13
RI0|_DFF_A|3|B I0|_DFF_A|A3 I0|_DFF_A|3|MID_SHUNT  2.7439617672
LI0|_DFF_A|3|RB I0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|4|1 I0|_DFF_A|A4 I0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|4|P I0|_DFF_A|4|MID_SERIES 0  2e-13
RI0|_DFF_A|4|B I0|_DFF_A|A4 I0|_DFF_A|4|MID_SHUNT  2.7439617672
LI0|_DFF_A|4|RB I0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|T|1 I0|_DFF_A|T1 I0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|T|P I0|_DFF_A|T|MID_SERIES 0  2e-13
RI0|_DFF_A|T|B I0|_DFF_A|T1 I0|_DFF_A|T|MID_SHUNT  2.7439617672
LI0|_DFF_A|T|RB I0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|45|1 I0|_DFF_A|T2 I0|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|45|B I0|_DFF_A|T2 I0|_DFF_A|45|MID_SHUNT  3.84154647408
LI0|_DFF_A|45|RB I0|_DFF_A|45|MID_SHUNT I0|_DFF_A|A4  2.1704737578552e-12
BI0|_DFF_A|6|1 I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|6|P I0|_DFF_A|6|MID_SERIES 0  2e-13
RI0|_DFF_A|6|B I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SHUNT  2.7439617672
LI0|_DFF_A|6|RB I0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_B|I_1|B I0|_DFF_B|A1 I0|_DFF_B|I_1|MID  2e-12
II0|_DFF_B|I_1|B 0 I0|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_3|B I0|_DFF_B|A3 I0|_DFF_B|I_3|MID  2e-12
II0|_DFF_B|I_3|B 0 I0|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_B|I_T|B I0|_DFF_B|T1 I0|_DFF_B|I_T|MID  2e-12
II0|_DFF_B|I_T|B 0 I0|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_6|B I0|_DFF_B|Q1 I0|_DFF_B|I_6|MID  2e-12
II0|_DFF_B|I_6|B 0 I0|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_B|1|1 I0|_DFF_B|A1 I0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|1|P I0|_DFF_B|1|MID_SERIES 0  2e-13
RI0|_DFF_B|1|B I0|_DFF_B|A1 I0|_DFF_B|1|MID_SHUNT  2.7439617672
LI0|_DFF_B|1|RB I0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|23|1 I0|_DFF_B|A2 I0|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|23|B I0|_DFF_B|A2 I0|_DFF_B|23|MID_SHUNT  3.84154647408
LI0|_DFF_B|23|RB I0|_DFF_B|23|MID_SHUNT I0|_DFF_B|A3  2.1704737578552e-12
BI0|_DFF_B|3|1 I0|_DFF_B|A3 I0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|3|P I0|_DFF_B|3|MID_SERIES 0  2e-13
RI0|_DFF_B|3|B I0|_DFF_B|A3 I0|_DFF_B|3|MID_SHUNT  2.7439617672
LI0|_DFF_B|3|RB I0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|4|1 I0|_DFF_B|A4 I0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|4|P I0|_DFF_B|4|MID_SERIES 0  2e-13
RI0|_DFF_B|4|B I0|_DFF_B|A4 I0|_DFF_B|4|MID_SHUNT  2.7439617672
LI0|_DFF_B|4|RB I0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|T|1 I0|_DFF_B|T1 I0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|T|P I0|_DFF_B|T|MID_SERIES 0  2e-13
RI0|_DFF_B|T|B I0|_DFF_B|T1 I0|_DFF_B|T|MID_SHUNT  2.7439617672
LI0|_DFF_B|T|RB I0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|45|1 I0|_DFF_B|T2 I0|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|45|B I0|_DFF_B|T2 I0|_DFF_B|45|MID_SHUNT  3.84154647408
LI0|_DFF_B|45|RB I0|_DFF_B|45|MID_SHUNT I0|_DFF_B|A4  2.1704737578552e-12
BI0|_DFF_B|6|1 I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|6|P I0|_DFF_B|6|MID_SERIES 0  2e-13
RI0|_DFF_B|6|B I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SHUNT  2.7439617672
LI0|_DFF_B|6|RB I0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI0|_XOR|I_A1|B I0|_XOR|A1 I0|_XOR|I_A1|MID  2e-12
II0|_XOR|I_A1|B 0 I0|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_A3|B I0|_XOR|A3 I0|_XOR|I_A3|MID  2e-12
II0|_XOR|I_A3|B 0 I0|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B1|B I0|_XOR|B1 I0|_XOR|I_B1|MID  2e-12
II0|_XOR|I_B1|B 0 I0|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B3|B I0|_XOR|B3 I0|_XOR|I_B3|MID  2e-12
II0|_XOR|I_B3|B 0 I0|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_Q1|B I0|_XOR|Q1 I0|_XOR|I_Q1|MID  2e-12
II0|_XOR|I_Q1|B 0 I0|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_XOR|A1|1 I0|_XOR|A1 I0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A1|P I0|_XOR|A1|MID_SERIES 0  5e-13
RI0|_XOR|A1|B I0|_XOR|A1 I0|_XOR|A1|MID_SHUNT  2.7439617672
LI0|_XOR|A1|RB I0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A2|1 I0|_XOR|A2 I0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A2|P I0|_XOR|A2|MID_SERIES 0  5e-13
RI0|_XOR|A2|B I0|_XOR|A2 I0|_XOR|A2|MID_SHUNT  2.7439617672
LI0|_XOR|A2|RB I0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A3|1 I0|_XOR|A2 I0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A3|P I0|_XOR|A3|MID_SERIES I0|_XOR|A3  1.2e-12
RI0|_XOR|A3|B I0|_XOR|A2 I0|_XOR|A3|MID_SHUNT  2.7439617672
LI0|_XOR|A3|RB I0|_XOR|A3|MID_SHUNT I0|_XOR|A3  2.050338398468e-12
BI0|_XOR|B1|1 I0|_XOR|B1 I0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B1|P I0|_XOR|B1|MID_SERIES 0  5e-13
RI0|_XOR|B1|B I0|_XOR|B1 I0|_XOR|B1|MID_SHUNT  2.7439617672
LI0|_XOR|B1|RB I0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B2|1 I0|_XOR|B2 I0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B2|P I0|_XOR|B2|MID_SERIES 0  5e-13
RI0|_XOR|B2|B I0|_XOR|B2 I0|_XOR|B2|MID_SHUNT  2.7439617672
LI0|_XOR|B2|RB I0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B3|1 I0|_XOR|B2 I0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B3|P I0|_XOR|B3|MID_SERIES I0|_XOR|B3  1.2e-12
RI0|_XOR|B3|B I0|_XOR|B2 I0|_XOR|B3|MID_SHUNT  2.7439617672
LI0|_XOR|B3|RB I0|_XOR|B3|MID_SHUNT I0|_XOR|B3  2.050338398468e-12
BI0|_XOR|T1|1 I0|_XOR|T1 I0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|T1|P I0|_XOR|T1|MID_SERIES 0  5e-13
RI0|_XOR|T1|B I0|_XOR|T1 I0|_XOR|T1|MID_SHUNT  2.7439617672
LI0|_XOR|T1|RB I0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|T2|1 I0|_XOR|T2 I0|_XOR|ABTQ JJMIT AREA=2.0
RI0|_XOR|T2|B I0|_XOR|T2 I0|_XOR|T2|MID_SHUNT  3.429952209
LI0|_XOR|T2|RB I0|_XOR|T2|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|AB|1 I0|_XOR|AB I0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI0|_XOR|AB|P I0|_XOR|AB|MID_SERIES I0|_XOR|ABTQ  1.2e-12
RI0|_XOR|AB|B I0|_XOR|AB I0|_XOR|AB|MID_SHUNT  3.429952209
LI0|_XOR|AB|RB I0|_XOR|AB|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|ABTQ|1 I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|ABTQ|P I0|_XOR|ABTQ|MID_SERIES 0  5e-13
RI0|_XOR|ABTQ|B I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI0|_XOR|ABTQ|RB I0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|Q1|1 I0|_XOR|Q1 I0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|Q1|P I0|_XOR|Q1|MID_SERIES 0  5e-13
RI0|_XOR|Q1|B I0|_XOR|Q1 I0|_XOR|Q1|MID_SHUNT  2.7439617672
LI0|_XOR|Q1|RB I0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI0|_AND|I_A1|B I0|_AND|A1 I0|_AND|I_A1|MID  2e-12
II0|_AND|I_A1|B 0 I0|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_B1|B I0|_AND|B1 I0|_AND|I_B1|MID  2e-12
II0|_AND|I_B1|B 0 I0|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q3|B I0|_AND|Q3 I0|_AND|I_Q3|MID  2e-12
II0|_AND|I_Q3|B 0 I0|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0|_AND|I_Q2|B I0|_AND|Q2 I0|_AND|I_Q2|MID  2e-12
II0|_AND|I_Q2|B 0 I0|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q1|B I0|_AND|Q1 I0|_AND|I_Q1|MID  2e-12
II0|_AND|I_Q1|B 0 I0|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_AND|A1|1 I0|_AND|A1 I0|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A1|P I0|_AND|A1|MID_SERIES 0  2e-13
RI0|_AND|A1|B I0|_AND|A1 I0|_AND|A1|MID_SHUNT  2.7439617672
LI0|_AND|A1|RB I0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A2|1 I0|_AND|A2 I0|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A2|P I0|_AND|A2|MID_SERIES 0  2e-13
RI0|_AND|A2|B I0|_AND|A2 I0|_AND|A2|MID_SHUNT  2.7439617672
LI0|_AND|A2|RB I0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A12|1 I0|_AND|A2 I0|_AND|A3 JJMIT AREA=1.7857142857142858
RI0|_AND|A12|B I0|_AND|A2 I0|_AND|A12|MID_SHUNT  3.84154647408
LI0|_AND|A12|RB I0|_AND|A12|MID_SHUNT I0|_AND|A3  2.1704737578552e-12
BI0|_AND|B1|1 I0|_AND|B1 I0|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B1|P I0|_AND|B1|MID_SERIES 0  2e-13
RI0|_AND|B1|B I0|_AND|B1 I0|_AND|B1|MID_SHUNT  2.7439617672
LI0|_AND|B1|RB I0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B2|1 I0|_AND|B2 I0|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B2|P I0|_AND|B2|MID_SERIES 0  2e-13
RI0|_AND|B2|B I0|_AND|B2 I0|_AND|B2|MID_SHUNT  2.7439617672
LI0|_AND|B2|RB I0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B12|1 I0|_AND|B2 I0|_AND|B3 JJMIT AREA=1.7857142857142858
RI0|_AND|B12|B I0|_AND|B2 I0|_AND|B12|MID_SHUNT  3.84154647408
LI0|_AND|B12|RB I0|_AND|B12|MID_SHUNT I0|_AND|B3  2.1704737578552e-12
BI0|_AND|Q2|1 I0|_AND|Q2 I0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q2|P I0|_AND|Q2|MID_SERIES 0  2e-13
RI0|_AND|Q2|B I0|_AND|Q2 I0|_AND|Q2|MID_SHUNT  2.7439617672
LI0|_AND|Q2|RB I0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|Q1|1 I0|_AND|Q1 I0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q1|P I0|_AND|Q1|MID_SERIES 0  2e-13
RI0|_AND|Q1|B I0|_AND|Q1 I0|_AND|Q1|MID_SHUNT  2.7439617672
LI0|_AND|Q1|RB I0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_A|I_D1|B I1|_SPL_A|D1 I1|_SPL_A|I_D1|MID  2e-12
II1|_SPL_A|I_D1|B 0 I1|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_D2|B I1|_SPL_A|D2 I1|_SPL_A|I_D2|MID  2e-12
II1|_SPL_A|I_D2|B 0 I1|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_A|I_Q1|B I1|_SPL_A|QA1 I1|_SPL_A|I_Q1|MID  2e-12
II1|_SPL_A|I_Q1|B 0 I1|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_Q2|B I1|_SPL_A|QB1 I1|_SPL_A|I_Q2|MID  2e-12
II1|_SPL_A|I_Q2|B 0 I1|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_A|1|1 I1|_SPL_A|D1 I1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|1|P I1|_SPL_A|1|MID_SERIES 0  2e-13
RI1|_SPL_A|1|B I1|_SPL_A|D1 I1|_SPL_A|1|MID_SHUNT  2.7439617672
LI1|_SPL_A|1|RB I1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|2|1 I1|_SPL_A|D2 I1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|2|P I1|_SPL_A|2|MID_SERIES 0  2e-13
RI1|_SPL_A|2|B I1|_SPL_A|D2 I1|_SPL_A|2|MID_SHUNT  2.7439617672
LI1|_SPL_A|2|RB I1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|A|1 I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|A|P I1|_SPL_A|A|MID_SERIES 0  2e-13
RI1|_SPL_A|A|B I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SHUNT  2.7439617672
LI1|_SPL_A|A|RB I1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|B|1 I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|B|P I1|_SPL_A|B|MID_SERIES 0  2e-13
RI1|_SPL_A|B|B I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SHUNT  2.7439617672
LI1|_SPL_A|B|RB I1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_B|I_D1|B I1|_SPL_B|D1 I1|_SPL_B|I_D1|MID  2e-12
II1|_SPL_B|I_D1|B 0 I1|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_D2|B I1|_SPL_B|D2 I1|_SPL_B|I_D2|MID  2e-12
II1|_SPL_B|I_D2|B 0 I1|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_B|I_Q1|B I1|_SPL_B|QA1 I1|_SPL_B|I_Q1|MID  2e-12
II1|_SPL_B|I_Q1|B 0 I1|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_Q2|B I1|_SPL_B|QB1 I1|_SPL_B|I_Q2|MID  2e-12
II1|_SPL_B|I_Q2|B 0 I1|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_B|1|1 I1|_SPL_B|D1 I1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|1|P I1|_SPL_B|1|MID_SERIES 0  2e-13
RI1|_SPL_B|1|B I1|_SPL_B|D1 I1|_SPL_B|1|MID_SHUNT  2.7439617672
LI1|_SPL_B|1|RB I1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|2|1 I1|_SPL_B|D2 I1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|2|P I1|_SPL_B|2|MID_SERIES 0  2e-13
RI1|_SPL_B|2|B I1|_SPL_B|D2 I1|_SPL_B|2|MID_SHUNT  2.7439617672
LI1|_SPL_B|2|RB I1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|A|1 I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|A|P I1|_SPL_B|A|MID_SERIES 0  2e-13
RI1|_SPL_B|A|B I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SHUNT  2.7439617672
LI1|_SPL_B|A|RB I1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|B|1 I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|B|P I1|_SPL_B|B|MID_SERIES 0  2e-13
RI1|_SPL_B|B|B I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SHUNT  2.7439617672
LI1|_SPL_B|B|RB I1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_A|I_1|B I1|_DFF_A|A1 I1|_DFF_A|I_1|MID  2e-12
II1|_DFF_A|I_1|B 0 I1|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_3|B I1|_DFF_A|A3 I1|_DFF_A|I_3|MID  2e-12
II1|_DFF_A|I_3|B 0 I1|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_A|I_T|B I1|_DFF_A|T1 I1|_DFF_A|I_T|MID  2e-12
II1|_DFF_A|I_T|B 0 I1|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_6|B I1|_DFF_A|Q1 I1|_DFF_A|I_6|MID  2e-12
II1|_DFF_A|I_6|B 0 I1|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_A|1|1 I1|_DFF_A|A1 I1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|1|P I1|_DFF_A|1|MID_SERIES 0  2e-13
RI1|_DFF_A|1|B I1|_DFF_A|A1 I1|_DFF_A|1|MID_SHUNT  2.7439617672
LI1|_DFF_A|1|RB I1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|23|1 I1|_DFF_A|A2 I1|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|23|B I1|_DFF_A|A2 I1|_DFF_A|23|MID_SHUNT  3.84154647408
LI1|_DFF_A|23|RB I1|_DFF_A|23|MID_SHUNT I1|_DFF_A|A3  2.1704737578552e-12
BI1|_DFF_A|3|1 I1|_DFF_A|A3 I1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|3|P I1|_DFF_A|3|MID_SERIES 0  2e-13
RI1|_DFF_A|3|B I1|_DFF_A|A3 I1|_DFF_A|3|MID_SHUNT  2.7439617672
LI1|_DFF_A|3|RB I1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|4|1 I1|_DFF_A|A4 I1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|4|P I1|_DFF_A|4|MID_SERIES 0  2e-13
RI1|_DFF_A|4|B I1|_DFF_A|A4 I1|_DFF_A|4|MID_SHUNT  2.7439617672
LI1|_DFF_A|4|RB I1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|T|1 I1|_DFF_A|T1 I1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|T|P I1|_DFF_A|T|MID_SERIES 0  2e-13
RI1|_DFF_A|T|B I1|_DFF_A|T1 I1|_DFF_A|T|MID_SHUNT  2.7439617672
LI1|_DFF_A|T|RB I1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|45|1 I1|_DFF_A|T2 I1|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|45|B I1|_DFF_A|T2 I1|_DFF_A|45|MID_SHUNT  3.84154647408
LI1|_DFF_A|45|RB I1|_DFF_A|45|MID_SHUNT I1|_DFF_A|A4  2.1704737578552e-12
BI1|_DFF_A|6|1 I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|6|P I1|_DFF_A|6|MID_SERIES 0  2e-13
RI1|_DFF_A|6|B I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SHUNT  2.7439617672
LI1|_DFF_A|6|RB I1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_B|I_1|B I1|_DFF_B|A1 I1|_DFF_B|I_1|MID  2e-12
II1|_DFF_B|I_1|B 0 I1|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_3|B I1|_DFF_B|A3 I1|_DFF_B|I_3|MID  2e-12
II1|_DFF_B|I_3|B 0 I1|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_B|I_T|B I1|_DFF_B|T1 I1|_DFF_B|I_T|MID  2e-12
II1|_DFF_B|I_T|B 0 I1|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_6|B I1|_DFF_B|Q1 I1|_DFF_B|I_6|MID  2e-12
II1|_DFF_B|I_6|B 0 I1|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_B|1|1 I1|_DFF_B|A1 I1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|1|P I1|_DFF_B|1|MID_SERIES 0  2e-13
RI1|_DFF_B|1|B I1|_DFF_B|A1 I1|_DFF_B|1|MID_SHUNT  2.7439617672
LI1|_DFF_B|1|RB I1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|23|1 I1|_DFF_B|A2 I1|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|23|B I1|_DFF_B|A2 I1|_DFF_B|23|MID_SHUNT  3.84154647408
LI1|_DFF_B|23|RB I1|_DFF_B|23|MID_SHUNT I1|_DFF_B|A3  2.1704737578552e-12
BI1|_DFF_B|3|1 I1|_DFF_B|A3 I1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|3|P I1|_DFF_B|3|MID_SERIES 0  2e-13
RI1|_DFF_B|3|B I1|_DFF_B|A3 I1|_DFF_B|3|MID_SHUNT  2.7439617672
LI1|_DFF_B|3|RB I1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|4|1 I1|_DFF_B|A4 I1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|4|P I1|_DFF_B|4|MID_SERIES 0  2e-13
RI1|_DFF_B|4|B I1|_DFF_B|A4 I1|_DFF_B|4|MID_SHUNT  2.7439617672
LI1|_DFF_B|4|RB I1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|T|1 I1|_DFF_B|T1 I1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|T|P I1|_DFF_B|T|MID_SERIES 0  2e-13
RI1|_DFF_B|T|B I1|_DFF_B|T1 I1|_DFF_B|T|MID_SHUNT  2.7439617672
LI1|_DFF_B|T|RB I1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|45|1 I1|_DFF_B|T2 I1|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|45|B I1|_DFF_B|T2 I1|_DFF_B|45|MID_SHUNT  3.84154647408
LI1|_DFF_B|45|RB I1|_DFF_B|45|MID_SHUNT I1|_DFF_B|A4  2.1704737578552e-12
BI1|_DFF_B|6|1 I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|6|P I1|_DFF_B|6|MID_SERIES 0  2e-13
RI1|_DFF_B|6|B I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SHUNT  2.7439617672
LI1|_DFF_B|6|RB I1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI1|_XOR|I_A1|B I1|_XOR|A1 I1|_XOR|I_A1|MID  2e-12
II1|_XOR|I_A1|B 0 I1|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_A3|B I1|_XOR|A3 I1|_XOR|I_A3|MID  2e-12
II1|_XOR|I_A3|B 0 I1|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B1|B I1|_XOR|B1 I1|_XOR|I_B1|MID  2e-12
II1|_XOR|I_B1|B 0 I1|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B3|B I1|_XOR|B3 I1|_XOR|I_B3|MID  2e-12
II1|_XOR|I_B3|B 0 I1|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_Q1|B I1|_XOR|Q1 I1|_XOR|I_Q1|MID  2e-12
II1|_XOR|I_Q1|B 0 I1|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_XOR|A1|1 I1|_XOR|A1 I1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A1|P I1|_XOR|A1|MID_SERIES 0  5e-13
RI1|_XOR|A1|B I1|_XOR|A1 I1|_XOR|A1|MID_SHUNT  2.7439617672
LI1|_XOR|A1|RB I1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A2|1 I1|_XOR|A2 I1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A2|P I1|_XOR|A2|MID_SERIES 0  5e-13
RI1|_XOR|A2|B I1|_XOR|A2 I1|_XOR|A2|MID_SHUNT  2.7439617672
LI1|_XOR|A2|RB I1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A3|1 I1|_XOR|A2 I1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A3|P I1|_XOR|A3|MID_SERIES I1|_XOR|A3  1.2e-12
RI1|_XOR|A3|B I1|_XOR|A2 I1|_XOR|A3|MID_SHUNT  2.7439617672
LI1|_XOR|A3|RB I1|_XOR|A3|MID_SHUNT I1|_XOR|A3  2.050338398468e-12
BI1|_XOR|B1|1 I1|_XOR|B1 I1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B1|P I1|_XOR|B1|MID_SERIES 0  5e-13
RI1|_XOR|B1|B I1|_XOR|B1 I1|_XOR|B1|MID_SHUNT  2.7439617672
LI1|_XOR|B1|RB I1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B2|1 I1|_XOR|B2 I1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B2|P I1|_XOR|B2|MID_SERIES 0  5e-13
RI1|_XOR|B2|B I1|_XOR|B2 I1|_XOR|B2|MID_SHUNT  2.7439617672
LI1|_XOR|B2|RB I1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B3|1 I1|_XOR|B2 I1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B3|P I1|_XOR|B3|MID_SERIES I1|_XOR|B3  1.2e-12
RI1|_XOR|B3|B I1|_XOR|B2 I1|_XOR|B3|MID_SHUNT  2.7439617672
LI1|_XOR|B3|RB I1|_XOR|B3|MID_SHUNT I1|_XOR|B3  2.050338398468e-12
BI1|_XOR|T1|1 I1|_XOR|T1 I1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|T1|P I1|_XOR|T1|MID_SERIES 0  5e-13
RI1|_XOR|T1|B I1|_XOR|T1 I1|_XOR|T1|MID_SHUNT  2.7439617672
LI1|_XOR|T1|RB I1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|T2|1 I1|_XOR|T2 I1|_XOR|ABTQ JJMIT AREA=2.0
RI1|_XOR|T2|B I1|_XOR|T2 I1|_XOR|T2|MID_SHUNT  3.429952209
LI1|_XOR|T2|RB I1|_XOR|T2|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|AB|1 I1|_XOR|AB I1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI1|_XOR|AB|P I1|_XOR|AB|MID_SERIES I1|_XOR|ABTQ  1.2e-12
RI1|_XOR|AB|B I1|_XOR|AB I1|_XOR|AB|MID_SHUNT  3.429952209
LI1|_XOR|AB|RB I1|_XOR|AB|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|ABTQ|1 I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|ABTQ|P I1|_XOR|ABTQ|MID_SERIES 0  5e-13
RI1|_XOR|ABTQ|B I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI1|_XOR|ABTQ|RB I1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|Q1|1 I1|_XOR|Q1 I1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|Q1|P I1|_XOR|Q1|MID_SERIES 0  5e-13
RI1|_XOR|Q1|B I1|_XOR|Q1 I1|_XOR|Q1|MID_SHUNT  2.7439617672
LI1|_XOR|Q1|RB I1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI1|_AND|I_A1|B I1|_AND|A1 I1|_AND|I_A1|MID  2e-12
II1|_AND|I_A1|B 0 I1|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_B1|B I1|_AND|B1 I1|_AND|I_B1|MID  2e-12
II1|_AND|I_B1|B 0 I1|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q3|B I1|_AND|Q3 I1|_AND|I_Q3|MID  2e-12
II1|_AND|I_Q3|B 0 I1|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1|_AND|I_Q2|B I1|_AND|Q2 I1|_AND|I_Q2|MID  2e-12
II1|_AND|I_Q2|B 0 I1|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q1|B I1|_AND|Q1 I1|_AND|I_Q1|MID  2e-12
II1|_AND|I_Q1|B 0 I1|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_AND|A1|1 I1|_AND|A1 I1|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A1|P I1|_AND|A1|MID_SERIES 0  2e-13
RI1|_AND|A1|B I1|_AND|A1 I1|_AND|A1|MID_SHUNT  2.7439617672
LI1|_AND|A1|RB I1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A2|1 I1|_AND|A2 I1|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A2|P I1|_AND|A2|MID_SERIES 0  2e-13
RI1|_AND|A2|B I1|_AND|A2 I1|_AND|A2|MID_SHUNT  2.7439617672
LI1|_AND|A2|RB I1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A12|1 I1|_AND|A2 I1|_AND|A3 JJMIT AREA=1.7857142857142858
RI1|_AND|A12|B I1|_AND|A2 I1|_AND|A12|MID_SHUNT  3.84154647408
LI1|_AND|A12|RB I1|_AND|A12|MID_SHUNT I1|_AND|A3  2.1704737578552e-12
BI1|_AND|B1|1 I1|_AND|B1 I1|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B1|P I1|_AND|B1|MID_SERIES 0  2e-13
RI1|_AND|B1|B I1|_AND|B1 I1|_AND|B1|MID_SHUNT  2.7439617672
LI1|_AND|B1|RB I1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B2|1 I1|_AND|B2 I1|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B2|P I1|_AND|B2|MID_SERIES 0  2e-13
RI1|_AND|B2|B I1|_AND|B2 I1|_AND|B2|MID_SHUNT  2.7439617672
LI1|_AND|B2|RB I1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B12|1 I1|_AND|B2 I1|_AND|B3 JJMIT AREA=1.7857142857142858
RI1|_AND|B12|B I1|_AND|B2 I1|_AND|B12|MID_SHUNT  3.84154647408
LI1|_AND|B12|RB I1|_AND|B12|MID_SHUNT I1|_AND|B3  2.1704737578552e-12
BI1|_AND|Q2|1 I1|_AND|Q2 I1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q2|P I1|_AND|Q2|MID_SERIES 0  2e-13
RI1|_AND|Q2|B I1|_AND|Q2 I1|_AND|Q2|MID_SHUNT  2.7439617672
LI1|_AND|Q2|RB I1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|Q1|1 I1|_AND|Q1 I1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q1|P I1|_AND|Q1|MID_SERIES 0  2e-13
RI1|_AND|Q1|B I1|_AND|Q1 I1|_AND|Q1|MID_SHUNT  2.7439617672
LI1|_AND|Q1|RB I1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_A|I_D1|B I2|_SPL_A|D1 I2|_SPL_A|I_D1|MID  2e-12
II2|_SPL_A|I_D1|B 0 I2|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_D2|B I2|_SPL_A|D2 I2|_SPL_A|I_D2|MID  2e-12
II2|_SPL_A|I_D2|B 0 I2|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_A|I_Q1|B I2|_SPL_A|QA1 I2|_SPL_A|I_Q1|MID  2e-12
II2|_SPL_A|I_Q1|B 0 I2|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_Q2|B I2|_SPL_A|QB1 I2|_SPL_A|I_Q2|MID  2e-12
II2|_SPL_A|I_Q2|B 0 I2|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_A|1|1 I2|_SPL_A|D1 I2|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|1|P I2|_SPL_A|1|MID_SERIES 0  2e-13
RI2|_SPL_A|1|B I2|_SPL_A|D1 I2|_SPL_A|1|MID_SHUNT  2.7439617672
LI2|_SPL_A|1|RB I2|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|2|1 I2|_SPL_A|D2 I2|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|2|P I2|_SPL_A|2|MID_SERIES 0  2e-13
RI2|_SPL_A|2|B I2|_SPL_A|D2 I2|_SPL_A|2|MID_SHUNT  2.7439617672
LI2|_SPL_A|2|RB I2|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|A|1 I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|A|P I2|_SPL_A|A|MID_SERIES 0  2e-13
RI2|_SPL_A|A|B I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SHUNT  2.7439617672
LI2|_SPL_A|A|RB I2|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|B|1 I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|B|P I2|_SPL_A|B|MID_SERIES 0  2e-13
RI2|_SPL_A|B|B I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SHUNT  2.7439617672
LI2|_SPL_A|B|RB I2|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_B|I_D1|B I2|_SPL_B|D1 I2|_SPL_B|I_D1|MID  2e-12
II2|_SPL_B|I_D1|B 0 I2|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_D2|B I2|_SPL_B|D2 I2|_SPL_B|I_D2|MID  2e-12
II2|_SPL_B|I_D2|B 0 I2|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_B|I_Q1|B I2|_SPL_B|QA1 I2|_SPL_B|I_Q1|MID  2e-12
II2|_SPL_B|I_Q1|B 0 I2|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_Q2|B I2|_SPL_B|QB1 I2|_SPL_B|I_Q2|MID  2e-12
II2|_SPL_B|I_Q2|B 0 I2|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_B|1|1 I2|_SPL_B|D1 I2|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|1|P I2|_SPL_B|1|MID_SERIES 0  2e-13
RI2|_SPL_B|1|B I2|_SPL_B|D1 I2|_SPL_B|1|MID_SHUNT  2.7439617672
LI2|_SPL_B|1|RB I2|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|2|1 I2|_SPL_B|D2 I2|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|2|P I2|_SPL_B|2|MID_SERIES 0  2e-13
RI2|_SPL_B|2|B I2|_SPL_B|D2 I2|_SPL_B|2|MID_SHUNT  2.7439617672
LI2|_SPL_B|2|RB I2|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|A|1 I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|A|P I2|_SPL_B|A|MID_SERIES 0  2e-13
RI2|_SPL_B|A|B I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SHUNT  2.7439617672
LI2|_SPL_B|A|RB I2|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|B|1 I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|B|P I2|_SPL_B|B|MID_SERIES 0  2e-13
RI2|_SPL_B|B|B I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SHUNT  2.7439617672
LI2|_SPL_B|B|RB I2|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_A|I_1|B I2|_DFF_A|A1 I2|_DFF_A|I_1|MID  2e-12
II2|_DFF_A|I_1|B 0 I2|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_3|B I2|_DFF_A|A3 I2|_DFF_A|I_3|MID  2e-12
II2|_DFF_A|I_3|B 0 I2|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_A|I_T|B I2|_DFF_A|T1 I2|_DFF_A|I_T|MID  2e-12
II2|_DFF_A|I_T|B 0 I2|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_6|B I2|_DFF_A|Q1 I2|_DFF_A|I_6|MID  2e-12
II2|_DFF_A|I_6|B 0 I2|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_A|1|1 I2|_DFF_A|A1 I2|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|1|P I2|_DFF_A|1|MID_SERIES 0  2e-13
RI2|_DFF_A|1|B I2|_DFF_A|A1 I2|_DFF_A|1|MID_SHUNT  2.7439617672
LI2|_DFF_A|1|RB I2|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|23|1 I2|_DFF_A|A2 I2|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|23|B I2|_DFF_A|A2 I2|_DFF_A|23|MID_SHUNT  3.84154647408
LI2|_DFF_A|23|RB I2|_DFF_A|23|MID_SHUNT I2|_DFF_A|A3  2.1704737578552e-12
BI2|_DFF_A|3|1 I2|_DFF_A|A3 I2|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|3|P I2|_DFF_A|3|MID_SERIES 0  2e-13
RI2|_DFF_A|3|B I2|_DFF_A|A3 I2|_DFF_A|3|MID_SHUNT  2.7439617672
LI2|_DFF_A|3|RB I2|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|4|1 I2|_DFF_A|A4 I2|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|4|P I2|_DFF_A|4|MID_SERIES 0  2e-13
RI2|_DFF_A|4|B I2|_DFF_A|A4 I2|_DFF_A|4|MID_SHUNT  2.7439617672
LI2|_DFF_A|4|RB I2|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|T|1 I2|_DFF_A|T1 I2|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|T|P I2|_DFF_A|T|MID_SERIES 0  2e-13
RI2|_DFF_A|T|B I2|_DFF_A|T1 I2|_DFF_A|T|MID_SHUNT  2.7439617672
LI2|_DFF_A|T|RB I2|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|45|1 I2|_DFF_A|T2 I2|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|45|B I2|_DFF_A|T2 I2|_DFF_A|45|MID_SHUNT  3.84154647408
LI2|_DFF_A|45|RB I2|_DFF_A|45|MID_SHUNT I2|_DFF_A|A4  2.1704737578552e-12
BI2|_DFF_A|6|1 I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|6|P I2|_DFF_A|6|MID_SERIES 0  2e-13
RI2|_DFF_A|6|B I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SHUNT  2.7439617672
LI2|_DFF_A|6|RB I2|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_B|I_1|B I2|_DFF_B|A1 I2|_DFF_B|I_1|MID  2e-12
II2|_DFF_B|I_1|B 0 I2|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_3|B I2|_DFF_B|A3 I2|_DFF_B|I_3|MID  2e-12
II2|_DFF_B|I_3|B 0 I2|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_B|I_T|B I2|_DFF_B|T1 I2|_DFF_B|I_T|MID  2e-12
II2|_DFF_B|I_T|B 0 I2|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_6|B I2|_DFF_B|Q1 I2|_DFF_B|I_6|MID  2e-12
II2|_DFF_B|I_6|B 0 I2|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_B|1|1 I2|_DFF_B|A1 I2|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|1|P I2|_DFF_B|1|MID_SERIES 0  2e-13
RI2|_DFF_B|1|B I2|_DFF_B|A1 I2|_DFF_B|1|MID_SHUNT  2.7439617672
LI2|_DFF_B|1|RB I2|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|23|1 I2|_DFF_B|A2 I2|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|23|B I2|_DFF_B|A2 I2|_DFF_B|23|MID_SHUNT  3.84154647408
LI2|_DFF_B|23|RB I2|_DFF_B|23|MID_SHUNT I2|_DFF_B|A3  2.1704737578552e-12
BI2|_DFF_B|3|1 I2|_DFF_B|A3 I2|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|3|P I2|_DFF_B|3|MID_SERIES 0  2e-13
RI2|_DFF_B|3|B I2|_DFF_B|A3 I2|_DFF_B|3|MID_SHUNT  2.7439617672
LI2|_DFF_B|3|RB I2|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|4|1 I2|_DFF_B|A4 I2|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|4|P I2|_DFF_B|4|MID_SERIES 0  2e-13
RI2|_DFF_B|4|B I2|_DFF_B|A4 I2|_DFF_B|4|MID_SHUNT  2.7439617672
LI2|_DFF_B|4|RB I2|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|T|1 I2|_DFF_B|T1 I2|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|T|P I2|_DFF_B|T|MID_SERIES 0  2e-13
RI2|_DFF_B|T|B I2|_DFF_B|T1 I2|_DFF_B|T|MID_SHUNT  2.7439617672
LI2|_DFF_B|T|RB I2|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|45|1 I2|_DFF_B|T2 I2|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|45|B I2|_DFF_B|T2 I2|_DFF_B|45|MID_SHUNT  3.84154647408
LI2|_DFF_B|45|RB I2|_DFF_B|45|MID_SHUNT I2|_DFF_B|A4  2.1704737578552e-12
BI2|_DFF_B|6|1 I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|6|P I2|_DFF_B|6|MID_SERIES 0  2e-13
RI2|_DFF_B|6|B I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SHUNT  2.7439617672
LI2|_DFF_B|6|RB I2|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI2|_XOR|I_A1|B I2|_XOR|A1 I2|_XOR|I_A1|MID  2e-12
II2|_XOR|I_A1|B 0 I2|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_A3|B I2|_XOR|A3 I2|_XOR|I_A3|MID  2e-12
II2|_XOR|I_A3|B 0 I2|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B1|B I2|_XOR|B1 I2|_XOR|I_B1|MID  2e-12
II2|_XOR|I_B1|B 0 I2|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B3|B I2|_XOR|B3 I2|_XOR|I_B3|MID  2e-12
II2|_XOR|I_B3|B 0 I2|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_Q1|B I2|_XOR|Q1 I2|_XOR|I_Q1|MID  2e-12
II2|_XOR|I_Q1|B 0 I2|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_XOR|A1|1 I2|_XOR|A1 I2|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A1|P I2|_XOR|A1|MID_SERIES 0  5e-13
RI2|_XOR|A1|B I2|_XOR|A1 I2|_XOR|A1|MID_SHUNT  2.7439617672
LI2|_XOR|A1|RB I2|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A2|1 I2|_XOR|A2 I2|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A2|P I2|_XOR|A2|MID_SERIES 0  5e-13
RI2|_XOR|A2|B I2|_XOR|A2 I2|_XOR|A2|MID_SHUNT  2.7439617672
LI2|_XOR|A2|RB I2|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A3|1 I2|_XOR|A2 I2|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A3|P I2|_XOR|A3|MID_SERIES I2|_XOR|A3  1.2e-12
RI2|_XOR|A3|B I2|_XOR|A2 I2|_XOR|A3|MID_SHUNT  2.7439617672
LI2|_XOR|A3|RB I2|_XOR|A3|MID_SHUNT I2|_XOR|A3  2.050338398468e-12
BI2|_XOR|B1|1 I2|_XOR|B1 I2|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B1|P I2|_XOR|B1|MID_SERIES 0  5e-13
RI2|_XOR|B1|B I2|_XOR|B1 I2|_XOR|B1|MID_SHUNT  2.7439617672
LI2|_XOR|B1|RB I2|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B2|1 I2|_XOR|B2 I2|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B2|P I2|_XOR|B2|MID_SERIES 0  5e-13
RI2|_XOR|B2|B I2|_XOR|B2 I2|_XOR|B2|MID_SHUNT  2.7439617672
LI2|_XOR|B2|RB I2|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B3|1 I2|_XOR|B2 I2|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B3|P I2|_XOR|B3|MID_SERIES I2|_XOR|B3  1.2e-12
RI2|_XOR|B3|B I2|_XOR|B2 I2|_XOR|B3|MID_SHUNT  2.7439617672
LI2|_XOR|B3|RB I2|_XOR|B3|MID_SHUNT I2|_XOR|B3  2.050338398468e-12
BI2|_XOR|T1|1 I2|_XOR|T1 I2|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|T1|P I2|_XOR|T1|MID_SERIES 0  5e-13
RI2|_XOR|T1|B I2|_XOR|T1 I2|_XOR|T1|MID_SHUNT  2.7439617672
LI2|_XOR|T1|RB I2|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|T2|1 I2|_XOR|T2 I2|_XOR|ABTQ JJMIT AREA=2.0
RI2|_XOR|T2|B I2|_XOR|T2 I2|_XOR|T2|MID_SHUNT  3.429952209
LI2|_XOR|T2|RB I2|_XOR|T2|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|AB|1 I2|_XOR|AB I2|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI2|_XOR|AB|P I2|_XOR|AB|MID_SERIES I2|_XOR|ABTQ  1.2e-12
RI2|_XOR|AB|B I2|_XOR|AB I2|_XOR|AB|MID_SHUNT  3.429952209
LI2|_XOR|AB|RB I2|_XOR|AB|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|ABTQ|1 I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|ABTQ|P I2|_XOR|ABTQ|MID_SERIES 0  5e-13
RI2|_XOR|ABTQ|B I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI2|_XOR|ABTQ|RB I2|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|Q1|1 I2|_XOR|Q1 I2|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|Q1|P I2|_XOR|Q1|MID_SERIES 0  5e-13
RI2|_XOR|Q1|B I2|_XOR|Q1 I2|_XOR|Q1|MID_SHUNT  2.7439617672
LI2|_XOR|Q1|RB I2|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI2|_AND|I_A1|B I2|_AND|A1 I2|_AND|I_A1|MID  2e-12
II2|_AND|I_A1|B 0 I2|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_B1|B I2|_AND|B1 I2|_AND|I_B1|MID  2e-12
II2|_AND|I_B1|B 0 I2|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q3|B I2|_AND|Q3 I2|_AND|I_Q3|MID  2e-12
II2|_AND|I_Q3|B 0 I2|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2|_AND|I_Q2|B I2|_AND|Q2 I2|_AND|I_Q2|MID  2e-12
II2|_AND|I_Q2|B 0 I2|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q1|B I2|_AND|Q1 I2|_AND|I_Q1|MID  2e-12
II2|_AND|I_Q1|B 0 I2|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_AND|A1|1 I2|_AND|A1 I2|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A1|P I2|_AND|A1|MID_SERIES 0  2e-13
RI2|_AND|A1|B I2|_AND|A1 I2|_AND|A1|MID_SHUNT  2.7439617672
LI2|_AND|A1|RB I2|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A2|1 I2|_AND|A2 I2|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A2|P I2|_AND|A2|MID_SERIES 0  2e-13
RI2|_AND|A2|B I2|_AND|A2 I2|_AND|A2|MID_SHUNT  2.7439617672
LI2|_AND|A2|RB I2|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A12|1 I2|_AND|A2 I2|_AND|A3 JJMIT AREA=1.7857142857142858
RI2|_AND|A12|B I2|_AND|A2 I2|_AND|A12|MID_SHUNT  3.84154647408
LI2|_AND|A12|RB I2|_AND|A12|MID_SHUNT I2|_AND|A3  2.1704737578552e-12
BI2|_AND|B1|1 I2|_AND|B1 I2|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B1|P I2|_AND|B1|MID_SERIES 0  2e-13
RI2|_AND|B1|B I2|_AND|B1 I2|_AND|B1|MID_SHUNT  2.7439617672
LI2|_AND|B1|RB I2|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B2|1 I2|_AND|B2 I2|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B2|P I2|_AND|B2|MID_SERIES 0  2e-13
RI2|_AND|B2|B I2|_AND|B2 I2|_AND|B2|MID_SHUNT  2.7439617672
LI2|_AND|B2|RB I2|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B12|1 I2|_AND|B2 I2|_AND|B3 JJMIT AREA=1.7857142857142858
RI2|_AND|B12|B I2|_AND|B2 I2|_AND|B12|MID_SHUNT  3.84154647408
LI2|_AND|B12|RB I2|_AND|B12|MID_SHUNT I2|_AND|B3  2.1704737578552e-12
BI2|_AND|Q2|1 I2|_AND|Q2 I2|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q2|P I2|_AND|Q2|MID_SERIES 0  2e-13
RI2|_AND|Q2|B I2|_AND|Q2 I2|_AND|Q2|MID_SHUNT  2.7439617672
LI2|_AND|Q2|RB I2|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|Q1|1 I2|_AND|Q1 I2|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q1|P I2|_AND|Q1|MID_SERIES 0  2e-13
RI2|_AND|Q1|B I2|_AND|Q1 I2|_AND|Q1|MID_SHUNT  2.7439617672
LI2|_AND|Q1|RB I2|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_A|I_D1|B I3|_SPL_A|D1 I3|_SPL_A|I_D1|MID  2e-12
II3|_SPL_A|I_D1|B 0 I3|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_D2|B I3|_SPL_A|D2 I3|_SPL_A|I_D2|MID  2e-12
II3|_SPL_A|I_D2|B 0 I3|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_A|I_Q1|B I3|_SPL_A|QA1 I3|_SPL_A|I_Q1|MID  2e-12
II3|_SPL_A|I_Q1|B 0 I3|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_Q2|B I3|_SPL_A|QB1 I3|_SPL_A|I_Q2|MID  2e-12
II3|_SPL_A|I_Q2|B 0 I3|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_A|1|1 I3|_SPL_A|D1 I3|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|1|P I3|_SPL_A|1|MID_SERIES 0  2e-13
RI3|_SPL_A|1|B I3|_SPL_A|D1 I3|_SPL_A|1|MID_SHUNT  2.7439617672
LI3|_SPL_A|1|RB I3|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|2|1 I3|_SPL_A|D2 I3|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|2|P I3|_SPL_A|2|MID_SERIES 0  2e-13
RI3|_SPL_A|2|B I3|_SPL_A|D2 I3|_SPL_A|2|MID_SHUNT  2.7439617672
LI3|_SPL_A|2|RB I3|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|A|1 I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|A|P I3|_SPL_A|A|MID_SERIES 0  2e-13
RI3|_SPL_A|A|B I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SHUNT  2.7439617672
LI3|_SPL_A|A|RB I3|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|B|1 I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|B|P I3|_SPL_A|B|MID_SERIES 0  2e-13
RI3|_SPL_A|B|B I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SHUNT  2.7439617672
LI3|_SPL_A|B|RB I3|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_B|I_D1|B I3|_SPL_B|D1 I3|_SPL_B|I_D1|MID  2e-12
II3|_SPL_B|I_D1|B 0 I3|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_D2|B I3|_SPL_B|D2 I3|_SPL_B|I_D2|MID  2e-12
II3|_SPL_B|I_D2|B 0 I3|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_B|I_Q1|B I3|_SPL_B|QA1 I3|_SPL_B|I_Q1|MID  2e-12
II3|_SPL_B|I_Q1|B 0 I3|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_Q2|B I3|_SPL_B|QB1 I3|_SPL_B|I_Q2|MID  2e-12
II3|_SPL_B|I_Q2|B 0 I3|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_B|1|1 I3|_SPL_B|D1 I3|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|1|P I3|_SPL_B|1|MID_SERIES 0  2e-13
RI3|_SPL_B|1|B I3|_SPL_B|D1 I3|_SPL_B|1|MID_SHUNT  2.7439617672
LI3|_SPL_B|1|RB I3|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|2|1 I3|_SPL_B|D2 I3|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|2|P I3|_SPL_B|2|MID_SERIES 0  2e-13
RI3|_SPL_B|2|B I3|_SPL_B|D2 I3|_SPL_B|2|MID_SHUNT  2.7439617672
LI3|_SPL_B|2|RB I3|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|A|1 I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|A|P I3|_SPL_B|A|MID_SERIES 0  2e-13
RI3|_SPL_B|A|B I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SHUNT  2.7439617672
LI3|_SPL_B|A|RB I3|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|B|1 I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|B|P I3|_SPL_B|B|MID_SERIES 0  2e-13
RI3|_SPL_B|B|B I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SHUNT  2.7439617672
LI3|_SPL_B|B|RB I3|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_A|I_1|B I3|_DFF_A|A1 I3|_DFF_A|I_1|MID  2e-12
II3|_DFF_A|I_1|B 0 I3|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_3|B I3|_DFF_A|A3 I3|_DFF_A|I_3|MID  2e-12
II3|_DFF_A|I_3|B 0 I3|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_A|I_T|B I3|_DFF_A|T1 I3|_DFF_A|I_T|MID  2e-12
II3|_DFF_A|I_T|B 0 I3|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_6|B I3|_DFF_A|Q1 I3|_DFF_A|I_6|MID  2e-12
II3|_DFF_A|I_6|B 0 I3|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_A|1|1 I3|_DFF_A|A1 I3|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|1|P I3|_DFF_A|1|MID_SERIES 0  2e-13
RI3|_DFF_A|1|B I3|_DFF_A|A1 I3|_DFF_A|1|MID_SHUNT  2.7439617672
LI3|_DFF_A|1|RB I3|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|23|1 I3|_DFF_A|A2 I3|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|23|B I3|_DFF_A|A2 I3|_DFF_A|23|MID_SHUNT  3.84154647408
LI3|_DFF_A|23|RB I3|_DFF_A|23|MID_SHUNT I3|_DFF_A|A3  2.1704737578552e-12
BI3|_DFF_A|3|1 I3|_DFF_A|A3 I3|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|3|P I3|_DFF_A|3|MID_SERIES 0  2e-13
RI3|_DFF_A|3|B I3|_DFF_A|A3 I3|_DFF_A|3|MID_SHUNT  2.7439617672
LI3|_DFF_A|3|RB I3|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|4|1 I3|_DFF_A|A4 I3|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|4|P I3|_DFF_A|4|MID_SERIES 0  2e-13
RI3|_DFF_A|4|B I3|_DFF_A|A4 I3|_DFF_A|4|MID_SHUNT  2.7439617672
LI3|_DFF_A|4|RB I3|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|T|1 I3|_DFF_A|T1 I3|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|T|P I3|_DFF_A|T|MID_SERIES 0  2e-13
RI3|_DFF_A|T|B I3|_DFF_A|T1 I3|_DFF_A|T|MID_SHUNT  2.7439617672
LI3|_DFF_A|T|RB I3|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|45|1 I3|_DFF_A|T2 I3|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|45|B I3|_DFF_A|T2 I3|_DFF_A|45|MID_SHUNT  3.84154647408
LI3|_DFF_A|45|RB I3|_DFF_A|45|MID_SHUNT I3|_DFF_A|A4  2.1704737578552e-12
BI3|_DFF_A|6|1 I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|6|P I3|_DFF_A|6|MID_SERIES 0  2e-13
RI3|_DFF_A|6|B I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SHUNT  2.7439617672
LI3|_DFF_A|6|RB I3|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_B|I_1|B I3|_DFF_B|A1 I3|_DFF_B|I_1|MID  2e-12
II3|_DFF_B|I_1|B 0 I3|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_3|B I3|_DFF_B|A3 I3|_DFF_B|I_3|MID  2e-12
II3|_DFF_B|I_3|B 0 I3|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_B|I_T|B I3|_DFF_B|T1 I3|_DFF_B|I_T|MID  2e-12
II3|_DFF_B|I_T|B 0 I3|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_6|B I3|_DFF_B|Q1 I3|_DFF_B|I_6|MID  2e-12
II3|_DFF_B|I_6|B 0 I3|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_B|1|1 I3|_DFF_B|A1 I3|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|1|P I3|_DFF_B|1|MID_SERIES 0  2e-13
RI3|_DFF_B|1|B I3|_DFF_B|A1 I3|_DFF_B|1|MID_SHUNT  2.7439617672
LI3|_DFF_B|1|RB I3|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|23|1 I3|_DFF_B|A2 I3|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|23|B I3|_DFF_B|A2 I3|_DFF_B|23|MID_SHUNT  3.84154647408
LI3|_DFF_B|23|RB I3|_DFF_B|23|MID_SHUNT I3|_DFF_B|A3  2.1704737578552e-12
BI3|_DFF_B|3|1 I3|_DFF_B|A3 I3|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|3|P I3|_DFF_B|3|MID_SERIES 0  2e-13
RI3|_DFF_B|3|B I3|_DFF_B|A3 I3|_DFF_B|3|MID_SHUNT  2.7439617672
LI3|_DFF_B|3|RB I3|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|4|1 I3|_DFF_B|A4 I3|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|4|P I3|_DFF_B|4|MID_SERIES 0  2e-13
RI3|_DFF_B|4|B I3|_DFF_B|A4 I3|_DFF_B|4|MID_SHUNT  2.7439617672
LI3|_DFF_B|4|RB I3|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|T|1 I3|_DFF_B|T1 I3|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|T|P I3|_DFF_B|T|MID_SERIES 0  2e-13
RI3|_DFF_B|T|B I3|_DFF_B|T1 I3|_DFF_B|T|MID_SHUNT  2.7439617672
LI3|_DFF_B|T|RB I3|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|45|1 I3|_DFF_B|T2 I3|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|45|B I3|_DFF_B|T2 I3|_DFF_B|45|MID_SHUNT  3.84154647408
LI3|_DFF_B|45|RB I3|_DFF_B|45|MID_SHUNT I3|_DFF_B|A4  2.1704737578552e-12
BI3|_DFF_B|6|1 I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|6|P I3|_DFF_B|6|MID_SERIES 0  2e-13
RI3|_DFF_B|6|B I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SHUNT  2.7439617672
LI3|_DFF_B|6|RB I3|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI3|_XOR|I_A1|B I3|_XOR|A1 I3|_XOR|I_A1|MID  2e-12
II3|_XOR|I_A1|B 0 I3|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_A3|B I3|_XOR|A3 I3|_XOR|I_A3|MID  2e-12
II3|_XOR|I_A3|B 0 I3|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B1|B I3|_XOR|B1 I3|_XOR|I_B1|MID  2e-12
II3|_XOR|I_B1|B 0 I3|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B3|B I3|_XOR|B3 I3|_XOR|I_B3|MID  2e-12
II3|_XOR|I_B3|B 0 I3|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_Q1|B I3|_XOR|Q1 I3|_XOR|I_Q1|MID  2e-12
II3|_XOR|I_Q1|B 0 I3|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_XOR|A1|1 I3|_XOR|A1 I3|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A1|P I3|_XOR|A1|MID_SERIES 0  5e-13
RI3|_XOR|A1|B I3|_XOR|A1 I3|_XOR|A1|MID_SHUNT  2.7439617672
LI3|_XOR|A1|RB I3|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A2|1 I3|_XOR|A2 I3|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A2|P I3|_XOR|A2|MID_SERIES 0  5e-13
RI3|_XOR|A2|B I3|_XOR|A2 I3|_XOR|A2|MID_SHUNT  2.7439617672
LI3|_XOR|A2|RB I3|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A3|1 I3|_XOR|A2 I3|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A3|P I3|_XOR|A3|MID_SERIES I3|_XOR|A3  1.2e-12
RI3|_XOR|A3|B I3|_XOR|A2 I3|_XOR|A3|MID_SHUNT  2.7439617672
LI3|_XOR|A3|RB I3|_XOR|A3|MID_SHUNT I3|_XOR|A3  2.050338398468e-12
BI3|_XOR|B1|1 I3|_XOR|B1 I3|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B1|P I3|_XOR|B1|MID_SERIES 0  5e-13
RI3|_XOR|B1|B I3|_XOR|B1 I3|_XOR|B1|MID_SHUNT  2.7439617672
LI3|_XOR|B1|RB I3|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B2|1 I3|_XOR|B2 I3|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B2|P I3|_XOR|B2|MID_SERIES 0  5e-13
RI3|_XOR|B2|B I3|_XOR|B2 I3|_XOR|B2|MID_SHUNT  2.7439617672
LI3|_XOR|B2|RB I3|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B3|1 I3|_XOR|B2 I3|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B3|P I3|_XOR|B3|MID_SERIES I3|_XOR|B3  1.2e-12
RI3|_XOR|B3|B I3|_XOR|B2 I3|_XOR|B3|MID_SHUNT  2.7439617672
LI3|_XOR|B3|RB I3|_XOR|B3|MID_SHUNT I3|_XOR|B3  2.050338398468e-12
BI3|_XOR|T1|1 I3|_XOR|T1 I3|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|T1|P I3|_XOR|T1|MID_SERIES 0  5e-13
RI3|_XOR|T1|B I3|_XOR|T1 I3|_XOR|T1|MID_SHUNT  2.7439617672
LI3|_XOR|T1|RB I3|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|T2|1 I3|_XOR|T2 I3|_XOR|ABTQ JJMIT AREA=2.0
RI3|_XOR|T2|B I3|_XOR|T2 I3|_XOR|T2|MID_SHUNT  3.429952209
LI3|_XOR|T2|RB I3|_XOR|T2|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|AB|1 I3|_XOR|AB I3|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI3|_XOR|AB|P I3|_XOR|AB|MID_SERIES I3|_XOR|ABTQ  1.2e-12
RI3|_XOR|AB|B I3|_XOR|AB I3|_XOR|AB|MID_SHUNT  3.429952209
LI3|_XOR|AB|RB I3|_XOR|AB|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|ABTQ|1 I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|ABTQ|P I3|_XOR|ABTQ|MID_SERIES 0  5e-13
RI3|_XOR|ABTQ|B I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI3|_XOR|ABTQ|RB I3|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|Q1|1 I3|_XOR|Q1 I3|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|Q1|P I3|_XOR|Q1|MID_SERIES 0  5e-13
RI3|_XOR|Q1|B I3|_XOR|Q1 I3|_XOR|Q1|MID_SHUNT  2.7439617672
LI3|_XOR|Q1|RB I3|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI3|_AND|I_A1|B I3|_AND|A1 I3|_AND|I_A1|MID  2e-12
II3|_AND|I_A1|B 0 I3|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_B1|B I3|_AND|B1 I3|_AND|I_B1|MID  2e-12
II3|_AND|I_B1|B 0 I3|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q3|B I3|_AND|Q3 I3|_AND|I_Q3|MID  2e-12
II3|_AND|I_Q3|B 0 I3|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3|_AND|I_Q2|B I3|_AND|Q2 I3|_AND|I_Q2|MID  2e-12
II3|_AND|I_Q2|B 0 I3|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q1|B I3|_AND|Q1 I3|_AND|I_Q1|MID  2e-12
II3|_AND|I_Q1|B 0 I3|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_AND|A1|1 I3|_AND|A1 I3|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A1|P I3|_AND|A1|MID_SERIES 0  2e-13
RI3|_AND|A1|B I3|_AND|A1 I3|_AND|A1|MID_SHUNT  2.7439617672
LI3|_AND|A1|RB I3|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A2|1 I3|_AND|A2 I3|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A2|P I3|_AND|A2|MID_SERIES 0  2e-13
RI3|_AND|A2|B I3|_AND|A2 I3|_AND|A2|MID_SHUNT  2.7439617672
LI3|_AND|A2|RB I3|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A12|1 I3|_AND|A2 I3|_AND|A3 JJMIT AREA=1.7857142857142858
RI3|_AND|A12|B I3|_AND|A2 I3|_AND|A12|MID_SHUNT  3.84154647408
LI3|_AND|A12|RB I3|_AND|A12|MID_SHUNT I3|_AND|A3  2.1704737578552e-12
BI3|_AND|B1|1 I3|_AND|B1 I3|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B1|P I3|_AND|B1|MID_SERIES 0  2e-13
RI3|_AND|B1|B I3|_AND|B1 I3|_AND|B1|MID_SHUNT  2.7439617672
LI3|_AND|B1|RB I3|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B2|1 I3|_AND|B2 I3|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B2|P I3|_AND|B2|MID_SERIES 0  2e-13
RI3|_AND|B2|B I3|_AND|B2 I3|_AND|B2|MID_SHUNT  2.7439617672
LI3|_AND|B2|RB I3|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B12|1 I3|_AND|B2 I3|_AND|B3 JJMIT AREA=1.7857142857142858
RI3|_AND|B12|B I3|_AND|B2 I3|_AND|B12|MID_SHUNT  3.84154647408
LI3|_AND|B12|RB I3|_AND|B12|MID_SHUNT I3|_AND|B3  2.1704737578552e-12
BI3|_AND|Q2|1 I3|_AND|Q2 I3|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q2|P I3|_AND|Q2|MID_SERIES 0  2e-13
RI3|_AND|Q2|B I3|_AND|Q2 I3|_AND|Q2|MID_SHUNT  2.7439617672
LI3|_AND|Q2|RB I3|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|Q1|1 I3|_AND|Q1 I3|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q1|P I3|_AND|Q1|MID_SERIES 0  2e-13
RI3|_AND|Q1|B I3|_AND|Q1 I3|_AND|Q1|MID_SHUNT  2.7439617672
LI3|_AND|Q1|RB I3|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|I_D1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|I_D1|MID  2e-12
ISPL_IP2_0|SPL1|I_D1|B 0 SPL_IP2_0|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL1|I_D2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|I_D2|MID  2e-12
ISPL_IP2_0|SPL1|I_D2|B 0 SPL_IP2_0|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_IP2_0|SPL1|I_Q1|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|I_Q1|MID  2e-12
ISPL_IP2_0|SPL1|I_Q1|B 0 SPL_IP2_0|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL1|I_Q2|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|I_Q2|MID  2e-12
ISPL_IP2_0|SPL1|I_Q2|B 0 SPL_IP2_0|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_IP2_0|SPL1|1|1 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|1|P SPL_IP2_0|SPL1|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|1|RB SPL_IP2_0|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|2|1 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|2|P SPL_IP2_0|SPL1|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|2|RB SPL_IP2_0|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|A|1 SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|A|P SPL_IP2_0|SPL1|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|A|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|A|RB SPL_IP2_0|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|B|1 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|B|P SPL_IP2_0|SPL1|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|B|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|B|RB SPL_IP2_0|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL2|I_D1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|I_D1|MID  2e-12
ISPL_IP2_0|SPL2|I_D1|B 0 SPL_IP2_0|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL2|I_D2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|I_D2|MID  2e-12
ISPL_IP2_0|SPL2|I_D2|B 0 SPL_IP2_0|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_IP2_0|SPL2|I_Q1|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|I_Q1|MID  2e-12
ISPL_IP2_0|SPL2|I_Q1|B 0 SPL_IP2_0|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL2|I_Q2|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|I_Q2|MID  2e-12
ISPL_IP2_0|SPL2|I_Q2|B 0 SPL_IP2_0|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_IP2_0|SPL2|1|1 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|1|P SPL_IP2_0|SPL2|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|1|RB SPL_IP2_0|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|2|1 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|2|P SPL_IP2_0|SPL2|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|2|RB SPL_IP2_0|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|A|1 SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|A|P SPL_IP2_0|SPL2|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|A|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|A|RB SPL_IP2_0|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|B|1 SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|B|P SPL_IP2_0|SPL2|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|B|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|B|RB SPL_IP2_0|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|I_1|B _PG0_01|P|A1 _PG0_01|P|I_1|MID  2e-12
I_PG0_01|P|I_1|B 0 _PG0_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_3|B _PG0_01|P|A3 _PG0_01|P|I_3|MID  2e-12
I_PG0_01|P|I_3|B 0 _PG0_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|P|I_T|B _PG0_01|P|T1 _PG0_01|P|I_T|MID  2e-12
I_PG0_01|P|I_T|B 0 _PG0_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_6|B _PG0_01|P|Q1 _PG0_01|P|I_6|MID  2e-12
I_PG0_01|P|I_6|B 0 _PG0_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|P|1|1 _PG0_01|P|A1 _PG0_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|1|P _PG0_01|P|1|MID_SERIES 0  2e-13
R_PG0_01|P|1|B _PG0_01|P|A1 _PG0_01|P|1|MID_SHUNT  2.7439617672
L_PG0_01|P|1|RB _PG0_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|23|1 _PG0_01|P|A2 _PG0_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|P|23|B _PG0_01|P|A2 _PG0_01|P|23|MID_SHUNT  3.84154647408
L_PG0_01|P|23|RB _PG0_01|P|23|MID_SHUNT _PG0_01|P|A3  2.1704737578552e-12
B_PG0_01|P|3|1 _PG0_01|P|A3 _PG0_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|3|P _PG0_01|P|3|MID_SERIES 0  2e-13
R_PG0_01|P|3|B _PG0_01|P|A3 _PG0_01|P|3|MID_SHUNT  2.7439617672
L_PG0_01|P|3|RB _PG0_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|4|1 _PG0_01|P|A4 _PG0_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|4|P _PG0_01|P|4|MID_SERIES 0  2e-13
R_PG0_01|P|4|B _PG0_01|P|A4 _PG0_01|P|4|MID_SHUNT  2.7439617672
L_PG0_01|P|4|RB _PG0_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|T|1 _PG0_01|P|T1 _PG0_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|T|P _PG0_01|P|T|MID_SERIES 0  2e-13
R_PG0_01|P|T|B _PG0_01|P|T1 _PG0_01|P|T|MID_SHUNT  2.7439617672
L_PG0_01|P|T|RB _PG0_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|45|1 _PG0_01|P|T2 _PG0_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|P|45|B _PG0_01|P|T2 _PG0_01|P|45|MID_SHUNT  3.84154647408
L_PG0_01|P|45|RB _PG0_01|P|45|MID_SHUNT _PG0_01|P|A4  2.1704737578552e-12
B_PG0_01|P|6|1 _PG0_01|P|Q1 _PG0_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|6|P _PG0_01|P|6|MID_SERIES 0  2e-13
R_PG0_01|P|6|B _PG0_01|P|Q1 _PG0_01|P|6|MID_SHUNT  2.7439617672
L_PG0_01|P|6|RB _PG0_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|G|I_1|B _PG0_01|G|A1 _PG0_01|G|I_1|MID  2e-12
I_PG0_01|G|I_1|B 0 _PG0_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_3|B _PG0_01|G|A3 _PG0_01|G|I_3|MID  2e-12
I_PG0_01|G|I_3|B 0 _PG0_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|G|I_T|B _PG0_01|G|T1 _PG0_01|G|I_T|MID  2e-12
I_PG0_01|G|I_T|B 0 _PG0_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_6|B _PG0_01|G|Q1 _PG0_01|G|I_6|MID  2e-12
I_PG0_01|G|I_6|B 0 _PG0_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|G|1|1 _PG0_01|G|A1 _PG0_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|1|P _PG0_01|G|1|MID_SERIES 0  2e-13
R_PG0_01|G|1|B _PG0_01|G|A1 _PG0_01|G|1|MID_SHUNT  2.7439617672
L_PG0_01|G|1|RB _PG0_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|23|1 _PG0_01|G|A2 _PG0_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|G|23|B _PG0_01|G|A2 _PG0_01|G|23|MID_SHUNT  3.84154647408
L_PG0_01|G|23|RB _PG0_01|G|23|MID_SHUNT _PG0_01|G|A3  2.1704737578552e-12
B_PG0_01|G|3|1 _PG0_01|G|A3 _PG0_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|3|P _PG0_01|G|3|MID_SERIES 0  2e-13
R_PG0_01|G|3|B _PG0_01|G|A3 _PG0_01|G|3|MID_SHUNT  2.7439617672
L_PG0_01|G|3|RB _PG0_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|4|1 _PG0_01|G|A4 _PG0_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|4|P _PG0_01|G|4|MID_SERIES 0  2e-13
R_PG0_01|G|4|B _PG0_01|G|A4 _PG0_01|G|4|MID_SHUNT  2.7439617672
L_PG0_01|G|4|RB _PG0_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|T|1 _PG0_01|G|T1 _PG0_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|T|P _PG0_01|G|T|MID_SERIES 0  2e-13
R_PG0_01|G|T|B _PG0_01|G|T1 _PG0_01|G|T|MID_SHUNT  2.7439617672
L_PG0_01|G|T|RB _PG0_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|45|1 _PG0_01|G|T2 _PG0_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|G|45|B _PG0_01|G|T2 _PG0_01|G|45|MID_SHUNT  3.84154647408
L_PG0_01|G|45|RB _PG0_01|G|45|MID_SHUNT _PG0_01|G|A4  2.1704737578552e-12
B_PG0_01|G|6|1 _PG0_01|G|Q1 _PG0_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|6|P _PG0_01|G|6|MID_SERIES 0  2e-13
R_PG0_01|G|6|B _PG0_01|G|Q1 _PG0_01|G|6|MID_SHUNT  2.7439617672
L_PG0_01|G|6|RB _PG0_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_SPL_G1|I_D1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|I_D1|MID  2e-12
I_PG1_01|_SPL_G1|I_D1|B 0 _PG1_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_D2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|I_D2|MID  2e-12
I_PG1_01|_SPL_G1|I_D2|B 0 _PG1_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG1_01|_SPL_G1|I_Q1|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|I_Q1|MID  2e-12
I_PG1_01|_SPL_G1|I_Q1|B 0 _PG1_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_Q2|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|I_Q2|MID  2e-12
I_PG1_01|_SPL_G1|I_Q2|B 0 _PG1_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG1_01|_SPL_G1|1|1 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|1|P _PG1_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|1|RB _PG1_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|2|1 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|2|P _PG1_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|2|RB _PG1_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|A|1 _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|A|P _PG1_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|A|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|A|RB _PG1_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|B|1 _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|B|P _PG1_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|B|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|B|RB _PG1_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_PG|I_A1|B _PG1_01|_PG|A1 _PG1_01|_PG|I_A1|MID  2e-12
I_PG1_01|_PG|I_A1|B 0 _PG1_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_B1|B _PG1_01|_PG|B1 _PG1_01|_PG|I_B1|MID  2e-12
I_PG1_01|_PG|I_B1|B 0 _PG1_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q3|B _PG1_01|_PG|Q3 _PG1_01|_PG|I_Q3|MID  2e-12
I_PG1_01|_PG|I_Q3|B 0 _PG1_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_PG|I_Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|I_Q2|MID  2e-12
I_PG1_01|_PG|I_Q2|B 0 _PG1_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|I_Q1|MID  2e-12
I_PG1_01|_PG|I_Q1|B 0 _PG1_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_PG|A1|1 _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A1|P _PG1_01|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01|_PG|A1|B _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A1|RB _PG1_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A2|1 _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A2|P _PG1_01|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01|_PG|A2|B _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A2|RB _PG1_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A12|1 _PG1_01|_PG|A2 _PG1_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|A12|B _PG1_01|_PG|A2 _PG1_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|A12|RB _PG1_01|_PG|A12|MID_SHUNT _PG1_01|_PG|A3  2.1704737578552e-12
B_PG1_01|_PG|B1|1 _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B1|P _PG1_01|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01|_PG|B1|B _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B1|RB _PG1_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B2|1 _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B2|P _PG1_01|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01|_PG|B2|B _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B2|RB _PG1_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B12|1 _PG1_01|_PG|B2 _PG1_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|B12|B _PG1_01|_PG|B2 _PG1_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|B12|RB _PG1_01|_PG|B12|MID_SHUNT _PG1_01|_PG|B3  2.1704737578552e-12
B_PG1_01|_PG|Q2|1 _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q2|P _PG1_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q2|RB _PG1_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|Q1|1 _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q1|P _PG1_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q1|RB _PG1_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_GG|I_A1|B _PG1_01|_GG|A1 _PG1_01|_GG|I_A1|MID  2e-12
I_PG1_01|_GG|I_A1|B 0 _PG1_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_B1|B _PG1_01|_GG|B1 _PG1_01|_GG|I_B1|MID  2e-12
I_PG1_01|_GG|I_B1|B 0 _PG1_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q3|B _PG1_01|_GG|Q3 _PG1_01|_GG|I_Q3|MID  2e-12
I_PG1_01|_GG|I_Q3|B 0 _PG1_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_GG|I_Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|I_Q2|MID  2e-12
I_PG1_01|_GG|I_Q2|B 0 _PG1_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|I_Q1|MID  2e-12
I_PG1_01|_GG|I_Q1|B 0 _PG1_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_GG|A1|1 _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A1|P _PG1_01|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01|_GG|A1|B _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A1|RB _PG1_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A2|1 _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A2|P _PG1_01|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01|_GG|A2|B _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A2|RB _PG1_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A12|1 _PG1_01|_GG|A2 _PG1_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|A12|B _PG1_01|_GG|A2 _PG1_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|A12|RB _PG1_01|_GG|A12|MID_SHUNT _PG1_01|_GG|A3  2.1704737578552e-12
B_PG1_01|_GG|B1|1 _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B1|P _PG1_01|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01|_GG|B1|B _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B1|RB _PG1_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B2|1 _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B2|P _PG1_01|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01|_GG|B2|B _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B2|RB _PG1_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B12|1 _PG1_01|_GG|B2 _PG1_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|B12|B _PG1_01|_GG|B2 _PG1_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|B12|RB _PG1_01|_GG|B12|MID_SHUNT _PG1_01|_GG|B3  2.1704737578552e-12
B_PG1_01|_GG|Q2|1 _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q2|P _PG1_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q2|RB _PG1_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|Q1|1 _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q1|P _PG1_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q1|RB _PG1_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_PG|I_1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|I_1|MID  2e-12
I_PG1_01|_DFF_PG|I_1|B 0 _PG1_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|I_3|MID  2e-12
I_PG1_01|_DFF_PG|I_3|B 0 _PG1_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_PG|I_T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|I_T|MID  2e-12
I_PG1_01|_DFF_PG|I_T|B 0 _PG1_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|I_6|MID  2e-12
I_PG1_01|_DFF_PG|I_6|B 0 _PG1_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_PG|1|1 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|1|P _PG1_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|1|RB _PG1_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|23|1 _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|23|B _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|23|RB _PG1_01|_DFF_PG|23|MID_SHUNT _PG1_01|_DFF_PG|A3  2.1704737578552e-12
B_PG1_01|_DFF_PG|3|1 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|3|P _PG1_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|3|RB _PG1_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|4|1 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|4|P _PG1_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|4|B _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|4|RB _PG1_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|T|1 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|T|P _PG1_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|T|RB _PG1_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|45|1 _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|45|B _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|45|RB _PG1_01|_DFF_PG|45|MID_SHUNT _PG1_01|_DFF_PG|A4  2.1704737578552e-12
B_PG1_01|_DFF_PG|6|1 _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|6|P _PG1_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|6|RB _PG1_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_GG|I_1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|I_1|MID  2e-12
I_PG1_01|_DFF_GG|I_1|B 0 _PG1_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|I_3|MID  2e-12
I_PG1_01|_DFF_GG|I_3|B 0 _PG1_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_GG|I_T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|I_T|MID  2e-12
I_PG1_01|_DFF_GG|I_T|B 0 _PG1_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|I_6|MID  2e-12
I_PG1_01|_DFF_GG|I_6|B 0 _PG1_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_GG|1|1 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|1|P _PG1_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|1|RB _PG1_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|23|1 _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|23|B _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|23|RB _PG1_01|_DFF_GG|23|MID_SHUNT _PG1_01|_DFF_GG|A3  2.1704737578552e-12
B_PG1_01|_DFF_GG|3|1 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|3|P _PG1_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|3|RB _PG1_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|4|1 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|4|P _PG1_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|4|B _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|4|RB _PG1_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|T|1 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|T|P _PG1_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|T|RB _PG1_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|45|1 _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|45|B _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|45|RB _PG1_01|_DFF_GG|45|MID_SHUNT _PG1_01|_DFF_GG|A4  2.1704737578552e-12
B_PG1_01|_DFF_GG|6|1 _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|6|P _PG1_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|6|RB _PG1_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_G|I_A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|I_A1|MID  2e-12
I_PG1_01|_AND_G|I_A1|B 0 _PG1_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|I_B1|MID  2e-12
I_PG1_01|_AND_G|I_B1|B 0 _PG1_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q3|B _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|I_Q3|MID  2e-12
I_PG1_01|_AND_G|I_Q3|B 0 _PG1_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_G|I_Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|I_Q2|MID  2e-12
I_PG1_01|_AND_G|I_Q2|B 0 _PG1_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|I_Q1|MID  2e-12
I_PG1_01|_AND_G|I_Q1|B 0 _PG1_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_G|A1|1 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A1|P _PG1_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A1|RB _PG1_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A2|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A2|P _PG1_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A2|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A2|RB _PG1_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A12|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|A12|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|A12|RB _PG1_01|_AND_G|A12|MID_SHUNT _PG1_01|_AND_G|A3  2.1704737578552e-12
B_PG1_01|_AND_G|B1|1 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B1|P _PG1_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B1|RB _PG1_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B2|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B2|P _PG1_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B2|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B2|RB _PG1_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B12|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|B12|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|B12|RB _PG1_01|_AND_G|B12|MID_SHUNT _PG1_01|_AND_G|B3  2.1704737578552e-12
B_PG1_01|_AND_G|Q2|1 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q2|P _PG1_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q2|RB _PG1_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|Q1|1 _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q1|P _PG1_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q1|RB _PG1_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|P|I_1|B _PG2_01|P|A1 _PG2_01|P|I_1|MID  2e-12
I_PG2_01|P|I_1|B 0 _PG2_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_3|B _PG2_01|P|A3 _PG2_01|P|I_3|MID  2e-12
I_PG2_01|P|I_3|B 0 _PG2_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|P|I_T|B _PG2_01|P|T1 _PG2_01|P|I_T|MID  2e-12
I_PG2_01|P|I_T|B 0 _PG2_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_6|B _PG2_01|P|Q1 _PG2_01|P|I_6|MID  2e-12
I_PG2_01|P|I_6|B 0 _PG2_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|P|1|1 _PG2_01|P|A1 _PG2_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|1|P _PG2_01|P|1|MID_SERIES 0  2e-13
R_PG2_01|P|1|B _PG2_01|P|A1 _PG2_01|P|1|MID_SHUNT  2.7439617672
L_PG2_01|P|1|RB _PG2_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|23|1 _PG2_01|P|A2 _PG2_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|P|23|B _PG2_01|P|A2 _PG2_01|P|23|MID_SHUNT  3.84154647408
L_PG2_01|P|23|RB _PG2_01|P|23|MID_SHUNT _PG2_01|P|A3  2.1704737578552e-12
B_PG2_01|P|3|1 _PG2_01|P|A3 _PG2_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|3|P _PG2_01|P|3|MID_SERIES 0  2e-13
R_PG2_01|P|3|B _PG2_01|P|A3 _PG2_01|P|3|MID_SHUNT  2.7439617672
L_PG2_01|P|3|RB _PG2_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|4|1 _PG2_01|P|A4 _PG2_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|4|P _PG2_01|P|4|MID_SERIES 0  2e-13
R_PG2_01|P|4|B _PG2_01|P|A4 _PG2_01|P|4|MID_SHUNT  2.7439617672
L_PG2_01|P|4|RB _PG2_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|T|1 _PG2_01|P|T1 _PG2_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|T|P _PG2_01|P|T|MID_SERIES 0  2e-13
R_PG2_01|P|T|B _PG2_01|P|T1 _PG2_01|P|T|MID_SHUNT  2.7439617672
L_PG2_01|P|T|RB _PG2_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|45|1 _PG2_01|P|T2 _PG2_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|P|45|B _PG2_01|P|T2 _PG2_01|P|45|MID_SHUNT  3.84154647408
L_PG2_01|P|45|RB _PG2_01|P|45|MID_SHUNT _PG2_01|P|A4  2.1704737578552e-12
B_PG2_01|P|6|1 _PG2_01|P|Q1 _PG2_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|6|P _PG2_01|P|6|MID_SERIES 0  2e-13
R_PG2_01|P|6|B _PG2_01|P|Q1 _PG2_01|P|6|MID_SHUNT  2.7439617672
L_PG2_01|P|6|RB _PG2_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|G|I_1|B _PG2_01|G|A1 _PG2_01|G|I_1|MID  2e-12
I_PG2_01|G|I_1|B 0 _PG2_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_3|B _PG2_01|G|A3 _PG2_01|G|I_3|MID  2e-12
I_PG2_01|G|I_3|B 0 _PG2_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|G|I_T|B _PG2_01|G|T1 _PG2_01|G|I_T|MID  2e-12
I_PG2_01|G|I_T|B 0 _PG2_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_6|B _PG2_01|G|Q1 _PG2_01|G|I_6|MID  2e-12
I_PG2_01|G|I_6|B 0 _PG2_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|G|1|1 _PG2_01|G|A1 _PG2_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|1|P _PG2_01|G|1|MID_SERIES 0  2e-13
R_PG2_01|G|1|B _PG2_01|G|A1 _PG2_01|G|1|MID_SHUNT  2.7439617672
L_PG2_01|G|1|RB _PG2_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|23|1 _PG2_01|G|A2 _PG2_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|G|23|B _PG2_01|G|A2 _PG2_01|G|23|MID_SHUNT  3.84154647408
L_PG2_01|G|23|RB _PG2_01|G|23|MID_SHUNT _PG2_01|G|A3  2.1704737578552e-12
B_PG2_01|G|3|1 _PG2_01|G|A3 _PG2_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|3|P _PG2_01|G|3|MID_SERIES 0  2e-13
R_PG2_01|G|3|B _PG2_01|G|A3 _PG2_01|G|3|MID_SHUNT  2.7439617672
L_PG2_01|G|3|RB _PG2_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|4|1 _PG2_01|G|A4 _PG2_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|4|P _PG2_01|G|4|MID_SERIES 0  2e-13
R_PG2_01|G|4|B _PG2_01|G|A4 _PG2_01|G|4|MID_SHUNT  2.7439617672
L_PG2_01|G|4|RB _PG2_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|T|1 _PG2_01|G|T1 _PG2_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|T|P _PG2_01|G|T|MID_SERIES 0  2e-13
R_PG2_01|G|T|B _PG2_01|G|T1 _PG2_01|G|T|MID_SHUNT  2.7439617672
L_PG2_01|G|T|RB _PG2_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|45|1 _PG2_01|G|T2 _PG2_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|G|45|B _PG2_01|G|T2 _PG2_01|G|45|MID_SHUNT  3.84154647408
L_PG2_01|G|45|RB _PG2_01|G|45|MID_SHUNT _PG2_01|G|A4  2.1704737578552e-12
B_PG2_01|G|6|1 _PG2_01|G|Q1 _PG2_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|6|P _PG2_01|G|6|MID_SERIES 0  2e-13
R_PG2_01|G|6|B _PG2_01|G|Q1 _PG2_01|G|6|MID_SHUNT  2.7439617672
L_PG2_01|G|6|RB _PG2_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_G1|I_D1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|I_D1|MID  2e-12
I_PG3_01|_SPL_G1|I_D1|B 0 _PG3_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_D2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|I_D2|MID  2e-12
I_PG3_01|_SPL_G1|I_D2|B 0 _PG3_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_G1|I_Q1|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|I_Q1|MID  2e-12
I_PG3_01|_SPL_G1|I_Q1|B 0 _PG3_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_Q2|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|I_Q2|MID  2e-12
I_PG3_01|_SPL_G1|I_Q2|B 0 _PG3_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_G1|1|1 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|1|P _PG3_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|1|RB _PG3_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|2|1 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|2|P _PG3_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|2|RB _PG3_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|A|1 _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|A|P _PG3_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|A|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|A|RB _PG3_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|B|1 _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|B|P _PG3_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|B|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|B|RB _PG3_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_P1|I_D1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|I_D1|MID  2e-12
I_PG3_01|_SPL_P1|I_D1|B 0 _PG3_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_D2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|I_D2|MID  2e-12
I_PG3_01|_SPL_P1|I_D2|B 0 _PG3_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_P1|I_Q1|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|I_Q1|MID  2e-12
I_PG3_01|_SPL_P1|I_Q1|B 0 _PG3_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_Q2|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|I_Q2|MID  2e-12
I_PG3_01|_SPL_P1|I_Q2|B 0 _PG3_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_P1|1|1 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|1|P _PG3_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|1|RB _PG3_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|2|1 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|2|P _PG3_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|2|RB _PG3_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|A|1 _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|A|P _PG3_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|A|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|A|RB _PG3_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|B|1 _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|B|P _PG3_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|B|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|B|RB _PG3_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_PG|I_A1|B _PG3_01|_PG|A1 _PG3_01|_PG|I_A1|MID  2e-12
I_PG3_01|_PG|I_A1|B 0 _PG3_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_B1|B _PG3_01|_PG|B1 _PG3_01|_PG|I_B1|MID  2e-12
I_PG3_01|_PG|I_B1|B 0 _PG3_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q3|B _PG3_01|_PG|Q3 _PG3_01|_PG|I_Q3|MID  2e-12
I_PG3_01|_PG|I_Q3|B 0 _PG3_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_PG|I_Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|I_Q2|MID  2e-12
I_PG3_01|_PG|I_Q2|B 0 _PG3_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|I_Q1|MID  2e-12
I_PG3_01|_PG|I_Q1|B 0 _PG3_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_PG|A1|1 _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A1|P _PG3_01|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01|_PG|A1|B _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A1|RB _PG3_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A2|1 _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A2|P _PG3_01|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01|_PG|A2|B _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A2|RB _PG3_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A12|1 _PG3_01|_PG|A2 _PG3_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|A12|B _PG3_01|_PG|A2 _PG3_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|A12|RB _PG3_01|_PG|A12|MID_SHUNT _PG3_01|_PG|A3  2.1704737578552e-12
B_PG3_01|_PG|B1|1 _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B1|P _PG3_01|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01|_PG|B1|B _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B1|RB _PG3_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B2|1 _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B2|P _PG3_01|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01|_PG|B2|B _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B2|RB _PG3_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B12|1 _PG3_01|_PG|B2 _PG3_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|B12|B _PG3_01|_PG|B2 _PG3_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|B12|RB _PG3_01|_PG|B12|MID_SHUNT _PG3_01|_PG|B3  2.1704737578552e-12
B_PG3_01|_PG|Q2|1 _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q2|P _PG3_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q2|RB _PG3_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|Q1|1 _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q1|P _PG3_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q1|RB _PG3_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_GG|I_A1|B _PG3_01|_GG|A1 _PG3_01|_GG|I_A1|MID  2e-12
I_PG3_01|_GG|I_A1|B 0 _PG3_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_B1|B _PG3_01|_GG|B1 _PG3_01|_GG|I_B1|MID  2e-12
I_PG3_01|_GG|I_B1|B 0 _PG3_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q3|B _PG3_01|_GG|Q3 _PG3_01|_GG|I_Q3|MID  2e-12
I_PG3_01|_GG|I_Q3|B 0 _PG3_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_GG|I_Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|I_Q2|MID  2e-12
I_PG3_01|_GG|I_Q2|B 0 _PG3_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|I_Q1|MID  2e-12
I_PG3_01|_GG|I_Q1|B 0 _PG3_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_GG|A1|1 _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A1|P _PG3_01|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01|_GG|A1|B _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A1|RB _PG3_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A2|1 _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A2|P _PG3_01|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01|_GG|A2|B _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A2|RB _PG3_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A12|1 _PG3_01|_GG|A2 _PG3_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|A12|B _PG3_01|_GG|A2 _PG3_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|A12|RB _PG3_01|_GG|A12|MID_SHUNT _PG3_01|_GG|A3  2.1704737578552e-12
B_PG3_01|_GG|B1|1 _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B1|P _PG3_01|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01|_GG|B1|B _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B1|RB _PG3_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B2|1 _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B2|P _PG3_01|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01|_GG|B2|B _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B2|RB _PG3_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B12|1 _PG3_01|_GG|B2 _PG3_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|B12|B _PG3_01|_GG|B2 _PG3_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|B12|RB _PG3_01|_GG|B12|MID_SHUNT _PG3_01|_GG|B3  2.1704737578552e-12
B_PG3_01|_GG|Q2|1 _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q2|P _PG3_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q2|RB _PG3_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|Q1|1 _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q1|P _PG3_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q1|RB _PG3_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P0|I_1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|I_1|MID  2e-12
I_PG3_01|_DFF_P0|I_1|B 0 _PG3_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|I_3|MID  2e-12
I_PG3_01|_DFF_P0|I_3|B 0 _PG3_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P0|I_T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|I_T|MID  2e-12
I_PG3_01|_DFF_P0|I_T|B 0 _PG3_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|I_6|MID  2e-12
I_PG3_01|_DFF_P0|I_6|B 0 _PG3_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P0|1|1 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|1|P _PG3_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|1|RB _PG3_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|23|1 _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|23|B _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|23|RB _PG3_01|_DFF_P0|23|MID_SHUNT _PG3_01|_DFF_P0|A3  2.1704737578552e-12
B_PG3_01|_DFF_P0|3|1 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|3|P _PG3_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|3|RB _PG3_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|4|1 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|4|P _PG3_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|4|B _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|4|RB _PG3_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|T|1 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|T|P _PG3_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|T|RB _PG3_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|45|1 _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|45|B _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|45|RB _PG3_01|_DFF_P0|45|MID_SHUNT _PG3_01|_DFF_P0|A4  2.1704737578552e-12
B_PG3_01|_DFF_P0|6|1 _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|6|P _PG3_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|6|RB _PG3_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P1|I_1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|I_1|MID  2e-12
I_PG3_01|_DFF_P1|I_1|B 0 _PG3_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|I_3|MID  2e-12
I_PG3_01|_DFF_P1|I_3|B 0 _PG3_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P1|I_T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|I_T|MID  2e-12
I_PG3_01|_DFF_P1|I_T|B 0 _PG3_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|I_6|MID  2e-12
I_PG3_01|_DFF_P1|I_6|B 0 _PG3_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P1|1|1 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|1|P _PG3_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|1|RB _PG3_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|23|1 _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|23|B _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|23|RB _PG3_01|_DFF_P1|23|MID_SHUNT _PG3_01|_DFF_P1|A3  2.1704737578552e-12
B_PG3_01|_DFF_P1|3|1 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|3|P _PG3_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|3|RB _PG3_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|4|1 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|4|P _PG3_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|4|B _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|4|RB _PG3_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|T|1 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|T|P _PG3_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|T|RB _PG3_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|45|1 _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|45|B _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|45|RB _PG3_01|_DFF_P1|45|MID_SHUNT _PG3_01|_DFF_P1|A4  2.1704737578552e-12
B_PG3_01|_DFF_P1|6|1 _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|6|P _PG3_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|6|RB _PG3_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_PG|I_1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|I_1|MID  2e-12
I_PG3_01|_DFF_PG|I_1|B 0 _PG3_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|I_3|MID  2e-12
I_PG3_01|_DFF_PG|I_3|B 0 _PG3_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_PG|I_T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|I_T|MID  2e-12
I_PG3_01|_DFF_PG|I_T|B 0 _PG3_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|I_6|MID  2e-12
I_PG3_01|_DFF_PG|I_6|B 0 _PG3_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_PG|1|1 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|1|P _PG3_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|1|RB _PG3_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|23|1 _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|23|B _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|23|RB _PG3_01|_DFF_PG|23|MID_SHUNT _PG3_01|_DFF_PG|A3  2.1704737578552e-12
B_PG3_01|_DFF_PG|3|1 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|3|P _PG3_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|3|RB _PG3_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|4|1 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|4|P _PG3_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|4|B _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|4|RB _PG3_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|T|1 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|T|P _PG3_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|T|RB _PG3_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|45|1 _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|45|B _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|45|RB _PG3_01|_DFF_PG|45|MID_SHUNT _PG3_01|_DFF_PG|A4  2.1704737578552e-12
B_PG3_01|_DFF_PG|6|1 _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|6|P _PG3_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|6|RB _PG3_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_GG|I_1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|I_1|MID  2e-12
I_PG3_01|_DFF_GG|I_1|B 0 _PG3_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|I_3|MID  2e-12
I_PG3_01|_DFF_GG|I_3|B 0 _PG3_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_GG|I_T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|I_T|MID  2e-12
I_PG3_01|_DFF_GG|I_T|B 0 _PG3_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|I_6|MID  2e-12
I_PG3_01|_DFF_GG|I_6|B 0 _PG3_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_GG|1|1 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|1|P _PG3_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|1|RB _PG3_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|23|1 _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|23|B _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|23|RB _PG3_01|_DFF_GG|23|MID_SHUNT _PG3_01|_DFF_GG|A3  2.1704737578552e-12
B_PG3_01|_DFF_GG|3|1 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|3|P _PG3_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|3|RB _PG3_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|4|1 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|4|P _PG3_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|4|B _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|4|RB _PG3_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|T|1 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|T|P _PG3_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|T|RB _PG3_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|45|1 _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|45|B _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|45|RB _PG3_01|_DFF_GG|45|MID_SHUNT _PG3_01|_DFF_GG|A4  2.1704737578552e-12
B_PG3_01|_DFF_GG|6|1 _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|6|P _PG3_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|6|RB _PG3_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_G|I_A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|I_A1|MID  2e-12
I_PG3_01|_AND_G|I_A1|B 0 _PG3_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|I_B1|MID  2e-12
I_PG3_01|_AND_G|I_B1|B 0 _PG3_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q3|B _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|I_Q3|MID  2e-12
I_PG3_01|_AND_G|I_Q3|B 0 _PG3_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_G|I_Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|I_Q2|MID  2e-12
I_PG3_01|_AND_G|I_Q2|B 0 _PG3_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|I_Q1|MID  2e-12
I_PG3_01|_AND_G|I_Q1|B 0 _PG3_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_G|A1|1 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A1|P _PG3_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A1|RB _PG3_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A2|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A2|P _PG3_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A2|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A2|RB _PG3_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A12|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|A12|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|A12|RB _PG3_01|_AND_G|A12|MID_SHUNT _PG3_01|_AND_G|A3  2.1704737578552e-12
B_PG3_01|_AND_G|B1|1 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B1|P _PG3_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B1|RB _PG3_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B2|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B2|P _PG3_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B2|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B2|RB _PG3_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B12|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|B12|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|B12|RB _PG3_01|_AND_G|B12|MID_SHUNT _PG3_01|_AND_G|B3  2.1704737578552e-12
B_PG3_01|_AND_G|Q2|1 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q2|P _PG3_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q2|RB _PG3_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|Q1|1 _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q1|P _PG3_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q1|RB _PG3_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_P|I_A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|I_A1|MID  2e-12
I_PG3_01|_AND_P|I_A1|B 0 _PG3_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|I_B1|MID  2e-12
I_PG3_01|_AND_P|I_B1|B 0 _PG3_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q3|B _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|I_Q3|MID  2e-12
I_PG3_01|_AND_P|I_Q3|B 0 _PG3_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_P|I_Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|I_Q2|MID  2e-12
I_PG3_01|_AND_P|I_Q2|B 0 _PG3_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|I_Q1|MID  2e-12
I_PG3_01|_AND_P|I_Q1|B 0 _PG3_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_P|A1|1 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A1|P _PG3_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A1|RB _PG3_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A2|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A2|P _PG3_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A2|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A2|RB _PG3_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A12|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|A12|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|A12|RB _PG3_01|_AND_P|A12|MID_SHUNT _PG3_01|_AND_P|A3  2.1704737578552e-12
B_PG3_01|_AND_P|B1|1 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B1|P _PG3_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B1|RB _PG3_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B2|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B2|P _PG3_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B2|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B2|RB _PG3_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B12|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|B12|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|B12|RB _PG3_01|_AND_P|B12|MID_SHUNT _PG3_01|_AND_P|B3  2.1704737578552e-12
B_PG3_01|_AND_P|Q2|1 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q2|P _PG3_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q2|RB _PG3_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|Q1|1 _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q1|P _PG3_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q1|RB _PG3_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL1|I_D1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|I_D1|MID  2e-12
ISPL_G1_1|SPL1|I_D1|B 0 SPL_G1_1|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_D2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|I_D2|MID  2e-12
ISPL_G1_1|SPL1|I_D2|B 0 SPL_G1_1|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL1|I_Q1|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|I_Q1|MID  2e-12
ISPL_G1_1|SPL1|I_Q1|B 0 SPL_G1_1|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_Q2|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|I_Q2|MID  2e-12
ISPL_G1_1|SPL1|I_Q2|B 0 SPL_G1_1|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL1|1|1 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|1|P SPL_G1_1|SPL1|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|1|RB SPL_G1_1|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|2|1 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|2|P SPL_G1_1|SPL1|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|2|RB SPL_G1_1|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|A|1 SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|A|P SPL_G1_1|SPL1|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|A|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|A|RB SPL_G1_1|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|B|1 SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|B|P SPL_G1_1|SPL1|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|B|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|B|RB SPL_G1_1|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL2|I_D1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|I_D1|MID  2e-12
ISPL_G1_1|SPL2|I_D1|B 0 SPL_G1_1|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_D2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|I_D2|MID  2e-12
ISPL_G1_1|SPL2|I_D2|B 0 SPL_G1_1|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL2|I_Q1|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|I_Q1|MID  2e-12
ISPL_G1_1|SPL2|I_Q1|B 0 SPL_G1_1|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_Q2|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|I_Q2|MID  2e-12
ISPL_G1_1|SPL2|I_Q2|B 0 SPL_G1_1|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL2|1|1 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|1|P SPL_G1_1|SPL2|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|1|RB SPL_G1_1|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|2|1 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|2|P SPL_G1_1|SPL2|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|2|RB SPL_G1_1|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|A|1 SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|A|P SPL_G1_1|SPL2|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|A|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|A|RB SPL_G1_1|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|B|1 SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|B|P SPL_G1_1|SPL2|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|B|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|B|RB SPL_G1_1|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|P|I_1|B _PG0_12|P|A1 _PG0_12|P|I_1|MID  2e-12
I_PG0_12|P|I_1|B 0 _PG0_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_3|B _PG0_12|P|A3 _PG0_12|P|I_3|MID  2e-12
I_PG0_12|P|I_3|B 0 _PG0_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|P|I_T|B _PG0_12|P|T1 _PG0_12|P|I_T|MID  2e-12
I_PG0_12|P|I_T|B 0 _PG0_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_6|B _PG0_12|P|Q1 _PG0_12|P|I_6|MID  2e-12
I_PG0_12|P|I_6|B 0 _PG0_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|P|1|1 _PG0_12|P|A1 _PG0_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|1|P _PG0_12|P|1|MID_SERIES 0  2e-13
R_PG0_12|P|1|B _PG0_12|P|A1 _PG0_12|P|1|MID_SHUNT  2.7439617672
L_PG0_12|P|1|RB _PG0_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|23|1 _PG0_12|P|A2 _PG0_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|P|23|B _PG0_12|P|A2 _PG0_12|P|23|MID_SHUNT  3.84154647408
L_PG0_12|P|23|RB _PG0_12|P|23|MID_SHUNT _PG0_12|P|A3  2.1704737578552e-12
B_PG0_12|P|3|1 _PG0_12|P|A3 _PG0_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|3|P _PG0_12|P|3|MID_SERIES 0  2e-13
R_PG0_12|P|3|B _PG0_12|P|A3 _PG0_12|P|3|MID_SHUNT  2.7439617672
L_PG0_12|P|3|RB _PG0_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|4|1 _PG0_12|P|A4 _PG0_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|4|P _PG0_12|P|4|MID_SERIES 0  2e-13
R_PG0_12|P|4|B _PG0_12|P|A4 _PG0_12|P|4|MID_SHUNT  2.7439617672
L_PG0_12|P|4|RB _PG0_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|T|1 _PG0_12|P|T1 _PG0_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|T|P _PG0_12|P|T|MID_SERIES 0  2e-13
R_PG0_12|P|T|B _PG0_12|P|T1 _PG0_12|P|T|MID_SHUNT  2.7439617672
L_PG0_12|P|T|RB _PG0_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|45|1 _PG0_12|P|T2 _PG0_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|P|45|B _PG0_12|P|T2 _PG0_12|P|45|MID_SHUNT  3.84154647408
L_PG0_12|P|45|RB _PG0_12|P|45|MID_SHUNT _PG0_12|P|A4  2.1704737578552e-12
B_PG0_12|P|6|1 _PG0_12|P|Q1 _PG0_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|6|P _PG0_12|P|6|MID_SERIES 0  2e-13
R_PG0_12|P|6|B _PG0_12|P|Q1 _PG0_12|P|6|MID_SHUNT  2.7439617672
L_PG0_12|P|6|RB _PG0_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|G|I_1|B _PG0_12|G|A1 _PG0_12|G|I_1|MID  2e-12
I_PG0_12|G|I_1|B 0 _PG0_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_3|B _PG0_12|G|A3 _PG0_12|G|I_3|MID  2e-12
I_PG0_12|G|I_3|B 0 _PG0_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|G|I_T|B _PG0_12|G|T1 _PG0_12|G|I_T|MID  2e-12
I_PG0_12|G|I_T|B 0 _PG0_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_6|B _PG0_12|G|Q1 _PG0_12|G|I_6|MID  2e-12
I_PG0_12|G|I_6|B 0 _PG0_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|G|1|1 _PG0_12|G|A1 _PG0_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|1|P _PG0_12|G|1|MID_SERIES 0  2e-13
R_PG0_12|G|1|B _PG0_12|G|A1 _PG0_12|G|1|MID_SHUNT  2.7439617672
L_PG0_12|G|1|RB _PG0_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|23|1 _PG0_12|G|A2 _PG0_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|G|23|B _PG0_12|G|A2 _PG0_12|G|23|MID_SHUNT  3.84154647408
L_PG0_12|G|23|RB _PG0_12|G|23|MID_SHUNT _PG0_12|G|A3  2.1704737578552e-12
B_PG0_12|G|3|1 _PG0_12|G|A3 _PG0_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|3|P _PG0_12|G|3|MID_SERIES 0  2e-13
R_PG0_12|G|3|B _PG0_12|G|A3 _PG0_12|G|3|MID_SHUNT  2.7439617672
L_PG0_12|G|3|RB _PG0_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|4|1 _PG0_12|G|A4 _PG0_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|4|P _PG0_12|G|4|MID_SERIES 0  2e-13
R_PG0_12|G|4|B _PG0_12|G|A4 _PG0_12|G|4|MID_SHUNT  2.7439617672
L_PG0_12|G|4|RB _PG0_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|T|1 _PG0_12|G|T1 _PG0_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|T|P _PG0_12|G|T|MID_SERIES 0  2e-13
R_PG0_12|G|T|B _PG0_12|G|T1 _PG0_12|G|T|MID_SHUNT  2.7439617672
L_PG0_12|G|T|RB _PG0_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|45|1 _PG0_12|G|T2 _PG0_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|G|45|B _PG0_12|G|T2 _PG0_12|G|45|MID_SHUNT  3.84154647408
L_PG0_12|G|45|RB _PG0_12|G|45|MID_SHUNT _PG0_12|G|A4  2.1704737578552e-12
B_PG0_12|G|6|1 _PG0_12|G|Q1 _PG0_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|6|P _PG0_12|G|6|MID_SERIES 0  2e-13
R_PG0_12|G|6|B _PG0_12|G|Q1 _PG0_12|G|6|MID_SHUNT  2.7439617672
L_PG0_12|G|6|RB _PG0_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|I_D1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|I_D1|MID  2e-12
I_PG2_12|_SPL_G1|I_D1|B 0 _PG2_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_D2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|I_D2|MID  2e-12
I_PG2_12|_SPL_G1|I_D2|B 0 _PG2_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG2_12|_SPL_G1|I_Q1|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|I_Q1|MID  2e-12
I_PG2_12|_SPL_G1|I_Q1|B 0 _PG2_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_Q2|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|I_Q2|MID  2e-12
I_PG2_12|_SPL_G1|I_Q2|B 0 _PG2_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG2_12|_SPL_G1|1|1 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|1|P _PG2_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|1|RB _PG2_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|2|1 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|2|P _PG2_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|2|RB _PG2_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|A|1 _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|A|P _PG2_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|A|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|A|RB _PG2_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|B|1 _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|B|P _PG2_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|B|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|B|RB _PG2_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_PG|I_A1|B _PG2_12|_PG|A1 _PG2_12|_PG|I_A1|MID  2e-12
I_PG2_12|_PG|I_A1|B 0 _PG2_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_B1|B _PG2_12|_PG|B1 _PG2_12|_PG|I_B1|MID  2e-12
I_PG2_12|_PG|I_B1|B 0 _PG2_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q3|B _PG2_12|_PG|Q3 _PG2_12|_PG|I_Q3|MID  2e-12
I_PG2_12|_PG|I_Q3|B 0 _PG2_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_PG|I_Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|I_Q2|MID  2e-12
I_PG2_12|_PG|I_Q2|B 0 _PG2_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|I_Q1|MID  2e-12
I_PG2_12|_PG|I_Q1|B 0 _PG2_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_PG|A1|1 _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A1|P _PG2_12|_PG|A1|MID_SERIES 0  2e-13
R_PG2_12|_PG|A1|B _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A1|RB _PG2_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A2|1 _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A2|P _PG2_12|_PG|A2|MID_SERIES 0  2e-13
R_PG2_12|_PG|A2|B _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A2|RB _PG2_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A12|1 _PG2_12|_PG|A2 _PG2_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|A12|B _PG2_12|_PG|A2 _PG2_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|A12|RB _PG2_12|_PG|A12|MID_SHUNT _PG2_12|_PG|A3  2.1704737578552e-12
B_PG2_12|_PG|B1|1 _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B1|P _PG2_12|_PG|B1|MID_SERIES 0  2e-13
R_PG2_12|_PG|B1|B _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B1|RB _PG2_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B2|1 _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B2|P _PG2_12|_PG|B2|MID_SERIES 0  2e-13
R_PG2_12|_PG|B2|B _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B2|RB _PG2_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B12|1 _PG2_12|_PG|B2 _PG2_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|B12|B _PG2_12|_PG|B2 _PG2_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|B12|RB _PG2_12|_PG|B12|MID_SHUNT _PG2_12|_PG|B3  2.1704737578552e-12
B_PG2_12|_PG|Q2|1 _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q2|P _PG2_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q2|RB _PG2_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|Q1|1 _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q1|P _PG2_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q1|RB _PG2_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_GG|I_A1|B _PG2_12|_GG|A1 _PG2_12|_GG|I_A1|MID  2e-12
I_PG2_12|_GG|I_A1|B 0 _PG2_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_B1|B _PG2_12|_GG|B1 _PG2_12|_GG|I_B1|MID  2e-12
I_PG2_12|_GG|I_B1|B 0 _PG2_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q3|B _PG2_12|_GG|Q3 _PG2_12|_GG|I_Q3|MID  2e-12
I_PG2_12|_GG|I_Q3|B 0 _PG2_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_GG|I_Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|I_Q2|MID  2e-12
I_PG2_12|_GG|I_Q2|B 0 _PG2_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|I_Q1|MID  2e-12
I_PG2_12|_GG|I_Q1|B 0 _PG2_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_GG|A1|1 _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A1|P _PG2_12|_GG|A1|MID_SERIES 0  2e-13
R_PG2_12|_GG|A1|B _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A1|RB _PG2_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A2|1 _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A2|P _PG2_12|_GG|A2|MID_SERIES 0  2e-13
R_PG2_12|_GG|A2|B _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A2|RB _PG2_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A12|1 _PG2_12|_GG|A2 _PG2_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|A12|B _PG2_12|_GG|A2 _PG2_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|A12|RB _PG2_12|_GG|A12|MID_SHUNT _PG2_12|_GG|A3  2.1704737578552e-12
B_PG2_12|_GG|B1|1 _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B1|P _PG2_12|_GG|B1|MID_SERIES 0  2e-13
R_PG2_12|_GG|B1|B _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B1|RB _PG2_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B2|1 _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B2|P _PG2_12|_GG|B2|MID_SERIES 0  2e-13
R_PG2_12|_GG|B2|B _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B2|RB _PG2_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B12|1 _PG2_12|_GG|B2 _PG2_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|B12|B _PG2_12|_GG|B2 _PG2_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|B12|RB _PG2_12|_GG|B12|MID_SHUNT _PG2_12|_GG|B3  2.1704737578552e-12
B_PG2_12|_GG|Q2|1 _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q2|P _PG2_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q2|RB _PG2_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|Q1|1 _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q1|P _PG2_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q1|RB _PG2_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_PG|I_1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|I_1|MID  2e-12
I_PG2_12|_DFF_PG|I_1|B 0 _PG2_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|I_3|MID  2e-12
I_PG2_12|_DFF_PG|I_3|B 0 _PG2_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_PG|I_T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|I_T|MID  2e-12
I_PG2_12|_DFF_PG|I_T|B 0 _PG2_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|I_6|MID  2e-12
I_PG2_12|_DFF_PG|I_6|B 0 _PG2_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_PG|1|1 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|1|P _PG2_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|1|RB _PG2_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|23|1 _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|23|B _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|23|RB _PG2_12|_DFF_PG|23|MID_SHUNT _PG2_12|_DFF_PG|A3  2.1704737578552e-12
B_PG2_12|_DFF_PG|3|1 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|3|P _PG2_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|3|RB _PG2_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|4|1 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|4|P _PG2_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|4|B _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|4|RB _PG2_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|T|1 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|T|P _PG2_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|T|RB _PG2_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|45|1 _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|45|B _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|45|RB _PG2_12|_DFF_PG|45|MID_SHUNT _PG2_12|_DFF_PG|A4  2.1704737578552e-12
B_PG2_12|_DFF_PG|6|1 _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|6|P _PG2_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|6|RB _PG2_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_GG|I_1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|I_1|MID  2e-12
I_PG2_12|_DFF_GG|I_1|B 0 _PG2_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|I_3|MID  2e-12
I_PG2_12|_DFF_GG|I_3|B 0 _PG2_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_GG|I_T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|I_T|MID  2e-12
I_PG2_12|_DFF_GG|I_T|B 0 _PG2_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|I_6|MID  2e-12
I_PG2_12|_DFF_GG|I_6|B 0 _PG2_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_GG|1|1 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|1|P _PG2_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|1|RB _PG2_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|23|1 _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|23|B _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|23|RB _PG2_12|_DFF_GG|23|MID_SHUNT _PG2_12|_DFF_GG|A3  2.1704737578552e-12
B_PG2_12|_DFF_GG|3|1 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|3|P _PG2_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|3|RB _PG2_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|4|1 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|4|P _PG2_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|4|B _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|4|RB _PG2_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|T|1 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|T|P _PG2_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|T|RB _PG2_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|45|1 _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|45|B _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|45|RB _PG2_12|_DFF_GG|45|MID_SHUNT _PG2_12|_DFF_GG|A4  2.1704737578552e-12
B_PG2_12|_DFF_GG|6|1 _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|6|P _PG2_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|6|RB _PG2_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_G|I_A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|I_A1|MID  2e-12
I_PG2_12|_AND_G|I_A1|B 0 _PG2_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|I_B1|MID  2e-12
I_PG2_12|_AND_G|I_B1|B 0 _PG2_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q3|B _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|I_Q3|MID  2e-12
I_PG2_12|_AND_G|I_Q3|B 0 _PG2_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_G|I_Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|I_Q2|MID  2e-12
I_PG2_12|_AND_G|I_Q2|B 0 _PG2_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|I_Q1|MID  2e-12
I_PG2_12|_AND_G|I_Q1|B 0 _PG2_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_G|A1|1 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A1|P _PG2_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A1|RB _PG2_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A2|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A2|P _PG2_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A2|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A2|RB _PG2_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A12|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|A12|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|A12|RB _PG2_12|_AND_G|A12|MID_SHUNT _PG2_12|_AND_G|A3  2.1704737578552e-12
B_PG2_12|_AND_G|B1|1 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B1|P _PG2_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B1|RB _PG2_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B2|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B2|P _PG2_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B2|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B2|RB _PG2_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B12|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|B12|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|B12|RB _PG2_12|_AND_G|B12|MID_SHUNT _PG2_12|_AND_G|B3  2.1704737578552e-12
B_PG2_12|_AND_G|Q2|1 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q2|P _PG2_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q2|RB _PG2_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|Q1|1 _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q1|P _PG2_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q1|RB _PG2_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_SPL_G1|I_D1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|I_D1|MID  2e-12
I_PG3_12|_SPL_G1|I_D1|B 0 _PG3_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_D2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|I_D2|MID  2e-12
I_PG3_12|_SPL_G1|I_D2|B 0 _PG3_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_12|_SPL_G1|I_Q1|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|I_Q1|MID  2e-12
I_PG3_12|_SPL_G1|I_Q1|B 0 _PG3_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_Q2|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|I_Q2|MID  2e-12
I_PG3_12|_SPL_G1|I_Q2|B 0 _PG3_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_12|_SPL_G1|1|1 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|1|P _PG3_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|1|RB _PG3_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|2|1 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|2|P _PG3_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|2|RB _PG3_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|A|1 _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|A|P _PG3_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|A|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|A|RB _PG3_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|B|1 _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|B|P _PG3_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|B|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|B|RB _PG3_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_PG|I_A1|B _PG3_12|_PG|A1 _PG3_12|_PG|I_A1|MID  2e-12
I_PG3_12|_PG|I_A1|B 0 _PG3_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_B1|B _PG3_12|_PG|B1 _PG3_12|_PG|I_B1|MID  2e-12
I_PG3_12|_PG|I_B1|B 0 _PG3_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q3|B _PG3_12|_PG|Q3 _PG3_12|_PG|I_Q3|MID  2e-12
I_PG3_12|_PG|I_Q3|B 0 _PG3_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_PG|I_Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|I_Q2|MID  2e-12
I_PG3_12|_PG|I_Q2|B 0 _PG3_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|I_Q1|MID  2e-12
I_PG3_12|_PG|I_Q1|B 0 _PG3_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_PG|A1|1 _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A1|P _PG3_12|_PG|A1|MID_SERIES 0  2e-13
R_PG3_12|_PG|A1|B _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A1|RB _PG3_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A2|1 _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A2|P _PG3_12|_PG|A2|MID_SERIES 0  2e-13
R_PG3_12|_PG|A2|B _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A2|RB _PG3_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A12|1 _PG3_12|_PG|A2 _PG3_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|A12|B _PG3_12|_PG|A2 _PG3_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|A12|RB _PG3_12|_PG|A12|MID_SHUNT _PG3_12|_PG|A3  2.1704737578552e-12
B_PG3_12|_PG|B1|1 _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B1|P _PG3_12|_PG|B1|MID_SERIES 0  2e-13
R_PG3_12|_PG|B1|B _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B1|RB _PG3_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B2|1 _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B2|P _PG3_12|_PG|B2|MID_SERIES 0  2e-13
R_PG3_12|_PG|B2|B _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B2|RB _PG3_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B12|1 _PG3_12|_PG|B2 _PG3_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|B12|B _PG3_12|_PG|B2 _PG3_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|B12|RB _PG3_12|_PG|B12|MID_SHUNT _PG3_12|_PG|B3  2.1704737578552e-12
B_PG3_12|_PG|Q2|1 _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q2|P _PG3_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q2|RB _PG3_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|Q1|1 _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q1|P _PG3_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q1|RB _PG3_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_GG|I_A1|B _PG3_12|_GG|A1 _PG3_12|_GG|I_A1|MID  2e-12
I_PG3_12|_GG|I_A1|B 0 _PG3_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_B1|B _PG3_12|_GG|B1 _PG3_12|_GG|I_B1|MID  2e-12
I_PG3_12|_GG|I_B1|B 0 _PG3_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q3|B _PG3_12|_GG|Q3 _PG3_12|_GG|I_Q3|MID  2e-12
I_PG3_12|_GG|I_Q3|B 0 _PG3_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_GG|I_Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|I_Q2|MID  2e-12
I_PG3_12|_GG|I_Q2|B 0 _PG3_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|I_Q1|MID  2e-12
I_PG3_12|_GG|I_Q1|B 0 _PG3_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_GG|A1|1 _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A1|P _PG3_12|_GG|A1|MID_SERIES 0  2e-13
R_PG3_12|_GG|A1|B _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A1|RB _PG3_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A2|1 _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A2|P _PG3_12|_GG|A2|MID_SERIES 0  2e-13
R_PG3_12|_GG|A2|B _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A2|RB _PG3_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A12|1 _PG3_12|_GG|A2 _PG3_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|A12|B _PG3_12|_GG|A2 _PG3_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|A12|RB _PG3_12|_GG|A12|MID_SHUNT _PG3_12|_GG|A3  2.1704737578552e-12
B_PG3_12|_GG|B1|1 _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B1|P _PG3_12|_GG|B1|MID_SERIES 0  2e-13
R_PG3_12|_GG|B1|B _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B1|RB _PG3_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B2|1 _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B2|P _PG3_12|_GG|B2|MID_SERIES 0  2e-13
R_PG3_12|_GG|B2|B _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B2|RB _PG3_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B12|1 _PG3_12|_GG|B2 _PG3_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|B12|B _PG3_12|_GG|B2 _PG3_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|B12|RB _PG3_12|_GG|B12|MID_SHUNT _PG3_12|_GG|B3  2.1704737578552e-12
B_PG3_12|_GG|Q2|1 _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q2|P _PG3_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q2|RB _PG3_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|Q1|1 _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q1|P _PG3_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q1|RB _PG3_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_PG|I_1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|I_1|MID  2e-12
I_PG3_12|_DFF_PG|I_1|B 0 _PG3_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|I_3|MID  2e-12
I_PG3_12|_DFF_PG|I_3|B 0 _PG3_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_PG|I_T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|I_T|MID  2e-12
I_PG3_12|_DFF_PG|I_T|B 0 _PG3_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|I_6|MID  2e-12
I_PG3_12|_DFF_PG|I_6|B 0 _PG3_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_PG|1|1 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|1|P _PG3_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|1|RB _PG3_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|23|1 _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|23|B _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|23|RB _PG3_12|_DFF_PG|23|MID_SHUNT _PG3_12|_DFF_PG|A3  2.1704737578552e-12
B_PG3_12|_DFF_PG|3|1 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|3|P _PG3_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|3|RB _PG3_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|4|1 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|4|P _PG3_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|4|B _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|4|RB _PG3_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|T|1 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|T|P _PG3_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|T|RB _PG3_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|45|1 _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|45|B _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|45|RB _PG3_12|_DFF_PG|45|MID_SHUNT _PG3_12|_DFF_PG|A4  2.1704737578552e-12
B_PG3_12|_DFF_PG|6|1 _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|6|P _PG3_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|6|RB _PG3_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_GG|I_1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|I_1|MID  2e-12
I_PG3_12|_DFF_GG|I_1|B 0 _PG3_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|I_3|MID  2e-12
I_PG3_12|_DFF_GG|I_3|B 0 _PG3_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_GG|I_T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|I_T|MID  2e-12
I_PG3_12|_DFF_GG|I_T|B 0 _PG3_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|I_6|MID  2e-12
I_PG3_12|_DFF_GG|I_6|B 0 _PG3_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_GG|1|1 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|1|P _PG3_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|1|RB _PG3_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|23|1 _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|23|B _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|23|RB _PG3_12|_DFF_GG|23|MID_SHUNT _PG3_12|_DFF_GG|A3  2.1704737578552e-12
B_PG3_12|_DFF_GG|3|1 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|3|P _PG3_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|3|RB _PG3_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|4|1 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|4|P _PG3_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|4|B _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|4|RB _PG3_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|T|1 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|T|P _PG3_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|T|RB _PG3_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|45|1 _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|45|B _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|45|RB _PG3_12|_DFF_GG|45|MID_SHUNT _PG3_12|_DFF_GG|A4  2.1704737578552e-12
B_PG3_12|_DFF_GG|6|1 _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|6|P _PG3_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|6|RB _PG3_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_G|I_A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|I_A1|MID  2e-12
I_PG3_12|_AND_G|I_A1|B 0 _PG3_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|I_B1|MID  2e-12
I_PG3_12|_AND_G|I_B1|B 0 _PG3_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q3|B _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|I_Q3|MID  2e-12
I_PG3_12|_AND_G|I_Q3|B 0 _PG3_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_G|I_Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|I_Q2|MID  2e-12
I_PG3_12|_AND_G|I_Q2|B 0 _PG3_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|I_Q1|MID  2e-12
I_PG3_12|_AND_G|I_Q1|B 0 _PG3_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_G|A1|1 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A1|P _PG3_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A1|RB _PG3_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A2|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A2|P _PG3_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A2|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A2|RB _PG3_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A12|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|A12|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|A12|RB _PG3_12|_AND_G|A12|MID_SHUNT _PG3_12|_AND_G|A3  2.1704737578552e-12
B_PG3_12|_AND_G|B1|1 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B1|P _PG3_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B1|RB _PG3_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B2|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B2|P _PG3_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B2|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B2|RB _PG3_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B12|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|B12|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|B12|RB _PG3_12|_AND_G|B12|MID_SHUNT _PG3_12|_AND_G|B3  2.1704737578552e-12
B_PG3_12|_AND_G|Q2|1 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q2|P _PG3_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q2|RB _PG3_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|Q1|1 _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q1|P _PG3_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q1|RB _PG3_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_S0
.print DEVI R_S1
.print DEVI R_S2
.print DEVI R_S3
.print DEVI R_S4
.print DEVI I_VEC|A0
.print DEVI I_VEC|A1
.print DEVI I_VEC|A2
.print DEVI I_VEC|A3
.print DEVI I_VEC|B0
.print DEVI I_VEC|B1
.print DEVI I_VEC|B2
.print DEVI I_VEC|B3
.print DEVI IT00|T
.print DEVI IT01|T
.print DEVI IT02|T
.print DEVI IT03|T
.print DEVI LSPL_IG0_0|1
.print DEVI LSPL_IG0_0|2
.print DEVI LSPL_IG0_0|3
.print DEVI LSPL_IG0_0|4
.print DEVI LSPL_IG0_0|5
.print DEVI LSPL_IG0_0|6
.print DEVI LSPL_IG0_0|7
.print DEVI LSPL_IP1_0|1
.print DEVI LSPL_IP1_0|2
.print DEVI LSPL_IP1_0|3
.print DEVI LSPL_IP1_0|4
.print DEVI LSPL_IP1_0|5
.print DEVI LSPL_IP1_0|6
.print DEVI LSPL_IP1_0|7
.print DEVI LSPL_IG2_0|1
.print DEVI LSPL_IG2_0|2
.print DEVI LSPL_IG2_0|3
.print DEVI LSPL_IG2_0|4
.print DEVI LSPL_IG2_0|5
.print DEVI LSPL_IG2_0|6
.print DEVI LSPL_IG2_0|7
.print DEVI LSPL_IP3_0|1
.print DEVI LSPL_IP3_0|2
.print DEVI LSPL_IP3_0|3
.print DEVI LSPL_IP3_0|4
.print DEVI LSPL_IP3_0|5
.print DEVI LSPL_IP3_0|6
.print DEVI LSPL_IP3_0|7
.print DEVI IT04|T
.print DEVI IT05|T
.print DEVI IT06|T
.print DEVI IT07|T
.print DEVI ID01|T
.print DEVI L_DFF_IP1_01|1
.print DEVI L_DFF_IP1_01|2
.print DEVI L_DFF_IP1_01|3
.print DEVI L_DFF_IP1_01|T
.print DEVI L_DFF_IP1_01|4
.print DEVI L_DFF_IP1_01|5
.print DEVI L_DFF_IP1_01|6
.print DEVI ID02|T
.print DEVI L_DFF_IP2_01|1
.print DEVI L_DFF_IP2_01|2
.print DEVI L_DFF_IP2_01|3
.print DEVI L_DFF_IP2_01|T
.print DEVI L_DFF_IP2_01|4
.print DEVI L_DFF_IP2_01|5
.print DEVI L_DFF_IP2_01|6
.print DEVI ID03|T
.print DEVI L_DFF_IP3_01|1
.print DEVI L_DFF_IP3_01|2
.print DEVI L_DFF_IP3_01|3
.print DEVI L_DFF_IP3_01|T
.print DEVI L_DFF_IP3_01|4
.print DEVI L_DFF_IP3_01|5
.print DEVI L_DFF_IP3_01|6
.print DEVI IT08|T
.print DEVI IT09|T
.print DEVI L_PG1_12|1
.print DEVI L_PG1_12|2
.print DEVI L_PG1_12|3
.print DEVI L_PG1_12|T
.print DEVI L_PG1_12|4
.print DEVI L_PG1_12|5
.print DEVI L_PG1_12|6
.print DEVI IT10|T
.print DEVI IT11|T
.print DEVI ID11|T
.print DEVI L_DFF_IP1_12|1
.print DEVI L_DFF_IP1_12|2
.print DEVI L_DFF_IP1_12|3
.print DEVI L_DFF_IP1_12|T
.print DEVI L_DFF_IP1_12|4
.print DEVI L_DFF_IP1_12|5
.print DEVI L_DFF_IP1_12|6
.print DEVI ID12|T
.print DEVI L_DFF_IP2_12|1
.print DEVI L_DFF_IP2_12|2
.print DEVI L_DFF_IP2_12|3
.print DEVI L_DFF_IP2_12|T
.print DEVI L_DFF_IP2_12|4
.print DEVI L_DFF_IP2_12|5
.print DEVI L_DFF_IP2_12|6
.print DEVI ID13|T
.print DEVI L_DFF_IP3_12|1
.print DEVI L_DFF_IP3_12|2
.print DEVI L_DFF_IP3_12|3
.print DEVI L_DFF_IP3_12|T
.print DEVI L_DFF_IP3_12|4
.print DEVI L_DFF_IP3_12|5
.print DEVI L_DFF_IP3_12|6
.print DEVI IT12|T
.print DEVI L_S0|1
.print DEVI L_S0|2
.print DEVI L_S0|3
.print DEVI L_S0|T
.print DEVI L_S0|4
.print DEVI L_S0|5
.print DEVI L_S0|6
.print DEVI IT13|T
.print DEVI L_S1|A1
.print DEVI L_S1|A2
.print DEVI L_S1|A3
.print DEVI L_S1|B1
.print DEVI L_S1|B2
.print DEVI L_S1|B3
.print DEVI L_S1|T1
.print DEVI L_S1|T2
.print DEVI L_S1|Q2
.print DEVI L_S1|Q1
.print DEVI IT14|T
.print DEVI L_S2|A1
.print DEVI L_S2|A2
.print DEVI L_S2|A3
.print DEVI L_S2|B1
.print DEVI L_S2|B2
.print DEVI L_S2|B3
.print DEVI L_S2|T1
.print DEVI L_S2|T2
.print DEVI L_S2|Q2
.print DEVI L_S2|Q1
.print DEVI IT15|T
.print DEVI L_S3|A1
.print DEVI L_S3|A2
.print DEVI L_S3|A3
.print DEVI L_S3|B1
.print DEVI L_S3|B2
.print DEVI L_S3|B3
.print DEVI L_S3|T1
.print DEVI L_S3|T2
.print DEVI L_S3|Q2
.print DEVI L_S3|Q1
.print DEVI IT16|T
.print DEVI L_S4|1
.print DEVI L_S4|2
.print DEVI L_S4|3
.print DEVI L_S4|T
.print DEVI L_S4|4
.print DEVI L_S4|5
.print DEVI L_S4|6
.print V _DFF_IP2_12|A4
.print V IP1_0_TO1
.print V _S0|A1
.print V _DFF_IP2_01|A2
.print V SPL_IG2_0|QA1
.print V IP1_0_RX
.print V T02
.print V I3|A1
.print V P0_2_RX
.print V _PTL_G3_2|A_PTL_RX
.print V _S3|T1
.print V _DFF_IP1_12|T1
.print V _S0|T1
.print V T01
.print V _PG3_01|GG
.print V IP1_0
.print V _PTL_IP1_0|A_PTL
.print V I2|A2
.print V G2_2_RX
.print V SPL_IP3_0|D2
.print V S1
.print V _PTL_IG1_0|A_PTL
.print V _S1|Q1
.print V _PG2_12|G1_COPY_1
.print V _PTL_G0_2|A_PTL_RX
.print V _DFF_IP3_12|T1
.print V _S1|ABTQ
.print V I1|A2
.print V _DFF_IP3_01|Q1
.print V A2
.print V SPL_IG2_0|D2
.print V IG3_0_RX
.print V S0
.print V IP2_0_TO3
.print V _DFF_IP1_12|Q1
.print V _DFF_IP2_01|A4
.print V IP3_2_OUT
.print V IP2_1_OUT_RX
.print V _S3|B1
.print V IP3_0_TO1
.print V _S4|A2
.print V _S1|T2
.print V IP2_1_OUT
.print V I3|B2
.print V IG1_0_RX
.print V IP3_0_OUT
.print V G1_2
.print V _S1|B3
.print V _PG3_01|PG
.print V P0_1
.print V _DFF_IP3_01|A3
.print V _PG3_01|P1_SYNC
.print V _DFF_IP1_01|A4
.print V IP1_1_OUT
.print V G1_1_TO3
.print V G1_1_RX
.print V G1_1
.print V _S4|T1
.print V _PG1_12|T2
.print V _PTL_G2_2|A_PTL_RX
.print V _DFF_IP1_01|T2
.print V T09
.print V _S2|A2
.print V _PTL_IP1_1|A_PTL
.print V _S3|A2
.print V IP2_0_RX
.print V _PG1_01|G1_COPY_1
.print V I0|A2
.print V _PG3_12|GG_SYNC
.print V _PG1_12|A4
.print V _S3|Q1
.print V G0_1
.print V _S1|B1
.print V SPL_IP3_0|QB1
.print V _DFF_IP3_12|A1
.print V SPL_IP3_0|QA1
.print V _PTL_A1|A_PTL
.print V _S0|A2
.print V I0|B2
.print V _PTL_A0|A_PTL
.print V _DFF_IP2_12|Q1
.print V _PG1_01|GG
.print V _DFF_IP3_12|T2
.print V _DFF_IP2_12|T2
.print V I1|A1_SYNC
.print V I0|B1
.print V I3|B1_SYNC
.print V SPL_IP1_0|QB1
.print V _PTL_P2_1|A_PTL
.print V _PG1_01|PG
.print V _PTL_P0_2|A_PTL
.print V _S2|A3
.print V _PTL_P3_1|A_PTL
.print V _PTL_IP2_2|A_PTL
.print V _PG1_01|GG_SYNC
.print V _S3|ABTQ
.print V SPL_G1_1|QTMP
.print V _DFF_IP1_01|T1
.print V _PG1_12|A3
.print V _PG2_12|PG_SYNC
.print V _DFF_IP1_01|A3
.print V _PTL_IG0_0|A_PTL
.print V G3_2_RX
.print V _S4|A1
.print V _DFF_IP1_01|Q1
.print V _PTL_IP2_1|A_PTL
.print V T12
.print V _S2|T1
.print V IG0_0_TO0
.print V IG0_0_TO1
.print V _PTL_G3_2|A_PTL
.print V _S4|A3
.print V _S2|AB
.print V A1_RX
.print V _DFF_IP1_12|A2
.print V G1_1_TO2
.print V G2_1
.print V A3_RX
.print V SPL_IG2_0|QB1
.print V IG2_0_RX
.print V _DFF_IP1_01|A1
.print V SPL_IP2_0|QTMP
.print V _S1|AB
.print V IP0_0_RX
.print V _PTL_B0|A_PTL
.print V _PG1_12|A1
.print V _PTL_G3_1|A_PTL
.print V _S4|T2
.print V _DFF_IP3_12|A4
.print V I0|A1
.print V SPL_IP1_0|D1
.print V I2|B1
.print V _DFF_IP3_01|T1
.print V _PTL_G1_2|A_PTL
.print V T11
.print V _PTL_P0_2|A_PTL_RX
.print V P3_1
.print V P0_2
.print V _DFF_IP3_01|T2
.print V _S0|A4
.print V T05
.print V _DFF_IP2_01|A1
.print V G0_2_RX
.print V P2_1
.print V D11
.print V G2_1_RX
.print V IP2_2_OUT
.print V I0|B1_SYNC
.print V T06
.print V _S2|T2
.print V _DFF_IP2_12|A2
.print V T07
.print V _DFF_IP3_12|A2
.print V _S2|B3
.print V _PG1_12|A2
.print V T16
.print V _S3|B3
.print V _DFF_IP2_12|A1
.print V B1_RX
.print V I1|B1
.print V G2_2
.print V A2_RX
.print V G0_2
.print V _PG3_12|G1_COPY_2
.print V SPL_IP1_0|JCT
.print V _PTL_G2_2|A_PTL
.print V I2|B1_SYNC
.print V G1_2_RX
.print V _PTL_G0_2|A_PTL
.print V _PTL_B3|A_PTL
.print V _PTL_G0_1|A_PTL
.print V _S0|Q1
.print V SPL_IP3_0|D1
.print V SPL_IG2_0|JCT
.print V _S3|A3
.print V A3
.print V _DFF_IP1_12|A3
.print V T08
.print V _DFF_IP1_01|A2
.print V IP3_0
.print V _PG3_01|P1_COPY_2
.print V I1|B2
.print V IP1_0_OUT
.print V SPL_IG2_0|D1
.print V IG0_0
.print V G3_2
.print V _DFF_IP3_12|A3
.print V T10
.print V I2|A1
.print V I1|B1_SYNC
.print V _PTL_A2|A_PTL
.print V _PTL_G1_1|A_PTL
.print V _PTL_IP3_2|A_PTL
.print V _PTL_IP1_2|A_PTL
.print V _PTL_G2_1|A_PTL
.print V IP0_0
.print V _DFF_IP1_12|A1
.print V IP3_0_RX
.print V _S1|T1
.print V _PG2_12|G1_COPY_2
.print V I3|A1_SYNC
.print V _PG3_01|P1_COPY_1
.print V D12
.print V _S3|A1
.print V _PTL_IP2_2|A_PTL_RX
.print V IP2_0
.print V IP2_2_OUT_RX
.print V D13
.print V IG2_0
.print V _PTL_IP2_0|A_PTL
.print V P3_1_RX
.print V B2_RX
.print V IG2_0_TO3
.print V D03
.print V _PG3_01|G1_COPY_1
.print V _S1|B2
.print V _PG3_12|PG_SYNC
.print V _DFF_IP1_12|T2
.print V _PTL_IP1_2|A_PTL_RX
.print V SPL_IG0_0|QA1
.print V S4
.print V _PG3_12|GG
.print V _DFF_IP2_01|A3
.print V _PG3_01|GG_SYNC
.print V _PTL_IP3_2|A_PTL_RX
.print V D02
.print V _PTL_IP3_1|A_PTL
.print V _S3|T2
.print V _PTL_IP0_0|A_PTL
.print V _PG3_01|G1_COPY_2
.print V _PG3_01|PG_SYNC
.print V P0_1_RX
.print V _DFF_IP3_12|Q1
.print V SPL_IP3_0|JCT
.print V _S2|ABTQ
.print V SPL_IG0_0|QB1
.print V _S0|A3
.print V G1_1_TO1
.print V B3
.print V _PG1_01|PG_SYNC
.print V _PG3_12|G1_COPY_1
.print V _DFF_IP2_01|T1
.print V D01
.print V IG1_0
.print V _S3|B2
.print V _PG2_12|GG
.print V IG3_0
.print V _S2|A1
.print V _PG1_01|G1_COPY_2
.print V B0_RX
.print V SPL_IG0_0|D1
.print V G0_1_RX
.print V T00
.print V B1
.print V IP2_0_OUT
.print V I3|A2
.print V T15
.print V P2_1_RX
.print V IP3_2_OUT_RX
.print V A0_RX
.print V _DFF_IP1_12|A4
.print V T13
.print V IP1_2_OUT_RX
.print V _PTL_B2|A_PTL
.print V _DFF_IP3_01|A2
.print V _PTL_IG3_0|A_PTL
.print V _DFF_IP2_01|Q1
.print V G3_1
.print V _PTL_IP3_0|A_PTL
.print V S3
.print V IP1_2_OUT
.print V _PG1_12|Q1
.print V _PTL_G1_2|A_PTL_RX
.print V I2|B2
.print V SPL_IP1_0|QA1
.print V T14
.print V IP1_1_OUT_RX
.print V B0
.print V _PTL_P0_1|A_PTL
.print V IG0_0_RX
.print V _S4|A4
.print V IG2_0_TO2
.print V _DFF_IP2_12|T1
.print V _PG1_12|T1
.print V IP3_1_OUT
.print V _PG3_12|PG
.print V _S1|A2
.print V _S3|AB
.print V _S1|A3
.print V I2|A1_SYNC
.print V IP2_0_TO2
.print V I0|A1_SYNC
.print V _DFF_IP3_01|A4
.print V _PG2_12|PG
.print V A1
.print V _DFF_IP2_01|T2
.print V S2
.print V _S4|Q1
.print V _PG3_01|P0_SYNC
.print V SPL_IG0_0|JCT
.print V _S0|T2
.print V _PTL_A3|A_PTL
.print V _S2|B2
.print V I3|B1
.print V _S2|B1
.print V _DFF_IP3_01|A1
.print V T04
.print V _S1|A1
.print V I1|A1
.print V SPL_IP1_0|D2
.print V _DFF_IP2_12|A3
.print V _PTL_B1|A_PTL
.print V _PG2_12|GG_SYNC
.print V SPL_IG0_0|D2
.print V B3_RX
.print V IP3_1_OUT_RX
.print V _PTL_IG2_0|A_PTL
.print V A0
.print V _S2|Q1
.print V T03
.print V G3_1_RX
.print V B2
