*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM TCLOCK=2e-10
.PARAM OS=5.0000000000000005e-12
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 54000E-12
R_P0_1 P0_1 0  1
R_G0_1 G0_1 0  1
R_P1_1_TO1 P1_1_TO1 0  1
R_P1_1_TO2 P1_1_TO2 0  1
R_P1_1_TO3 P1_1_TO3 0  1
R_G1_1_TO1 G1_1_TO1 0  1
R_G1_1_TO2 G1_1_TO2 0  1
R_G1_1_TO3 G1_1_TO3 0  1
R_P2_1 P2_1 0  1
R_G2_1 G2_1 0  1
R_P3_1 P3_1 0  1
R_G3_1 G3_1 0  1
R_IP1_1 IP1_1_OUT 0  1
R_IP2_1 IP2_1_OUT 0  1
R_IP3_1 IP3_1_OUT 0  1
IA0_|A 0 A0_  PWL(0 0 3.55e-11 0 3.7e-11 0.0013786 3.85e-11 0 4.355e-10 0 4.37e-10 0.0013786 4.385e-10 0 8.355e-10 0 8.37e-10 0.0013786 8.385e-10 0 1.2355e-09 0 1.237e-09 0.0013786 1.2385e-09 0 1.6355e-09 0 1.637e-09 0.0013786 1.6385e-09 0 2.0355e-09 0 2.037e-09 0.0013786 2.0385e-09 0 2.4355e-09 0 2.437e-09 0.0013786 2.4385e-09 0 2.8355e-09 0 2.837e-09 0.0013786 2.8385e-09 0 3.2355e-09 0 3.237e-09 0.0013786 3.2385e-09 0 3.6355e-09 0 3.637e-09 0.0013786 3.6385e-09 0 4.0355e-09 0 4.037e-09 0.0013786 4.0385e-09 0 4.4355e-09 0 4.437e-09 0.0013786 4.4385e-09 0 4.8355e-09 0 4.837e-09 0.0013786 4.8385e-09 0 5.2355e-09 0 5.237e-09 0.0013786 5.2385e-09 0 5.6355e-09 0 5.637e-09 0.0013786 5.6385e-09 0 6.0355e-09 0 6.037e-09 0.0013786 6.0385e-09 0 6.4355e-09 0 6.437e-09 0.0013786 6.4385e-09 0 6.8355e-09 0 6.837e-09 0.0013786 6.8385e-09 0 7.2355e-09 0 7.237e-09 0.0013786 7.2385e-09 0 7.6355e-09 0 7.637e-09 0.0013786 7.6385e-09 0 8.0355e-09 0 8.037e-09 0.0013786 8.0385e-09 0 8.4355e-09 0 8.437e-09 0.0013786 8.4385e-09 0 8.8355e-09 0 8.837e-09 0.0013786 8.8385e-09 0 9.2355e-09 0 9.237e-09 0.0013786 9.2385e-09 0 9.6355e-09 0 9.637e-09 0.0013786 9.6385e-09 0 1.00355e-08 0 1.0037e-08 0.0013786 1.00385e-08 0 1.04355e-08 0 1.0437e-08 0.0013786 1.04385e-08 0 1.08355e-08 0 1.0837e-08 0.0013786 1.08385e-08 0 1.12355e-08 0 1.1237e-08 0.0013786 1.12385e-08 0 1.16355e-08 0 1.1637e-08 0.0013786 1.16385e-08 0 1.20355e-08 0 1.2037e-08 0.0013786 1.20385e-08 0 1.24355e-08 0 1.2437e-08 0.0013786 1.24385e-08 0 1.28355e-08 0 1.2837e-08 0.0013786 1.28385e-08 0 1.32355e-08 0 1.3237e-08 0.0013786 1.32385e-08 0 1.36355e-08 0 1.3637e-08 0.0013786 1.36385e-08 0 1.40355e-08 0 1.4037e-08 0.0013786 1.40385e-08 0 1.44355e-08 0 1.4437e-08 0.0013786 1.44385e-08 0 1.48355e-08 0 1.4837e-08 0.0013786 1.48385e-08 0 1.52355e-08 0 1.5237e-08 0.0013786 1.52385e-08 0 1.56355e-08 0 1.5637e-08 0.0013786 1.56385e-08 0 1.60355e-08 0 1.6037e-08 0.0013786 1.60385e-08 0 1.64355e-08 0 1.6437e-08 0.0013786 1.64385e-08 0 1.68355e-08 0 1.6837e-08 0.0013786 1.68385e-08 0 1.72355e-08 0 1.7237e-08 0.0013786 1.72385e-08 0 1.76355e-08 0 1.7637e-08 0.0013786 1.76385e-08 0 1.80355e-08 0 1.8037e-08 0.0013786 1.80385e-08 0 1.84355e-08 0 1.8437e-08 0.0013786 1.84385e-08 0 1.88355e-08 0 1.8837e-08 0.0013786 1.88385e-08 0 1.92355e-08 0 1.9237e-08 0.0013786 1.92385e-08 0 1.96355e-08 0 1.9637e-08 0.0013786 1.96385e-08 0 2.00355e-08 0 2.0037e-08 0.0013786 2.00385e-08 0 2.04355e-08 0 2.0437e-08 0.0013786 2.04385e-08 0 2.08355e-08 0 2.0837e-08 0.0013786 2.08385e-08 0 2.12355e-08 0 2.1237e-08 0.0013786 2.12385e-08 0 2.16355e-08 0 2.1637e-08 0.0013786 2.16385e-08 0 2.20355e-08 0 2.2037e-08 0.0013786 2.20385e-08 0 2.24355e-08 0 2.2437e-08 0.0013786 2.24385e-08 0 2.28355e-08 0 2.2837e-08 0.0013786 2.28385e-08 0 2.32355e-08 0 2.3237e-08 0.0013786 2.32385e-08 0 2.36355e-08 0 2.3637e-08 0.0013786 2.36385e-08 0 2.40355e-08 0 2.4037e-08 0.0013786 2.40385e-08 0 2.44355e-08 0 2.4437e-08 0.0013786 2.44385e-08 0 2.48355e-08 0 2.4837e-08 0.0013786 2.48385e-08 0 2.52355e-08 0 2.5237e-08 0.0013786 2.52385e-08 0 2.56355e-08 0 2.5637e-08 0.0013786 2.56385e-08 0 2.60355e-08 0 2.6037e-08 0.0013786 2.60385e-08 0 2.64355e-08 0 2.6437e-08 0.0013786 2.64385e-08 0 2.68355e-08 0 2.6837e-08 0.0013786 2.68385e-08 0 2.72355e-08 0 2.7237e-08 0.0013786 2.72385e-08 0 2.76355e-08 0 2.7637e-08 0.0013786 2.76385e-08 0 2.80355e-08 0 2.8037e-08 0.0013786 2.80385e-08 0 2.84355e-08 0 2.8437e-08 0.0013786 2.84385e-08 0 2.88355e-08 0 2.8837e-08 0.0013786 2.88385e-08 0 2.92355e-08 0 2.9237e-08 0.0013786 2.92385e-08 0 2.96355e-08 0 2.9637e-08 0.0013786 2.96385e-08 0 3.00355e-08 0 3.0037e-08 0.0013786 3.00385e-08 0 3.04355e-08 0 3.0437e-08 0.0013786 3.04385e-08 0 3.08355e-08 0 3.0837e-08 0.0013786 3.08385e-08 0 3.12355e-08 0 3.1237e-08 0.0013786 3.12385e-08 0 3.16355e-08 0 3.1637e-08 0.0013786 3.16385e-08 0 3.20355e-08 0 3.2037e-08 0.0013786 3.20385e-08 0 3.24355e-08 0 3.2437e-08 0.0013786 3.24385e-08 0 3.28355e-08 0 3.2837e-08 0.0013786 3.28385e-08 0 3.32355e-08 0 3.3237e-08 0.0013786 3.32385e-08 0 3.36355e-08 0 3.3637e-08 0.0013786 3.36385e-08 0 3.40355e-08 0 3.4037e-08 0.0013786 3.40385e-08 0 3.44355e-08 0 3.4437e-08 0.0013786 3.44385e-08 0 3.48355e-08 0 3.4837e-08 0.0013786 3.48385e-08 0 3.52355e-08 0 3.5237e-08 0.0013786 3.52385e-08 0 3.56355e-08 0 3.5637e-08 0.0013786 3.56385e-08 0 3.60355e-08 0 3.6037e-08 0.0013786 3.60385e-08 0 3.64355e-08 0 3.6437e-08 0.0013786 3.64385e-08 0 3.68355e-08 0 3.6837e-08 0.0013786 3.68385e-08 0 3.72355e-08 0 3.7237e-08 0.0013786 3.72385e-08 0 3.76355e-08 0 3.7637e-08 0.0013786 3.76385e-08 0 3.80355e-08 0 3.8037e-08 0.0013786 3.80385e-08 0 3.84355e-08 0 3.8437e-08 0.0013786 3.84385e-08 0 3.88355e-08 0 3.8837e-08 0.0013786 3.88385e-08 0 3.92355e-08 0 3.9237e-08 0.0013786 3.92385e-08 0 3.96355e-08 0 3.9637e-08 0.0013786 3.96385e-08 0 4.00355e-08 0 4.0037e-08 0.0013786 4.00385e-08 0 4.04355e-08 0 4.0437e-08 0.0013786 4.04385e-08 0 4.08355e-08 0 4.0837e-08 0.0013786 4.08385e-08 0 4.12355e-08 0 4.1237e-08 0.0013786 4.12385e-08 0 4.16355e-08 0 4.1637e-08 0.0013786 4.16385e-08 0 4.20355e-08 0 4.2037e-08 0.0013786 4.20385e-08 0 4.24355e-08 0 4.2437e-08 0.0013786 4.24385e-08 0 4.28355e-08 0 4.2837e-08 0.0013786 4.28385e-08 0 4.32355e-08 0 4.3237e-08 0.0013786 4.32385e-08 0 4.36355e-08 0 4.3637e-08 0.0013786 4.36385e-08 0 4.40355e-08 0 4.4037e-08 0.0013786 4.40385e-08 0 4.44355e-08 0 4.4437e-08 0.0013786 4.44385e-08 0 4.48355e-08 0 4.4837e-08 0.0013786 4.48385e-08 0 4.52355e-08 0 4.5237e-08 0.0013786 4.52385e-08 0 4.56355e-08 0 4.5637e-08 0.0013786 4.56385e-08 0 4.60355e-08 0 4.6037e-08 0.0013786 4.60385e-08 0 4.64355e-08 0 4.6437e-08 0.0013786 4.64385e-08 0 4.68355e-08 0 4.6837e-08 0.0013786 4.68385e-08 0 4.72355e-08 0 4.7237e-08 0.0013786 4.72385e-08 0 4.76355e-08 0 4.7637e-08 0.0013786 4.76385e-08 0 4.80355e-08 0 4.8037e-08 0.0013786 4.80385e-08 0 4.84355e-08 0 4.8437e-08 0.0013786 4.84385e-08 0 4.88355e-08 0 4.8837e-08 0.0013786 4.88385e-08 0 4.92355e-08 0 4.9237e-08 0.0013786 4.92385e-08 0 4.96355e-08 0 4.9637e-08 0.0013786 4.96385e-08 0 5.00355e-08 0 5.0037e-08 0.0013786 5.00385e-08 0 5.04355e-08 0 5.0437e-08 0.0013786 5.04385e-08 0 5.08355e-08 0 5.0837e-08 0.0013786 5.08385e-08 0)
IB0_|B 0 B0_  PWL(0 0 5.15e-11 0 5.3e-11 0.0013786 5.45e-11 0 2.515e-10 0 2.53e-10 0.0013786 2.545e-10 0 8.515e-10 0 8.53e-10 0.0013786 8.545e-10 0 1.0515e-09 0 1.053e-09 0.0013786 1.0545e-09 0 1.6515e-09 0 1.653e-09 0.0013786 1.6545e-09 0 1.8515e-09 0 1.853e-09 0.0013786 1.8545e-09 0 2.4515e-09 0 2.453e-09 0.0013786 2.4545e-09 0 2.6515e-09 0 2.653e-09 0.0013786 2.6545e-09 0 3.2515e-09 0 3.253e-09 0.0013786 3.2545e-09 0 3.4515e-09 0 3.453e-09 0.0013786 3.4545e-09 0 4.0515e-09 0 4.053e-09 0.0013786 4.0545e-09 0 4.2515e-09 0 4.253e-09 0.0013786 4.2545e-09 0 4.8515e-09 0 4.853e-09 0.0013786 4.8545e-09 0 5.0515e-09 0 5.053e-09 0.0013786 5.0545e-09 0 5.6515e-09 0 5.653e-09 0.0013786 5.6545e-09 0 5.8515e-09 0 5.853e-09 0.0013786 5.8545e-09 0 6.4515e-09 0 6.453e-09 0.0013786 6.4545e-09 0 6.6515e-09 0 6.653e-09 0.0013786 6.6545e-09 0 7.2515e-09 0 7.253e-09 0.0013786 7.2545e-09 0 7.4515e-09 0 7.453e-09 0.0013786 7.4545e-09 0 8.0515e-09 0 8.053e-09 0.0013786 8.0545e-09 0 8.2515e-09 0 8.253e-09 0.0013786 8.2545e-09 0 8.8515e-09 0 8.853e-09 0.0013786 8.8545e-09 0 9.0515e-09 0 9.053e-09 0.0013786 9.0545e-09 0 9.6515e-09 0 9.653e-09 0.0013786 9.6545e-09 0 9.8515e-09 0 9.853e-09 0.0013786 9.8545e-09 0 1.04515e-08 0 1.0453e-08 0.0013786 1.04545e-08 0 1.06515e-08 0 1.0653e-08 0.0013786 1.06545e-08 0 1.12515e-08 0 1.1253e-08 0.0013786 1.12545e-08 0 1.14515e-08 0 1.1453e-08 0.0013786 1.14545e-08 0 1.20515e-08 0 1.2053e-08 0.0013786 1.20545e-08 0 1.22515e-08 0 1.2253e-08 0.0013786 1.22545e-08 0 1.28515e-08 0 1.2853e-08 0.0013786 1.28545e-08 0 1.30515e-08 0 1.3053e-08 0.0013786 1.30545e-08 0 1.36515e-08 0 1.3653e-08 0.0013786 1.36545e-08 0 1.38515e-08 0 1.3853e-08 0.0013786 1.38545e-08 0 1.44515e-08 0 1.4453e-08 0.0013786 1.44545e-08 0 1.46515e-08 0 1.4653e-08 0.0013786 1.46545e-08 0 1.52515e-08 0 1.5253e-08 0.0013786 1.52545e-08 0 1.54515e-08 0 1.5453e-08 0.0013786 1.54545e-08 0 1.60515e-08 0 1.6053e-08 0.0013786 1.60545e-08 0 1.62515e-08 0 1.6253e-08 0.0013786 1.62545e-08 0 1.68515e-08 0 1.6853e-08 0.0013786 1.68545e-08 0 1.70515e-08 0 1.7053e-08 0.0013786 1.70545e-08 0 1.76515e-08 0 1.7653e-08 0.0013786 1.76545e-08 0 1.78515e-08 0 1.7853e-08 0.0013786 1.78545e-08 0 1.84515e-08 0 1.8453e-08 0.0013786 1.84545e-08 0 1.86515e-08 0 1.8653e-08 0.0013786 1.86545e-08 0 1.92515e-08 0 1.9253e-08 0.0013786 1.92545e-08 0 1.94515e-08 0 1.9453e-08 0.0013786 1.94545e-08 0 2.00515e-08 0 2.0053e-08 0.0013786 2.00545e-08 0 2.02515e-08 0 2.0253e-08 0.0013786 2.02545e-08 0 2.08515e-08 0 2.0853e-08 0.0013786 2.08545e-08 0 2.10515e-08 0 2.1053e-08 0.0013786 2.10545e-08 0 2.16515e-08 0 2.1653e-08 0.0013786 2.16545e-08 0 2.18515e-08 0 2.1853e-08 0.0013786 2.18545e-08 0 2.24515e-08 0 2.2453e-08 0.0013786 2.24545e-08 0 2.26515e-08 0 2.2653e-08 0.0013786 2.26545e-08 0 2.32515e-08 0 2.3253e-08 0.0013786 2.32545e-08 0 2.34515e-08 0 2.3453e-08 0.0013786 2.34545e-08 0 2.40515e-08 0 2.4053e-08 0.0013786 2.40545e-08 0 2.42515e-08 0 2.4253e-08 0.0013786 2.42545e-08 0 2.48515e-08 0 2.4853e-08 0.0013786 2.48545e-08 0 2.50515e-08 0 2.5053e-08 0.0013786 2.50545e-08 0 2.56515e-08 0 2.5653e-08 0.0013786 2.56545e-08 0 2.58515e-08 0 2.5853e-08 0.0013786 2.58545e-08 0 2.64515e-08 0 2.6453e-08 0.0013786 2.64545e-08 0 2.66515e-08 0 2.6653e-08 0.0013786 2.66545e-08 0 2.72515e-08 0 2.7253e-08 0.0013786 2.72545e-08 0 2.74515e-08 0 2.7453e-08 0.0013786 2.74545e-08 0 2.80515e-08 0 2.8053e-08 0.0013786 2.80545e-08 0 2.82515e-08 0 2.8253e-08 0.0013786 2.82545e-08 0 2.88515e-08 0 2.8853e-08 0.0013786 2.88545e-08 0 2.90515e-08 0 2.9053e-08 0.0013786 2.90545e-08 0 2.96515e-08 0 2.9653e-08 0.0013786 2.96545e-08 0 2.98515e-08 0 2.9853e-08 0.0013786 2.98545e-08 0 3.04515e-08 0 3.0453e-08 0.0013786 3.04545e-08 0 3.06515e-08 0 3.0653e-08 0.0013786 3.06545e-08 0 3.12515e-08 0 3.1253e-08 0.0013786 3.12545e-08 0 3.14515e-08 0 3.1453e-08 0.0013786 3.14545e-08 0 3.20515e-08 0 3.2053e-08 0.0013786 3.20545e-08 0 3.22515e-08 0 3.2253e-08 0.0013786 3.22545e-08 0 3.28515e-08 0 3.2853e-08 0.0013786 3.28545e-08 0 3.30515e-08 0 3.3053e-08 0.0013786 3.30545e-08 0 3.36515e-08 0 3.3653e-08 0.0013786 3.36545e-08 0 3.38515e-08 0 3.3853e-08 0.0013786 3.38545e-08 0 3.44515e-08 0 3.4453e-08 0.0013786 3.44545e-08 0 3.46515e-08 0 3.4653e-08 0.0013786 3.46545e-08 0 3.52515e-08 0 3.5253e-08 0.0013786 3.52545e-08 0 3.54515e-08 0 3.5453e-08 0.0013786 3.54545e-08 0 3.60515e-08 0 3.6053e-08 0.0013786 3.60545e-08 0 3.62515e-08 0 3.6253e-08 0.0013786 3.62545e-08 0 3.68515e-08 0 3.6853e-08 0.0013786 3.68545e-08 0 3.70515e-08 0 3.7053e-08 0.0013786 3.70545e-08 0 3.76515e-08 0 3.7653e-08 0.0013786 3.76545e-08 0 3.78515e-08 0 3.7853e-08 0.0013786 3.78545e-08 0 3.84515e-08 0 3.8453e-08 0.0013786 3.84545e-08 0 3.86515e-08 0 3.8653e-08 0.0013786 3.86545e-08 0 3.92515e-08 0 3.9253e-08 0.0013786 3.92545e-08 0 3.94515e-08 0 3.9453e-08 0.0013786 3.94545e-08 0 4.00515e-08 0 4.0053e-08 0.0013786 4.00545e-08 0 4.02515e-08 0 4.0253e-08 0.0013786 4.02545e-08 0 4.08515e-08 0 4.0853e-08 0.0013786 4.08545e-08 0 4.10515e-08 0 4.1053e-08 0.0013786 4.10545e-08 0 4.16515e-08 0 4.1653e-08 0.0013786 4.16545e-08 0 4.18515e-08 0 4.1853e-08 0.0013786 4.18545e-08 0 4.24515e-08 0 4.2453e-08 0.0013786 4.24545e-08 0 4.26515e-08 0 4.2653e-08 0.0013786 4.26545e-08 0 4.32515e-08 0 4.3253e-08 0.0013786 4.32545e-08 0 4.34515e-08 0 4.3453e-08 0.0013786 4.34545e-08 0 4.40515e-08 0 4.4053e-08 0.0013786 4.40545e-08 0 4.42515e-08 0 4.4253e-08 0.0013786 4.42545e-08 0 4.48515e-08 0 4.4853e-08 0.0013786 4.48545e-08 0 4.50515e-08 0 4.5053e-08 0.0013786 4.50545e-08 0 4.56515e-08 0 4.5653e-08 0.0013786 4.56545e-08 0 4.58515e-08 0 4.5853e-08 0.0013786 4.58545e-08 0 4.64515e-08 0 4.6453e-08 0.0013786 4.64545e-08 0 4.66515e-08 0 4.6653e-08 0.0013786 4.66545e-08 0 4.72515e-08 0 4.7253e-08 0.0013786 4.72545e-08 0 4.74515e-08 0 4.7453e-08 0.0013786 4.74545e-08 0 4.80515e-08 0 4.8053e-08 0.0013786 4.80545e-08 0 4.82515e-08 0 4.8253e-08 0.0013786 4.82545e-08 0 4.88515e-08 0 4.8853e-08 0.0013786 4.88545e-08 0 4.90515e-08 0 4.9053e-08 0.0013786 4.90545e-08 0 4.96515e-08 0 4.9653e-08 0.0013786 4.96545e-08 0 4.98515e-08 0 4.9853e-08 0.0013786 4.98545e-08 0 5.04515e-08 0 5.0453e-08 0.0013786 5.04545e-08 0 5.06515e-08 0 5.0653e-08 0.0013786 5.06545e-08 0)
IA1_|C 0 A1_  PWL(0 0 6.75e-11 0 6.9e-11 0.0013786 7.05e-11 0 2.675e-10 0 2.69e-10 0.0013786 2.705e-10 0 4.675e-10 0 4.69e-10 0.0013786 4.705e-10 0 6.675e-10 0 6.69e-10 0.0013786 6.705e-10 0 1.6675e-09 0 1.669e-09 0.0013786 1.6705e-09 0 1.8675e-09 0 1.869e-09 0.0013786 1.8705e-09 0 2.0675e-09 0 2.069e-09 0.0013786 2.0705e-09 0 2.2675e-09 0 2.269e-09 0.0013786 2.2705e-09 0 3.2675e-09 0 3.269e-09 0.0013786 3.2705e-09 0 3.4675e-09 0 3.469e-09 0.0013786 3.4705e-09 0 3.6675e-09 0 3.669e-09 0.0013786 3.6705e-09 0 3.8675e-09 0 3.869e-09 0.0013786 3.8705e-09 0 4.8675e-09 0 4.869e-09 0.0013786 4.8705e-09 0 5.0675e-09 0 5.069e-09 0.0013786 5.0705e-09 0 5.2675e-09 0 5.269e-09 0.0013786 5.2705e-09 0 5.4675e-09 0 5.469e-09 0.0013786 5.4705e-09 0 6.4675e-09 0 6.469e-09 0.0013786 6.4705e-09 0 6.6675e-09 0 6.669e-09 0.0013786 6.6705e-09 0 6.8675e-09 0 6.869e-09 0.0013786 6.8705e-09 0 7.0675e-09 0 7.069e-09 0.0013786 7.0705e-09 0 8.0675e-09 0 8.069e-09 0.0013786 8.0705e-09 0 8.2675e-09 0 8.269e-09 0.0013786 8.2705e-09 0 8.4675e-09 0 8.469e-09 0.0013786 8.4705e-09 0 8.6675e-09 0 8.669e-09 0.0013786 8.6705e-09 0 9.6675e-09 0 9.669e-09 0.0013786 9.6705e-09 0 9.8675e-09 0 9.869e-09 0.0013786 9.8705e-09 0 1.00675e-08 0 1.0069e-08 0.0013786 1.00705e-08 0 1.02675e-08 0 1.0269e-08 0.0013786 1.02705e-08 0 1.12675e-08 0 1.1269e-08 0.0013786 1.12705e-08 0 1.14675e-08 0 1.1469e-08 0.0013786 1.14705e-08 0 1.16675e-08 0 1.1669e-08 0.0013786 1.16705e-08 0 1.18675e-08 0 1.1869e-08 0.0013786 1.18705e-08 0 1.28675e-08 0 1.2869e-08 0.0013786 1.28705e-08 0 1.30675e-08 0 1.3069e-08 0.0013786 1.30705e-08 0 1.32675e-08 0 1.3269e-08 0.0013786 1.32705e-08 0 1.34675e-08 0 1.3469e-08 0.0013786 1.34705e-08 0 1.44675e-08 0 1.4469e-08 0.0013786 1.44705e-08 0 1.46675e-08 0 1.4669e-08 0.0013786 1.46705e-08 0 1.48675e-08 0 1.4869e-08 0.0013786 1.48705e-08 0 1.50675e-08 0 1.5069e-08 0.0013786 1.50705e-08 0 1.60675e-08 0 1.6069e-08 0.0013786 1.60705e-08 0 1.62675e-08 0 1.6269e-08 0.0013786 1.62705e-08 0 1.64675e-08 0 1.6469e-08 0.0013786 1.64705e-08 0 1.66675e-08 0 1.6669e-08 0.0013786 1.66705e-08 0 1.76675e-08 0 1.7669e-08 0.0013786 1.76705e-08 0 1.78675e-08 0 1.7869e-08 0.0013786 1.78705e-08 0 1.80675e-08 0 1.8069e-08 0.0013786 1.80705e-08 0 1.82675e-08 0 1.8269e-08 0.0013786 1.82705e-08 0 1.92675e-08 0 1.9269e-08 0.0013786 1.92705e-08 0 1.94675e-08 0 1.9469e-08 0.0013786 1.94705e-08 0 1.96675e-08 0 1.9669e-08 0.0013786 1.96705e-08 0 1.98675e-08 0 1.9869e-08 0.0013786 1.98705e-08 0 2.08675e-08 0 2.0869e-08 0.0013786 2.08705e-08 0 2.10675e-08 0 2.1069e-08 0.0013786 2.10705e-08 0 2.12675e-08 0 2.1269e-08 0.0013786 2.12705e-08 0 2.14675e-08 0 2.1469e-08 0.0013786 2.14705e-08 0 2.24675e-08 0 2.2469e-08 0.0013786 2.24705e-08 0 2.26675e-08 0 2.2669e-08 0.0013786 2.26705e-08 0 2.28675e-08 0 2.2869e-08 0.0013786 2.28705e-08 0 2.30675e-08 0 2.3069e-08 0.0013786 2.30705e-08 0 2.40675e-08 0 2.4069e-08 0.0013786 2.40705e-08 0 2.42675e-08 0 2.4269e-08 0.0013786 2.42705e-08 0 2.44675e-08 0 2.4469e-08 0.0013786 2.44705e-08 0 2.46675e-08 0 2.4669e-08 0.0013786 2.46705e-08 0 2.56675e-08 0 2.5669e-08 0.0013786 2.56705e-08 0 2.58675e-08 0 2.5869e-08 0.0013786 2.58705e-08 0 2.60675e-08 0 2.6069e-08 0.0013786 2.60705e-08 0 2.62675e-08 0 2.6269e-08 0.0013786 2.62705e-08 0 2.72675e-08 0 2.7269e-08 0.0013786 2.72705e-08 0 2.74675e-08 0 2.7469e-08 0.0013786 2.74705e-08 0 2.76675e-08 0 2.7669e-08 0.0013786 2.76705e-08 0 2.78675e-08 0 2.7869e-08 0.0013786 2.78705e-08 0 2.88675e-08 0 2.8869e-08 0.0013786 2.88705e-08 0 2.90675e-08 0 2.9069e-08 0.0013786 2.90705e-08 0 2.92675e-08 0 2.9269e-08 0.0013786 2.92705e-08 0 2.94675e-08 0 2.9469e-08 0.0013786 2.94705e-08 0 3.04675e-08 0 3.0469e-08 0.0013786 3.04705e-08 0 3.06675e-08 0 3.0669e-08 0.0013786 3.06705e-08 0 3.08675e-08 0 3.0869e-08 0.0013786 3.08705e-08 0 3.10675e-08 0 3.1069e-08 0.0013786 3.10705e-08 0 3.20675e-08 0 3.2069e-08 0.0013786 3.20705e-08 0 3.22675e-08 0 3.2269e-08 0.0013786 3.22705e-08 0 3.24675e-08 0 3.2469e-08 0.0013786 3.24705e-08 0 3.26675e-08 0 3.2669e-08 0.0013786 3.26705e-08 0 3.36675e-08 0 3.3669e-08 0.0013786 3.36705e-08 0 3.38675e-08 0 3.3869e-08 0.0013786 3.38705e-08 0 3.40675e-08 0 3.4069e-08 0.0013786 3.40705e-08 0 3.42675e-08 0 3.4269e-08 0.0013786 3.42705e-08 0 3.52675e-08 0 3.5269e-08 0.0013786 3.52705e-08 0 3.54675e-08 0 3.5469e-08 0.0013786 3.54705e-08 0 3.56675e-08 0 3.5669e-08 0.0013786 3.56705e-08 0 3.58675e-08 0 3.5869e-08 0.0013786 3.58705e-08 0 3.68675e-08 0 3.6869e-08 0.0013786 3.68705e-08 0 3.70675e-08 0 3.7069e-08 0.0013786 3.70705e-08 0 3.72675e-08 0 3.7269e-08 0.0013786 3.72705e-08 0 3.74675e-08 0 3.7469e-08 0.0013786 3.74705e-08 0 3.84675e-08 0 3.8469e-08 0.0013786 3.84705e-08 0 3.86675e-08 0 3.8669e-08 0.0013786 3.86705e-08 0 3.88675e-08 0 3.8869e-08 0.0013786 3.88705e-08 0 3.90675e-08 0 3.9069e-08 0.0013786 3.90705e-08 0 4.00675e-08 0 4.0069e-08 0.0013786 4.00705e-08 0 4.02675e-08 0 4.0269e-08 0.0013786 4.02705e-08 0 4.04675e-08 0 4.0469e-08 0.0013786 4.04705e-08 0 4.06675e-08 0 4.0669e-08 0.0013786 4.06705e-08 0 4.16675e-08 0 4.1669e-08 0.0013786 4.16705e-08 0 4.18675e-08 0 4.1869e-08 0.0013786 4.18705e-08 0 4.20675e-08 0 4.2069e-08 0.0013786 4.20705e-08 0 4.22675e-08 0 4.2269e-08 0.0013786 4.22705e-08 0 4.32675e-08 0 4.3269e-08 0.0013786 4.32705e-08 0 4.34675e-08 0 4.3469e-08 0.0013786 4.34705e-08 0 4.36675e-08 0 4.3669e-08 0.0013786 4.36705e-08 0 4.38675e-08 0 4.3869e-08 0.0013786 4.38705e-08 0 4.48675e-08 0 4.4869e-08 0.0013786 4.48705e-08 0 4.50675e-08 0 4.5069e-08 0.0013786 4.50705e-08 0 4.52675e-08 0 4.5269e-08 0.0013786 4.52705e-08 0 4.54675e-08 0 4.5469e-08 0.0013786 4.54705e-08 0 4.64675e-08 0 4.6469e-08 0.0013786 4.64705e-08 0 4.66675e-08 0 4.6669e-08 0.0013786 4.66705e-08 0 4.68675e-08 0 4.6869e-08 0.0013786 4.68705e-08 0 4.70675e-08 0 4.7069e-08 0.0013786 4.70705e-08 0 4.80675e-08 0 4.8069e-08 0.0013786 4.80705e-08 0 4.82675e-08 0 4.8269e-08 0.0013786 4.82705e-08 0 4.84675e-08 0 4.8469e-08 0.0013786 4.84705e-08 0 4.86675e-08 0 4.8669e-08 0.0013786 4.86705e-08 0 4.96675e-08 0 4.9669e-08 0.0013786 4.96705e-08 0 4.98675e-08 0 4.9869e-08 0.0013786 4.98705e-08 0 5.00675e-08 0 5.0069e-08 0.0013786 5.00705e-08 0 5.02675e-08 0 5.0269e-08 0.0013786 5.02705e-08 0)
IB1_|D 0 B1_  PWL(0 0 8.35e-11 0 8.5e-11 0.0013786 8.65e-11 0 2.835e-10 0 2.85e-10 0.0013786 2.865e-10 0 4.835e-10 0 4.85e-10 0.0013786 4.865e-10 0 6.835e-10 0 6.85e-10 0.0013786 6.865e-10 0 8.835e-10 0 8.85e-10 0.0013786 8.865e-10 0 1.0835e-09 0 1.085e-09 0.0013786 1.0865e-09 0 1.2835e-09 0 1.285e-09 0.0013786 1.2865e-09 0 1.4835e-09 0 1.485e-09 0.0013786 1.4865e-09 0 3.2835e-09 0 3.285e-09 0.0013786 3.2865e-09 0 3.4835e-09 0 3.485e-09 0.0013786 3.4865e-09 0 3.6835e-09 0 3.685e-09 0.0013786 3.6865e-09 0 3.8835e-09 0 3.885e-09 0.0013786 3.8865e-09 0 4.0835e-09 0 4.085e-09 0.0013786 4.0865e-09 0 4.2835e-09 0 4.285e-09 0.0013786 4.2865e-09 0 4.4835e-09 0 4.485e-09 0.0013786 4.4865e-09 0 4.6835e-09 0 4.685e-09 0.0013786 4.6865e-09 0 6.4835e-09 0 6.485e-09 0.0013786 6.4865e-09 0 6.6835e-09 0 6.685e-09 0.0013786 6.6865e-09 0 6.8835e-09 0 6.885e-09 0.0013786 6.8865e-09 0 7.0835e-09 0 7.085e-09 0.0013786 7.0865e-09 0 7.2835e-09 0 7.285e-09 0.0013786 7.2865e-09 0 7.4835e-09 0 7.485e-09 0.0013786 7.4865e-09 0 7.6835e-09 0 7.685e-09 0.0013786 7.6865e-09 0 7.8835e-09 0 7.885e-09 0.0013786 7.8865e-09 0 9.6835e-09 0 9.685e-09 0.0013786 9.6865e-09 0 9.8835e-09 0 9.885e-09 0.0013786 9.8865e-09 0 1.00835e-08 0 1.0085e-08 0.0013786 1.00865e-08 0 1.02835e-08 0 1.0285e-08 0.0013786 1.02865e-08 0 1.04835e-08 0 1.0485e-08 0.0013786 1.04865e-08 0 1.06835e-08 0 1.0685e-08 0.0013786 1.06865e-08 0 1.08835e-08 0 1.0885e-08 0.0013786 1.08865e-08 0 1.10835e-08 0 1.1085e-08 0.0013786 1.10865e-08 0 1.28835e-08 0 1.2885e-08 0.0013786 1.28865e-08 0 1.30835e-08 0 1.3085e-08 0.0013786 1.30865e-08 0 1.32835e-08 0 1.3285e-08 0.0013786 1.32865e-08 0 1.34835e-08 0 1.3485e-08 0.0013786 1.34865e-08 0 1.36835e-08 0 1.3685e-08 0.0013786 1.36865e-08 0 1.38835e-08 0 1.3885e-08 0.0013786 1.38865e-08 0 1.40835e-08 0 1.4085e-08 0.0013786 1.40865e-08 0 1.42835e-08 0 1.4285e-08 0.0013786 1.42865e-08 0 1.60835e-08 0 1.6085e-08 0.0013786 1.60865e-08 0 1.62835e-08 0 1.6285e-08 0.0013786 1.62865e-08 0 1.64835e-08 0 1.6485e-08 0.0013786 1.64865e-08 0 1.66835e-08 0 1.6685e-08 0.0013786 1.66865e-08 0 1.68835e-08 0 1.6885e-08 0.0013786 1.68865e-08 0 1.70835e-08 0 1.7085e-08 0.0013786 1.70865e-08 0 1.72835e-08 0 1.7285e-08 0.0013786 1.72865e-08 0 1.74835e-08 0 1.7485e-08 0.0013786 1.74865e-08 0 1.92835e-08 0 1.9285e-08 0.0013786 1.92865e-08 0 1.94835e-08 0 1.9485e-08 0.0013786 1.94865e-08 0 1.96835e-08 0 1.9685e-08 0.0013786 1.96865e-08 0 1.98835e-08 0 1.9885e-08 0.0013786 1.98865e-08 0 2.00835e-08 0 2.0085e-08 0.0013786 2.00865e-08 0 2.02835e-08 0 2.0285e-08 0.0013786 2.02865e-08 0 2.04835e-08 0 2.0485e-08 0.0013786 2.04865e-08 0 2.06835e-08 0 2.0685e-08 0.0013786 2.06865e-08 0 2.24835e-08 0 2.2485e-08 0.0013786 2.24865e-08 0 2.26835e-08 0 2.2685e-08 0.0013786 2.26865e-08 0 2.28835e-08 0 2.2885e-08 0.0013786 2.28865e-08 0 2.30835e-08 0 2.3085e-08 0.0013786 2.30865e-08 0 2.32835e-08 0 2.3285e-08 0.0013786 2.32865e-08 0 2.34835e-08 0 2.3485e-08 0.0013786 2.34865e-08 0 2.36835e-08 0 2.3685e-08 0.0013786 2.36865e-08 0 2.38835e-08 0 2.3885e-08 0.0013786 2.38865e-08 0 2.56835e-08 0 2.5685e-08 0.0013786 2.56865e-08 0 2.58835e-08 0 2.5885e-08 0.0013786 2.58865e-08 0 2.60835e-08 0 2.6085e-08 0.0013786 2.60865e-08 0 2.62835e-08 0 2.6285e-08 0.0013786 2.62865e-08 0 2.64835e-08 0 2.6485e-08 0.0013786 2.64865e-08 0 2.66835e-08 0 2.6685e-08 0.0013786 2.66865e-08 0 2.68835e-08 0 2.6885e-08 0.0013786 2.68865e-08 0 2.70835e-08 0 2.7085e-08 0.0013786 2.70865e-08 0 2.88835e-08 0 2.8885e-08 0.0013786 2.88865e-08 0 2.90835e-08 0 2.9085e-08 0.0013786 2.90865e-08 0 2.92835e-08 0 2.9285e-08 0.0013786 2.92865e-08 0 2.94835e-08 0 2.9485e-08 0.0013786 2.94865e-08 0 2.96835e-08 0 2.9685e-08 0.0013786 2.96865e-08 0 2.98835e-08 0 2.9885e-08 0.0013786 2.98865e-08 0 3.00835e-08 0 3.0085e-08 0.0013786 3.00865e-08 0 3.02835e-08 0 3.0285e-08 0.0013786 3.02865e-08 0 3.20835e-08 0 3.2085e-08 0.0013786 3.20865e-08 0 3.22835e-08 0 3.2285e-08 0.0013786 3.22865e-08 0 3.24835e-08 0 3.2485e-08 0.0013786 3.24865e-08 0 3.26835e-08 0 3.2685e-08 0.0013786 3.26865e-08 0 3.28835e-08 0 3.2885e-08 0.0013786 3.28865e-08 0 3.30835e-08 0 3.3085e-08 0.0013786 3.30865e-08 0 3.32835e-08 0 3.3285e-08 0.0013786 3.32865e-08 0 3.34835e-08 0 3.3485e-08 0.0013786 3.34865e-08 0 3.52835e-08 0 3.5285e-08 0.0013786 3.52865e-08 0 3.54835e-08 0 3.5485e-08 0.0013786 3.54865e-08 0 3.56835e-08 0 3.5685e-08 0.0013786 3.56865e-08 0 3.58835e-08 0 3.5885e-08 0.0013786 3.58865e-08 0 3.60835e-08 0 3.6085e-08 0.0013786 3.60865e-08 0 3.62835e-08 0 3.6285e-08 0.0013786 3.62865e-08 0 3.64835e-08 0 3.6485e-08 0.0013786 3.64865e-08 0 3.66835e-08 0 3.6685e-08 0.0013786 3.66865e-08 0 3.84835e-08 0 3.8485e-08 0.0013786 3.84865e-08 0 3.86835e-08 0 3.8685e-08 0.0013786 3.86865e-08 0 3.88835e-08 0 3.8885e-08 0.0013786 3.88865e-08 0 3.90835e-08 0 3.9085e-08 0.0013786 3.90865e-08 0 3.92835e-08 0 3.9285e-08 0.0013786 3.92865e-08 0 3.94835e-08 0 3.9485e-08 0.0013786 3.94865e-08 0 3.96835e-08 0 3.9685e-08 0.0013786 3.96865e-08 0 3.98835e-08 0 3.9885e-08 0.0013786 3.98865e-08 0 4.16835e-08 0 4.1685e-08 0.0013786 4.16865e-08 0 4.18835e-08 0 4.1885e-08 0.0013786 4.18865e-08 0 4.20835e-08 0 4.2085e-08 0.0013786 4.20865e-08 0 4.22835e-08 0 4.2285e-08 0.0013786 4.22865e-08 0 4.24835e-08 0 4.2485e-08 0.0013786 4.24865e-08 0 4.26835e-08 0 4.2685e-08 0.0013786 4.26865e-08 0 4.28835e-08 0 4.2885e-08 0.0013786 4.28865e-08 0 4.30835e-08 0 4.3085e-08 0.0013786 4.30865e-08 0 4.48835e-08 0 4.4885e-08 0.0013786 4.48865e-08 0 4.50835e-08 0 4.5085e-08 0.0013786 4.50865e-08 0 4.52835e-08 0 4.5285e-08 0.0013786 4.52865e-08 0 4.54835e-08 0 4.5485e-08 0.0013786 4.54865e-08 0 4.56835e-08 0 4.5685e-08 0.0013786 4.56865e-08 0 4.58835e-08 0 4.5885e-08 0.0013786 4.58865e-08 0 4.60835e-08 0 4.6085e-08 0.0013786 4.60865e-08 0 4.62835e-08 0 4.6285e-08 0.0013786 4.62865e-08 0 4.80835e-08 0 4.8085e-08 0.0013786 4.80865e-08 0 4.82835e-08 0 4.8285e-08 0.0013786 4.82865e-08 0 4.84835e-08 0 4.8485e-08 0.0013786 4.84865e-08 0 4.86835e-08 0 4.8685e-08 0.0013786 4.86865e-08 0 4.88835e-08 0 4.8885e-08 0.0013786 4.88865e-08 0 4.90835e-08 0 4.9085e-08 0.0013786 4.90865e-08 0 4.92835e-08 0 4.9285e-08 0.0013786 4.92865e-08 0 4.94835e-08 0 4.9485e-08 0.0013786 4.94865e-08 0)
IA2_|E 0 A2_  PWL(0 0 9.95e-11 0 1.01e-10 0.0013786 1.025e-10 0 2.995e-10 0 3.01e-10 0.0013786 3.025e-10 0 4.995e-10 0 5.01e-10 0.0013786 5.025e-10 0 6.995e-10 0 7.01e-10 0.0013786 7.025e-10 0 8.995e-10 0 9.01e-10 0.0013786 9.025e-10 0 1.0995e-09 0 1.101e-09 0.0013786 1.1025e-09 0 1.2995e-09 0 1.301e-09 0.0013786 1.3025e-09 0 1.4995e-09 0 1.501e-09 0.0013786 1.5025e-09 0 1.6995e-09 0 1.701e-09 0.0013786 1.7025e-09 0 1.8995e-09 0 1.901e-09 0.0013786 1.9025e-09 0 2.0995e-09 0 2.101e-09 0.0013786 2.1025e-09 0 2.2995e-09 0 2.301e-09 0.0013786 2.3025e-09 0 2.4995e-09 0 2.501e-09 0.0013786 2.5025e-09 0 2.6995e-09 0 2.701e-09 0.0013786 2.7025e-09 0 2.8995e-09 0 2.901e-09 0.0013786 2.9025e-09 0 3.0995e-09 0 3.101e-09 0.0013786 3.1025e-09 0 6.4995e-09 0 6.501e-09 0.0013786 6.5025e-09 0 6.6995e-09 0 6.701e-09 0.0013786 6.7025e-09 0 6.8995e-09 0 6.901e-09 0.0013786 6.9025e-09 0 7.0995e-09 0 7.101e-09 0.0013786 7.1025e-09 0 7.2995e-09 0 7.301e-09 0.0013786 7.3025e-09 0 7.4995e-09 0 7.501e-09 0.0013786 7.5025e-09 0 7.6995e-09 0 7.701e-09 0.0013786 7.7025e-09 0 7.8995e-09 0 7.901e-09 0.0013786 7.9025e-09 0 8.0995e-09 0 8.101e-09 0.0013786 8.1025e-09 0 8.2995e-09 0 8.301e-09 0.0013786 8.3025e-09 0 8.4995e-09 0 8.501e-09 0.0013786 8.5025e-09 0 8.6995e-09 0 8.701e-09 0.0013786 8.7025e-09 0 8.8995e-09 0 8.901e-09 0.0013786 8.9025e-09 0 9.0995e-09 0 9.101e-09 0.0013786 9.1025e-09 0 9.2995e-09 0 9.301e-09 0.0013786 9.3025e-09 0 9.4995e-09 0 9.501e-09 0.0013786 9.5025e-09 0 1.28995e-08 0 1.2901e-08 0.0013786 1.29025e-08 0 1.30995e-08 0 1.3101e-08 0.0013786 1.31025e-08 0 1.32995e-08 0 1.3301e-08 0.0013786 1.33025e-08 0 1.34995e-08 0 1.3501e-08 0.0013786 1.35025e-08 0 1.36995e-08 0 1.3701e-08 0.0013786 1.37025e-08 0 1.38995e-08 0 1.3901e-08 0.0013786 1.39025e-08 0 1.40995e-08 0 1.4101e-08 0.0013786 1.41025e-08 0 1.42995e-08 0 1.4301e-08 0.0013786 1.43025e-08 0 1.44995e-08 0 1.4501e-08 0.0013786 1.45025e-08 0 1.46995e-08 0 1.4701e-08 0.0013786 1.47025e-08 0 1.48995e-08 0 1.4901e-08 0.0013786 1.49025e-08 0 1.50995e-08 0 1.5101e-08 0.0013786 1.51025e-08 0 1.52995e-08 0 1.5301e-08 0.0013786 1.53025e-08 0 1.54995e-08 0 1.5501e-08 0.0013786 1.55025e-08 0 1.56995e-08 0 1.5701e-08 0.0013786 1.57025e-08 0 1.58995e-08 0 1.5901e-08 0.0013786 1.59025e-08 0 1.92995e-08 0 1.9301e-08 0.0013786 1.93025e-08 0 1.94995e-08 0 1.9501e-08 0.0013786 1.95025e-08 0 1.96995e-08 0 1.9701e-08 0.0013786 1.97025e-08 0 1.98995e-08 0 1.9901e-08 0.0013786 1.99025e-08 0 2.00995e-08 0 2.0101e-08 0.0013786 2.01025e-08 0 2.02995e-08 0 2.0301e-08 0.0013786 2.03025e-08 0 2.04995e-08 0 2.0501e-08 0.0013786 2.05025e-08 0 2.06995e-08 0 2.0701e-08 0.0013786 2.07025e-08 0 2.08995e-08 0 2.0901e-08 0.0013786 2.09025e-08 0 2.10995e-08 0 2.1101e-08 0.0013786 2.11025e-08 0 2.12995e-08 0 2.1301e-08 0.0013786 2.13025e-08 0 2.14995e-08 0 2.1501e-08 0.0013786 2.15025e-08 0 2.16995e-08 0 2.1701e-08 0.0013786 2.17025e-08 0 2.18995e-08 0 2.1901e-08 0.0013786 2.19025e-08 0 2.20995e-08 0 2.2101e-08 0.0013786 2.21025e-08 0 2.22995e-08 0 2.2301e-08 0.0013786 2.23025e-08 0 2.56995e-08 0 2.5701e-08 0.0013786 2.57025e-08 0 2.58995e-08 0 2.5901e-08 0.0013786 2.59025e-08 0 2.60995e-08 0 2.6101e-08 0.0013786 2.61025e-08 0 2.62995e-08 0 2.6301e-08 0.0013786 2.63025e-08 0 2.64995e-08 0 2.6501e-08 0.0013786 2.65025e-08 0 2.66995e-08 0 2.6701e-08 0.0013786 2.67025e-08 0 2.68995e-08 0 2.6901e-08 0.0013786 2.69025e-08 0 2.70995e-08 0 2.7101e-08 0.0013786 2.71025e-08 0 2.72995e-08 0 2.7301e-08 0.0013786 2.73025e-08 0 2.74995e-08 0 2.7501e-08 0.0013786 2.75025e-08 0 2.76995e-08 0 2.7701e-08 0.0013786 2.77025e-08 0 2.78995e-08 0 2.7901e-08 0.0013786 2.79025e-08 0 2.80995e-08 0 2.8101e-08 0.0013786 2.81025e-08 0 2.82995e-08 0 2.8301e-08 0.0013786 2.83025e-08 0 2.84995e-08 0 2.8501e-08 0.0013786 2.85025e-08 0 2.86995e-08 0 2.8701e-08 0.0013786 2.87025e-08 0 3.20995e-08 0 3.2101e-08 0.0013786 3.21025e-08 0 3.22995e-08 0 3.2301e-08 0.0013786 3.23025e-08 0 3.24995e-08 0 3.2501e-08 0.0013786 3.25025e-08 0 3.26995e-08 0 3.2701e-08 0.0013786 3.27025e-08 0 3.28995e-08 0 3.2901e-08 0.0013786 3.29025e-08 0 3.30995e-08 0 3.3101e-08 0.0013786 3.31025e-08 0 3.32995e-08 0 3.3301e-08 0.0013786 3.33025e-08 0 3.34995e-08 0 3.3501e-08 0.0013786 3.35025e-08 0 3.36995e-08 0 3.3701e-08 0.0013786 3.37025e-08 0 3.38995e-08 0 3.3901e-08 0.0013786 3.39025e-08 0 3.40995e-08 0 3.4101e-08 0.0013786 3.41025e-08 0 3.42995e-08 0 3.4301e-08 0.0013786 3.43025e-08 0 3.44995e-08 0 3.4501e-08 0.0013786 3.45025e-08 0 3.46995e-08 0 3.4701e-08 0.0013786 3.47025e-08 0 3.48995e-08 0 3.4901e-08 0.0013786 3.49025e-08 0 3.50995e-08 0 3.5101e-08 0.0013786 3.51025e-08 0 3.84995e-08 0 3.8501e-08 0.0013786 3.85025e-08 0 3.86995e-08 0 3.8701e-08 0.0013786 3.87025e-08 0 3.88995e-08 0 3.8901e-08 0.0013786 3.89025e-08 0 3.90995e-08 0 3.9101e-08 0.0013786 3.91025e-08 0 3.92995e-08 0 3.9301e-08 0.0013786 3.93025e-08 0 3.94995e-08 0 3.9501e-08 0.0013786 3.95025e-08 0 3.96995e-08 0 3.9701e-08 0.0013786 3.97025e-08 0 3.98995e-08 0 3.9901e-08 0.0013786 3.99025e-08 0 4.00995e-08 0 4.0101e-08 0.0013786 4.01025e-08 0 4.02995e-08 0 4.0301e-08 0.0013786 4.03025e-08 0 4.04995e-08 0 4.0501e-08 0.0013786 4.05025e-08 0 4.06995e-08 0 4.0701e-08 0.0013786 4.07025e-08 0 4.08995e-08 0 4.0901e-08 0.0013786 4.09025e-08 0 4.10995e-08 0 4.1101e-08 0.0013786 4.11025e-08 0 4.12995e-08 0 4.1301e-08 0.0013786 4.13025e-08 0 4.14995e-08 0 4.1501e-08 0.0013786 4.15025e-08 0 4.48995e-08 0 4.4901e-08 0.0013786 4.49025e-08 0 4.50995e-08 0 4.5101e-08 0.0013786 4.51025e-08 0 4.52995e-08 0 4.5301e-08 0.0013786 4.53025e-08 0 4.54995e-08 0 4.5501e-08 0.0013786 4.55025e-08 0 4.56995e-08 0 4.5701e-08 0.0013786 4.57025e-08 0 4.58995e-08 0 4.5901e-08 0.0013786 4.59025e-08 0 4.60995e-08 0 4.6101e-08 0.0013786 4.61025e-08 0 4.62995e-08 0 4.6301e-08 0.0013786 4.63025e-08 0 4.64995e-08 0 4.6501e-08 0.0013786 4.65025e-08 0 4.66995e-08 0 4.6701e-08 0.0013786 4.67025e-08 0 4.68995e-08 0 4.6901e-08 0.0013786 4.69025e-08 0 4.70995e-08 0 4.7101e-08 0.0013786 4.71025e-08 0 4.72995e-08 0 4.7301e-08 0.0013786 4.73025e-08 0 4.74995e-08 0 4.7501e-08 0.0013786 4.75025e-08 0 4.76995e-08 0 4.7701e-08 0.0013786 4.77025e-08 0 4.78995e-08 0 4.7901e-08 0.0013786 4.79025e-08 0)
IB2_|F 0 B2_  PWL(0 0 1.155e-10 0 1.17e-10 0.0013786 1.185e-10 0 3.155e-10 0 3.17e-10 0.0013786 3.185e-10 0 5.155e-10 0 5.17e-10 0.0013786 5.185e-10 0 7.155e-10 0 7.17e-10 0.0013786 7.185e-10 0 9.155e-10 0 9.17e-10 0.0013786 9.185e-10 0 1.1155e-09 0 1.117e-09 0.0013786 1.1185e-09 0 1.3155e-09 0 1.317e-09 0.0013786 1.3185e-09 0 1.5155e-09 0 1.517e-09 0.0013786 1.5185e-09 0 1.7155e-09 0 1.717e-09 0.0013786 1.7185e-09 0 1.9155e-09 0 1.917e-09 0.0013786 1.9185e-09 0 2.1155e-09 0 2.117e-09 0.0013786 2.1185e-09 0 2.3155e-09 0 2.317e-09 0.0013786 2.3185e-09 0 2.5155e-09 0 2.517e-09 0.0013786 2.5185e-09 0 2.7155e-09 0 2.717e-09 0.0013786 2.7185e-09 0 2.9155e-09 0 2.917e-09 0.0013786 2.9185e-09 0 3.1155e-09 0 3.117e-09 0.0013786 3.1185e-09 0 3.3155e-09 0 3.317e-09 0.0013786 3.3185e-09 0 3.5155e-09 0 3.517e-09 0.0013786 3.5185e-09 0 3.7155e-09 0 3.717e-09 0.0013786 3.7185e-09 0 3.9155e-09 0 3.917e-09 0.0013786 3.9185e-09 0 4.1155e-09 0 4.117e-09 0.0013786 4.1185e-09 0 4.3155e-09 0 4.317e-09 0.0013786 4.3185e-09 0 4.5155e-09 0 4.517e-09 0.0013786 4.5185e-09 0 4.7155e-09 0 4.717e-09 0.0013786 4.7185e-09 0 4.9155e-09 0 4.917e-09 0.0013786 4.9185e-09 0 5.1155e-09 0 5.117e-09 0.0013786 5.1185e-09 0 5.3155e-09 0 5.317e-09 0.0013786 5.3185e-09 0 5.5155e-09 0 5.517e-09 0.0013786 5.5185e-09 0 5.7155e-09 0 5.717e-09 0.0013786 5.7185e-09 0 5.9155e-09 0 5.917e-09 0.0013786 5.9185e-09 0 6.1155e-09 0 6.117e-09 0.0013786 6.1185e-09 0 6.3155e-09 0 6.317e-09 0.0013786 6.3185e-09 0 1.29155e-08 0 1.2917e-08 0.0013786 1.29185e-08 0 1.31155e-08 0 1.3117e-08 0.0013786 1.31185e-08 0 1.33155e-08 0 1.3317e-08 0.0013786 1.33185e-08 0 1.35155e-08 0 1.3517e-08 0.0013786 1.35185e-08 0 1.37155e-08 0 1.3717e-08 0.0013786 1.37185e-08 0 1.39155e-08 0 1.3917e-08 0.0013786 1.39185e-08 0 1.41155e-08 0 1.4117e-08 0.0013786 1.41185e-08 0 1.43155e-08 0 1.4317e-08 0.0013786 1.43185e-08 0 1.45155e-08 0 1.4517e-08 0.0013786 1.45185e-08 0 1.47155e-08 0 1.4717e-08 0.0013786 1.47185e-08 0 1.49155e-08 0 1.4917e-08 0.0013786 1.49185e-08 0 1.51155e-08 0 1.5117e-08 0.0013786 1.51185e-08 0 1.53155e-08 0 1.5317e-08 0.0013786 1.53185e-08 0 1.55155e-08 0 1.5517e-08 0.0013786 1.55185e-08 0 1.57155e-08 0 1.5717e-08 0.0013786 1.57185e-08 0 1.59155e-08 0 1.5917e-08 0.0013786 1.59185e-08 0 1.61155e-08 0 1.6117e-08 0.0013786 1.61185e-08 0 1.63155e-08 0 1.6317e-08 0.0013786 1.63185e-08 0 1.65155e-08 0 1.6517e-08 0.0013786 1.65185e-08 0 1.67155e-08 0 1.6717e-08 0.0013786 1.67185e-08 0 1.69155e-08 0 1.6917e-08 0.0013786 1.69185e-08 0 1.71155e-08 0 1.7117e-08 0.0013786 1.71185e-08 0 1.73155e-08 0 1.7317e-08 0.0013786 1.73185e-08 0 1.75155e-08 0 1.7517e-08 0.0013786 1.75185e-08 0 1.77155e-08 0 1.7717e-08 0.0013786 1.77185e-08 0 1.79155e-08 0 1.7917e-08 0.0013786 1.79185e-08 0 1.81155e-08 0 1.8117e-08 0.0013786 1.81185e-08 0 1.83155e-08 0 1.8317e-08 0.0013786 1.83185e-08 0 1.85155e-08 0 1.8517e-08 0.0013786 1.85185e-08 0 1.87155e-08 0 1.8717e-08 0.0013786 1.87185e-08 0 1.89155e-08 0 1.8917e-08 0.0013786 1.89185e-08 0 1.91155e-08 0 1.9117e-08 0.0013786 1.91185e-08 0 2.57155e-08 0 2.5717e-08 0.0013786 2.57185e-08 0 2.59155e-08 0 2.5917e-08 0.0013786 2.59185e-08 0 2.61155e-08 0 2.6117e-08 0.0013786 2.61185e-08 0 2.63155e-08 0 2.6317e-08 0.0013786 2.63185e-08 0 2.65155e-08 0 2.6517e-08 0.0013786 2.65185e-08 0 2.67155e-08 0 2.6717e-08 0.0013786 2.67185e-08 0 2.69155e-08 0 2.6917e-08 0.0013786 2.69185e-08 0 2.71155e-08 0 2.7117e-08 0.0013786 2.71185e-08 0 2.73155e-08 0 2.7317e-08 0.0013786 2.73185e-08 0 2.75155e-08 0 2.7517e-08 0.0013786 2.75185e-08 0 2.77155e-08 0 2.7717e-08 0.0013786 2.77185e-08 0 2.79155e-08 0 2.7917e-08 0.0013786 2.79185e-08 0 2.81155e-08 0 2.8117e-08 0.0013786 2.81185e-08 0 2.83155e-08 0 2.8317e-08 0.0013786 2.83185e-08 0 2.85155e-08 0 2.8517e-08 0.0013786 2.85185e-08 0 2.87155e-08 0 2.8717e-08 0.0013786 2.87185e-08 0 2.89155e-08 0 2.8917e-08 0.0013786 2.89185e-08 0 2.91155e-08 0 2.9117e-08 0.0013786 2.91185e-08 0 2.93155e-08 0 2.9317e-08 0.0013786 2.93185e-08 0 2.95155e-08 0 2.9517e-08 0.0013786 2.95185e-08 0 2.97155e-08 0 2.9717e-08 0.0013786 2.97185e-08 0 2.99155e-08 0 2.9917e-08 0.0013786 2.99185e-08 0 3.01155e-08 0 3.0117e-08 0.0013786 3.01185e-08 0 3.03155e-08 0 3.0317e-08 0.0013786 3.03185e-08 0 3.05155e-08 0 3.0517e-08 0.0013786 3.05185e-08 0 3.07155e-08 0 3.0717e-08 0.0013786 3.07185e-08 0 3.09155e-08 0 3.0917e-08 0.0013786 3.09185e-08 0 3.11155e-08 0 3.1117e-08 0.0013786 3.11185e-08 0 3.13155e-08 0 3.1317e-08 0.0013786 3.13185e-08 0 3.15155e-08 0 3.1517e-08 0.0013786 3.15185e-08 0 3.17155e-08 0 3.1717e-08 0.0013786 3.17185e-08 0 3.19155e-08 0 3.1917e-08 0.0013786 3.19185e-08 0 3.85155e-08 0 3.8517e-08 0.0013786 3.85185e-08 0 3.87155e-08 0 3.8717e-08 0.0013786 3.87185e-08 0 3.89155e-08 0 3.8917e-08 0.0013786 3.89185e-08 0 3.91155e-08 0 3.9117e-08 0.0013786 3.91185e-08 0 3.93155e-08 0 3.9317e-08 0.0013786 3.93185e-08 0 3.95155e-08 0 3.9517e-08 0.0013786 3.95185e-08 0 3.97155e-08 0 3.9717e-08 0.0013786 3.97185e-08 0 3.99155e-08 0 3.9917e-08 0.0013786 3.99185e-08 0 4.01155e-08 0 4.0117e-08 0.0013786 4.01185e-08 0 4.03155e-08 0 4.0317e-08 0.0013786 4.03185e-08 0 4.05155e-08 0 4.0517e-08 0.0013786 4.05185e-08 0 4.07155e-08 0 4.0717e-08 0.0013786 4.07185e-08 0 4.09155e-08 0 4.0917e-08 0.0013786 4.09185e-08 0 4.11155e-08 0 4.1117e-08 0.0013786 4.11185e-08 0 4.13155e-08 0 4.1317e-08 0.0013786 4.13185e-08 0 4.15155e-08 0 4.1517e-08 0.0013786 4.15185e-08 0 4.17155e-08 0 4.1717e-08 0.0013786 4.17185e-08 0 4.19155e-08 0 4.1917e-08 0.0013786 4.19185e-08 0 4.21155e-08 0 4.2117e-08 0.0013786 4.21185e-08 0 4.23155e-08 0 4.2317e-08 0.0013786 4.23185e-08 0 4.25155e-08 0 4.2517e-08 0.0013786 4.25185e-08 0 4.27155e-08 0 4.2717e-08 0.0013786 4.27185e-08 0 4.29155e-08 0 4.2917e-08 0.0013786 4.29185e-08 0 4.31155e-08 0 4.3117e-08 0.0013786 4.31185e-08 0 4.33155e-08 0 4.3317e-08 0.0013786 4.33185e-08 0 4.35155e-08 0 4.3517e-08 0.0013786 4.35185e-08 0 4.37155e-08 0 4.3717e-08 0.0013786 4.37185e-08 0 4.39155e-08 0 4.3917e-08 0.0013786 4.39185e-08 0 4.41155e-08 0 4.4117e-08 0.0013786 4.41185e-08 0 4.43155e-08 0 4.4317e-08 0.0013786 4.43185e-08 0 4.45155e-08 0 4.4517e-08 0.0013786 4.45185e-08 0 4.47155e-08 0 4.4717e-08 0.0013786 4.47185e-08 0)
IA3_|G 0 A3_  PWL(0 0 1.315e-10 0 1.33e-10 0.0013786 1.345e-10 0 3.315e-10 0 3.33e-10 0.0013786 3.345e-10 0 5.315e-10 0 5.33e-10 0.0013786 5.345e-10 0 7.315e-10 0 7.33e-10 0.0013786 7.345e-10 0 9.315e-10 0 9.33e-10 0.0013786 9.345e-10 0 1.1315e-09 0 1.133e-09 0.0013786 1.1345e-09 0 1.3315e-09 0 1.333e-09 0.0013786 1.3345e-09 0 1.5315e-09 0 1.533e-09 0.0013786 1.5345e-09 0 1.7315e-09 0 1.733e-09 0.0013786 1.7345e-09 0 1.9315e-09 0 1.933e-09 0.0013786 1.9345e-09 0 2.1315e-09 0 2.133e-09 0.0013786 2.1345e-09 0 2.3315e-09 0 2.333e-09 0.0013786 2.3345e-09 0 2.5315e-09 0 2.533e-09 0.0013786 2.5345e-09 0 2.7315e-09 0 2.733e-09 0.0013786 2.7345e-09 0 2.9315e-09 0 2.933e-09 0.0013786 2.9345e-09 0 3.1315e-09 0 3.133e-09 0.0013786 3.1345e-09 0 3.3315e-09 0 3.333e-09 0.0013786 3.3345e-09 0 3.5315e-09 0 3.533e-09 0.0013786 3.5345e-09 0 3.7315e-09 0 3.733e-09 0.0013786 3.7345e-09 0 3.9315e-09 0 3.933e-09 0.0013786 3.9345e-09 0 4.1315e-09 0 4.133e-09 0.0013786 4.1345e-09 0 4.3315e-09 0 4.333e-09 0.0013786 4.3345e-09 0 4.5315e-09 0 4.533e-09 0.0013786 4.5345e-09 0 4.7315e-09 0 4.733e-09 0.0013786 4.7345e-09 0 4.9315e-09 0 4.933e-09 0.0013786 4.9345e-09 0 5.1315e-09 0 5.133e-09 0.0013786 5.1345e-09 0 5.3315e-09 0 5.333e-09 0.0013786 5.3345e-09 0 5.5315e-09 0 5.533e-09 0.0013786 5.5345e-09 0 5.7315e-09 0 5.733e-09 0.0013786 5.7345e-09 0 5.9315e-09 0 5.933e-09 0.0013786 5.9345e-09 0 6.1315e-09 0 6.133e-09 0.0013786 6.1345e-09 0 6.3315e-09 0 6.333e-09 0.0013786 6.3345e-09 0 6.5315e-09 0 6.533e-09 0.0013786 6.5345e-09 0 6.7315e-09 0 6.733e-09 0.0013786 6.7345e-09 0 6.9315e-09 0 6.933e-09 0.0013786 6.9345e-09 0 7.1315e-09 0 7.133e-09 0.0013786 7.1345e-09 0 7.3315e-09 0 7.333e-09 0.0013786 7.3345e-09 0 7.5315e-09 0 7.533e-09 0.0013786 7.5345e-09 0 7.7315e-09 0 7.733e-09 0.0013786 7.7345e-09 0 7.9315e-09 0 7.933e-09 0.0013786 7.9345e-09 0 8.1315e-09 0 8.133e-09 0.0013786 8.1345e-09 0 8.3315e-09 0 8.333e-09 0.0013786 8.3345e-09 0 8.5315e-09 0 8.533e-09 0.0013786 8.5345e-09 0 8.7315e-09 0 8.733e-09 0.0013786 8.7345e-09 0 8.9315e-09 0 8.933e-09 0.0013786 8.9345e-09 0 9.1315e-09 0 9.133e-09 0.0013786 9.1345e-09 0 9.3315e-09 0 9.333e-09 0.0013786 9.3345e-09 0 9.5315e-09 0 9.533e-09 0.0013786 9.5345e-09 0 9.7315e-09 0 9.733e-09 0.0013786 9.7345e-09 0 9.9315e-09 0 9.933e-09 0.0013786 9.9345e-09 0 1.01315e-08 0 1.0133e-08 0.0013786 1.01345e-08 0 1.03315e-08 0 1.0333e-08 0.0013786 1.03345e-08 0 1.05315e-08 0 1.0533e-08 0.0013786 1.05345e-08 0 1.07315e-08 0 1.0733e-08 0.0013786 1.07345e-08 0 1.09315e-08 0 1.0933e-08 0.0013786 1.09345e-08 0 1.11315e-08 0 1.1133e-08 0.0013786 1.11345e-08 0 1.13315e-08 0 1.1333e-08 0.0013786 1.13345e-08 0 1.15315e-08 0 1.1533e-08 0.0013786 1.15345e-08 0 1.17315e-08 0 1.1733e-08 0.0013786 1.17345e-08 0 1.19315e-08 0 1.1933e-08 0.0013786 1.19345e-08 0 1.21315e-08 0 1.2133e-08 0.0013786 1.21345e-08 0 1.23315e-08 0 1.2333e-08 0.0013786 1.23345e-08 0 1.25315e-08 0 1.2533e-08 0.0013786 1.25345e-08 0 1.27315e-08 0 1.2733e-08 0.0013786 1.27345e-08 0 2.57315e-08 0 2.5733e-08 0.0013786 2.57345e-08 0 2.59315e-08 0 2.5933e-08 0.0013786 2.59345e-08 0 2.61315e-08 0 2.6133e-08 0.0013786 2.61345e-08 0 2.63315e-08 0 2.6333e-08 0.0013786 2.63345e-08 0 2.65315e-08 0 2.6533e-08 0.0013786 2.65345e-08 0 2.67315e-08 0 2.6733e-08 0.0013786 2.67345e-08 0 2.69315e-08 0 2.6933e-08 0.0013786 2.69345e-08 0 2.71315e-08 0 2.7133e-08 0.0013786 2.71345e-08 0 2.73315e-08 0 2.7333e-08 0.0013786 2.73345e-08 0 2.75315e-08 0 2.7533e-08 0.0013786 2.75345e-08 0 2.77315e-08 0 2.7733e-08 0.0013786 2.77345e-08 0 2.79315e-08 0 2.7933e-08 0.0013786 2.79345e-08 0 2.81315e-08 0 2.8133e-08 0.0013786 2.81345e-08 0 2.83315e-08 0 2.8333e-08 0.0013786 2.83345e-08 0 2.85315e-08 0 2.8533e-08 0.0013786 2.85345e-08 0 2.87315e-08 0 2.8733e-08 0.0013786 2.87345e-08 0 2.89315e-08 0 2.8933e-08 0.0013786 2.89345e-08 0 2.91315e-08 0 2.9133e-08 0.0013786 2.91345e-08 0 2.93315e-08 0 2.9333e-08 0.0013786 2.93345e-08 0 2.95315e-08 0 2.9533e-08 0.0013786 2.95345e-08 0 2.97315e-08 0 2.9733e-08 0.0013786 2.97345e-08 0 2.99315e-08 0 2.9933e-08 0.0013786 2.99345e-08 0 3.01315e-08 0 3.0133e-08 0.0013786 3.01345e-08 0 3.03315e-08 0 3.0333e-08 0.0013786 3.03345e-08 0 3.05315e-08 0 3.0533e-08 0.0013786 3.05345e-08 0 3.07315e-08 0 3.0733e-08 0.0013786 3.07345e-08 0 3.09315e-08 0 3.0933e-08 0.0013786 3.09345e-08 0 3.11315e-08 0 3.1133e-08 0.0013786 3.11345e-08 0 3.13315e-08 0 3.1333e-08 0.0013786 3.13345e-08 0 3.15315e-08 0 3.1533e-08 0.0013786 3.15345e-08 0 3.17315e-08 0 3.1733e-08 0.0013786 3.17345e-08 0 3.19315e-08 0 3.1933e-08 0.0013786 3.19345e-08 0 3.21315e-08 0 3.2133e-08 0.0013786 3.21345e-08 0 3.23315e-08 0 3.2333e-08 0.0013786 3.23345e-08 0 3.25315e-08 0 3.2533e-08 0.0013786 3.25345e-08 0 3.27315e-08 0 3.2733e-08 0.0013786 3.27345e-08 0 3.29315e-08 0 3.2933e-08 0.0013786 3.29345e-08 0 3.31315e-08 0 3.3133e-08 0.0013786 3.31345e-08 0 3.33315e-08 0 3.3333e-08 0.0013786 3.33345e-08 0 3.35315e-08 0 3.3533e-08 0.0013786 3.35345e-08 0 3.37315e-08 0 3.3733e-08 0.0013786 3.37345e-08 0 3.39315e-08 0 3.3933e-08 0.0013786 3.39345e-08 0 3.41315e-08 0 3.4133e-08 0.0013786 3.41345e-08 0 3.43315e-08 0 3.4333e-08 0.0013786 3.43345e-08 0 3.45315e-08 0 3.4533e-08 0.0013786 3.45345e-08 0 3.47315e-08 0 3.4733e-08 0.0013786 3.47345e-08 0 3.49315e-08 0 3.4933e-08 0.0013786 3.49345e-08 0 3.51315e-08 0 3.5133e-08 0.0013786 3.51345e-08 0 3.53315e-08 0 3.5333e-08 0.0013786 3.53345e-08 0 3.55315e-08 0 3.5533e-08 0.0013786 3.55345e-08 0 3.57315e-08 0 3.5733e-08 0.0013786 3.57345e-08 0 3.59315e-08 0 3.5933e-08 0.0013786 3.59345e-08 0 3.61315e-08 0 3.6133e-08 0.0013786 3.61345e-08 0 3.63315e-08 0 3.6333e-08 0.0013786 3.63345e-08 0 3.65315e-08 0 3.6533e-08 0.0013786 3.65345e-08 0 3.67315e-08 0 3.6733e-08 0.0013786 3.67345e-08 0 3.69315e-08 0 3.6933e-08 0.0013786 3.69345e-08 0 3.71315e-08 0 3.7133e-08 0.0013786 3.71345e-08 0 3.73315e-08 0 3.7333e-08 0.0013786 3.73345e-08 0 3.75315e-08 0 3.7533e-08 0.0013786 3.75345e-08 0 3.77315e-08 0 3.7733e-08 0.0013786 3.77345e-08 0 3.79315e-08 0 3.7933e-08 0.0013786 3.79345e-08 0 3.81315e-08 0 3.8133e-08 0.0013786 3.81345e-08 0 3.83315e-08 0 3.8333e-08 0.0013786 3.83345e-08 0)
IB3_|H 0 B3_  PWL(0 0 1.475e-10 0 1.49e-10 0.0013786 1.505e-10 0 3.475e-10 0 3.49e-10 0.0013786 3.505e-10 0 5.475e-10 0 5.49e-10 0.0013786 5.505e-10 0 7.475e-10 0 7.49e-10 0.0013786 7.505e-10 0 9.475e-10 0 9.49e-10 0.0013786 9.505e-10 0 1.1475e-09 0 1.149e-09 0.0013786 1.1505e-09 0 1.3475e-09 0 1.349e-09 0.0013786 1.3505e-09 0 1.5475e-09 0 1.549e-09 0.0013786 1.5505e-09 0 1.7475e-09 0 1.749e-09 0.0013786 1.7505e-09 0 1.9475e-09 0 1.949e-09 0.0013786 1.9505e-09 0 2.1475e-09 0 2.149e-09 0.0013786 2.1505e-09 0 2.3475e-09 0 2.349e-09 0.0013786 2.3505e-09 0 2.5475e-09 0 2.549e-09 0.0013786 2.5505e-09 0 2.7475e-09 0 2.749e-09 0.0013786 2.7505e-09 0 2.9475e-09 0 2.949e-09 0.0013786 2.9505e-09 0 3.1475e-09 0 3.149e-09 0.0013786 3.1505e-09 0 3.3475e-09 0 3.349e-09 0.0013786 3.3505e-09 0 3.5475e-09 0 3.549e-09 0.0013786 3.5505e-09 0 3.7475e-09 0 3.749e-09 0.0013786 3.7505e-09 0 3.9475e-09 0 3.949e-09 0.0013786 3.9505e-09 0 4.1475e-09 0 4.149e-09 0.0013786 4.1505e-09 0 4.3475e-09 0 4.349e-09 0.0013786 4.3505e-09 0 4.5475e-09 0 4.549e-09 0.0013786 4.5505e-09 0 4.7475e-09 0 4.749e-09 0.0013786 4.7505e-09 0 4.9475e-09 0 4.949e-09 0.0013786 4.9505e-09 0 5.1475e-09 0 5.149e-09 0.0013786 5.1505e-09 0 5.3475e-09 0 5.349e-09 0.0013786 5.3505e-09 0 5.5475e-09 0 5.549e-09 0.0013786 5.5505e-09 0 5.7475e-09 0 5.749e-09 0.0013786 5.7505e-09 0 5.9475e-09 0 5.949e-09 0.0013786 5.9505e-09 0 6.1475e-09 0 6.149e-09 0.0013786 6.1505e-09 0 6.3475e-09 0 6.349e-09 0.0013786 6.3505e-09 0 6.5475e-09 0 6.549e-09 0.0013786 6.5505e-09 0 6.7475e-09 0 6.749e-09 0.0013786 6.7505e-09 0 6.9475e-09 0 6.949e-09 0.0013786 6.9505e-09 0 7.1475e-09 0 7.149e-09 0.0013786 7.1505e-09 0 7.3475e-09 0 7.349e-09 0.0013786 7.3505e-09 0 7.5475e-09 0 7.549e-09 0.0013786 7.5505e-09 0 7.7475e-09 0 7.749e-09 0.0013786 7.7505e-09 0 7.9475e-09 0 7.949e-09 0.0013786 7.9505e-09 0 8.1475e-09 0 8.149e-09 0.0013786 8.1505e-09 0 8.3475e-09 0 8.349e-09 0.0013786 8.3505e-09 0 8.5475e-09 0 8.549e-09 0.0013786 8.5505e-09 0 8.7475e-09 0 8.749e-09 0.0013786 8.7505e-09 0 8.9475e-09 0 8.949e-09 0.0013786 8.9505e-09 0 9.1475e-09 0 9.149e-09 0.0013786 9.1505e-09 0 9.3475e-09 0 9.349e-09 0.0013786 9.3505e-09 0 9.5475e-09 0 9.549e-09 0.0013786 9.5505e-09 0 9.7475e-09 0 9.749e-09 0.0013786 9.7505e-09 0 9.9475e-09 0 9.949e-09 0.0013786 9.9505e-09 0 1.01475e-08 0 1.0149e-08 0.0013786 1.01505e-08 0 1.03475e-08 0 1.0349e-08 0.0013786 1.03505e-08 0 1.05475e-08 0 1.0549e-08 0.0013786 1.05505e-08 0 1.07475e-08 0 1.0749e-08 0.0013786 1.07505e-08 0 1.09475e-08 0 1.0949e-08 0.0013786 1.09505e-08 0 1.11475e-08 0 1.1149e-08 0.0013786 1.11505e-08 0 1.13475e-08 0 1.1349e-08 0.0013786 1.13505e-08 0 1.15475e-08 0 1.1549e-08 0.0013786 1.15505e-08 0 1.17475e-08 0 1.1749e-08 0.0013786 1.17505e-08 0 1.19475e-08 0 1.1949e-08 0.0013786 1.19505e-08 0 1.21475e-08 0 1.2149e-08 0.0013786 1.21505e-08 0 1.23475e-08 0 1.2349e-08 0.0013786 1.23505e-08 0 1.25475e-08 0 1.2549e-08 0.0013786 1.25505e-08 0 1.27475e-08 0 1.2749e-08 0.0013786 1.27505e-08 0 1.29475e-08 0 1.2949e-08 0.0013786 1.29505e-08 0 1.31475e-08 0 1.3149e-08 0.0013786 1.31505e-08 0 1.33475e-08 0 1.3349e-08 0.0013786 1.33505e-08 0 1.35475e-08 0 1.3549e-08 0.0013786 1.35505e-08 0 1.37475e-08 0 1.3749e-08 0.0013786 1.37505e-08 0 1.39475e-08 0 1.3949e-08 0.0013786 1.39505e-08 0 1.41475e-08 0 1.4149e-08 0.0013786 1.41505e-08 0 1.43475e-08 0 1.4349e-08 0.0013786 1.43505e-08 0 1.45475e-08 0 1.4549e-08 0.0013786 1.45505e-08 0 1.47475e-08 0 1.4749e-08 0.0013786 1.47505e-08 0 1.49475e-08 0 1.4949e-08 0.0013786 1.49505e-08 0 1.51475e-08 0 1.5149e-08 0.0013786 1.51505e-08 0 1.53475e-08 0 1.5349e-08 0.0013786 1.53505e-08 0 1.55475e-08 0 1.5549e-08 0.0013786 1.55505e-08 0 1.57475e-08 0 1.5749e-08 0.0013786 1.57505e-08 0 1.59475e-08 0 1.5949e-08 0.0013786 1.59505e-08 0 1.61475e-08 0 1.6149e-08 0.0013786 1.61505e-08 0 1.63475e-08 0 1.6349e-08 0.0013786 1.63505e-08 0 1.65475e-08 0 1.6549e-08 0.0013786 1.65505e-08 0 1.67475e-08 0 1.6749e-08 0.0013786 1.67505e-08 0 1.69475e-08 0 1.6949e-08 0.0013786 1.69505e-08 0 1.71475e-08 0 1.7149e-08 0.0013786 1.71505e-08 0 1.73475e-08 0 1.7349e-08 0.0013786 1.73505e-08 0 1.75475e-08 0 1.7549e-08 0.0013786 1.75505e-08 0 1.77475e-08 0 1.7749e-08 0.0013786 1.77505e-08 0 1.79475e-08 0 1.7949e-08 0.0013786 1.79505e-08 0 1.81475e-08 0 1.8149e-08 0.0013786 1.81505e-08 0 1.83475e-08 0 1.8349e-08 0.0013786 1.83505e-08 0 1.85475e-08 0 1.8549e-08 0.0013786 1.85505e-08 0 1.87475e-08 0 1.8749e-08 0.0013786 1.87505e-08 0 1.89475e-08 0 1.8949e-08 0.0013786 1.89505e-08 0 1.91475e-08 0 1.9149e-08 0.0013786 1.91505e-08 0 1.93475e-08 0 1.9349e-08 0.0013786 1.93505e-08 0 1.95475e-08 0 1.9549e-08 0.0013786 1.95505e-08 0 1.97475e-08 0 1.9749e-08 0.0013786 1.97505e-08 0 1.99475e-08 0 1.9949e-08 0.0013786 1.99505e-08 0 2.01475e-08 0 2.0149e-08 0.0013786 2.01505e-08 0 2.03475e-08 0 2.0349e-08 0.0013786 2.03505e-08 0 2.05475e-08 0 2.0549e-08 0.0013786 2.05505e-08 0 2.07475e-08 0 2.0749e-08 0.0013786 2.07505e-08 0 2.09475e-08 0 2.0949e-08 0.0013786 2.09505e-08 0 2.11475e-08 0 2.1149e-08 0.0013786 2.11505e-08 0 2.13475e-08 0 2.1349e-08 0.0013786 2.13505e-08 0 2.15475e-08 0 2.1549e-08 0.0013786 2.15505e-08 0 2.17475e-08 0 2.1749e-08 0.0013786 2.17505e-08 0 2.19475e-08 0 2.1949e-08 0.0013786 2.19505e-08 0 2.21475e-08 0 2.2149e-08 0.0013786 2.21505e-08 0 2.23475e-08 0 2.2349e-08 0.0013786 2.23505e-08 0 2.25475e-08 0 2.2549e-08 0.0013786 2.25505e-08 0 2.27475e-08 0 2.2749e-08 0.0013786 2.27505e-08 0 2.29475e-08 0 2.2949e-08 0.0013786 2.29505e-08 0 2.31475e-08 0 2.3149e-08 0.0013786 2.31505e-08 0 2.33475e-08 0 2.3349e-08 0.0013786 2.33505e-08 0 2.35475e-08 0 2.3549e-08 0.0013786 2.35505e-08 0 2.37475e-08 0 2.3749e-08 0.0013786 2.37505e-08 0 2.39475e-08 0 2.3949e-08 0.0013786 2.39505e-08 0 2.41475e-08 0 2.4149e-08 0.0013786 2.41505e-08 0 2.43475e-08 0 2.4349e-08 0.0013786 2.43505e-08 0 2.45475e-08 0 2.4549e-08 0.0013786 2.45505e-08 0 2.47475e-08 0 2.4749e-08 0.0013786 2.47505e-08 0 2.49475e-08 0 2.4949e-08 0.0013786 2.49505e-08 0 2.51475e-08 0 2.5149e-08 0.0013786 2.51505e-08 0 2.53475e-08 0 2.5349e-08 0.0013786 2.53505e-08 0 2.55475e-08 0 2.5549e-08 0.0013786 2.55505e-08 0)
IT00_|T 0 T00_  PWL(0 0 1.85e-11 0 2e-11 0.0041358 2.15e-11 0 2.185e-10 0 2.2e-10 0.0041358 2.215e-10 0 4.185e-10 0 4.2e-10 0.0041358 4.215e-10 0 6.185e-10 0 6.2e-10 0.0041358 6.215e-10 0 8.185e-10 0 8.2e-10 0.0041358 8.215e-10 0 1.0185e-09 0 1.02e-09 0.0041358 1.0215e-09 0 1.2185e-09 0 1.22e-09 0.0041358 1.2215e-09 0 1.4185e-09 0 1.42e-09 0.0041358 1.4215e-09 0 1.6185e-09 0 1.62e-09 0.0041358 1.6215e-09 0 1.8185e-09 0 1.82e-09 0.0041358 1.8215e-09 0 2.0185e-09 0 2.02e-09 0.0041358 2.0215e-09 0 2.2185e-09 0 2.22e-09 0.0041358 2.2215e-09 0 2.4185e-09 0 2.42e-09 0.0041358 2.4215e-09 0 2.6185e-09 0 2.62e-09 0.0041358 2.6215e-09 0 2.8185e-09 0 2.82e-09 0.0041358 2.8215e-09 0 3.0185e-09 0 3.02e-09 0.0041358 3.0215e-09 0 3.2185e-09 0 3.22e-09 0.0041358 3.2215e-09 0 3.4185e-09 0 3.42e-09 0.0041358 3.4215e-09 0 3.6185e-09 0 3.62e-09 0.0041358 3.6215e-09 0 3.8185e-09 0 3.82e-09 0.0041358 3.8215e-09 0 4.0185e-09 0 4.02e-09 0.0041358 4.0215e-09 0 4.2185e-09 0 4.22e-09 0.0041358 4.2215e-09 0 4.4185e-09 0 4.42e-09 0.0041358 4.4215e-09 0 4.6185e-09 0 4.62e-09 0.0041358 4.6215e-09 0 4.8185e-09 0 4.82e-09 0.0041358 4.8215e-09 0 5.0185e-09 0 5.02e-09 0.0041358 5.0215e-09 0 5.2185e-09 0 5.22e-09 0.0041358 5.2215e-09 0 5.4185e-09 0 5.42e-09 0.0041358 5.4215e-09 0 5.6185e-09 0 5.62e-09 0.0041358 5.6215e-09 0 5.8185e-09 0 5.82e-09 0.0041358 5.8215e-09 0 6.0185e-09 0 6.02e-09 0.0041358 6.0215e-09 0 6.2185e-09 0 6.22e-09 0.0041358 6.2215e-09 0 6.4185e-09 0 6.42e-09 0.0041358 6.4215e-09 0 6.6185e-09 0 6.62e-09 0.0041358 6.6215e-09 0 6.8185e-09 0 6.82e-09 0.0041358 6.8215e-09 0 7.0185e-09 0 7.02e-09 0.0041358 7.0215e-09 0 7.2185e-09 0 7.22e-09 0.0041358 7.2215e-09 0 7.4185e-09 0 7.42e-09 0.0041358 7.4215e-09 0 7.6185e-09 0 7.62e-09 0.0041358 7.6215e-09 0 7.8185e-09 0 7.82e-09 0.0041358 7.8215e-09 0 8.0185e-09 0 8.02e-09 0.0041358 8.0215e-09 0 8.2185e-09 0 8.22e-09 0.0041358 8.2215e-09 0 8.4185e-09 0 8.42e-09 0.0041358 8.4215e-09 0 8.6185e-09 0 8.62e-09 0.0041358 8.6215e-09 0 8.8185e-09 0 8.82e-09 0.0041358 8.8215e-09 0 9.0185e-09 0 9.02e-09 0.0041358 9.0215e-09 0 9.2185e-09 0 9.22e-09 0.0041358 9.2215e-09 0 9.4185e-09 0 9.42e-09 0.0041358 9.4215e-09 0 9.6185e-09 0 9.62e-09 0.0041358 9.6215e-09 0 9.8185e-09 0 9.82e-09 0.0041358 9.8215e-09 0 1.00185e-08 0 1.002e-08 0.0041358 1.00215e-08 0 1.02185e-08 0 1.022e-08 0.0041358 1.02215e-08 0 1.04185e-08 0 1.042e-08 0.0041358 1.04215e-08 0 1.06185e-08 0 1.062e-08 0.0041358 1.06215e-08 0 1.08185e-08 0 1.082e-08 0.0041358 1.08215e-08 0 1.10185e-08 0 1.102e-08 0.0041358 1.10215e-08 0 1.12185e-08 0 1.122e-08 0.0041358 1.12215e-08 0 1.14185e-08 0 1.142e-08 0.0041358 1.14215e-08 0 1.16185e-08 0 1.162e-08 0.0041358 1.16215e-08 0 1.18185e-08 0 1.182e-08 0.0041358 1.18215e-08 0 1.20185e-08 0 1.202e-08 0.0041358 1.20215e-08 0 1.22185e-08 0 1.222e-08 0.0041358 1.22215e-08 0 1.24185e-08 0 1.242e-08 0.0041358 1.24215e-08 0 1.26185e-08 0 1.262e-08 0.0041358 1.26215e-08 0 1.28185e-08 0 1.282e-08 0.0041358 1.28215e-08 0 1.30185e-08 0 1.302e-08 0.0041358 1.30215e-08 0 1.32185e-08 0 1.322e-08 0.0041358 1.32215e-08 0 1.34185e-08 0 1.342e-08 0.0041358 1.34215e-08 0 1.36185e-08 0 1.362e-08 0.0041358 1.36215e-08 0 1.38185e-08 0 1.382e-08 0.0041358 1.38215e-08 0 1.40185e-08 0 1.402e-08 0.0041358 1.40215e-08 0 1.42185e-08 0 1.422e-08 0.0041358 1.42215e-08 0 1.44185e-08 0 1.442e-08 0.0041358 1.44215e-08 0 1.46185e-08 0 1.462e-08 0.0041358 1.46215e-08 0 1.48185e-08 0 1.482e-08 0.0041358 1.48215e-08 0 1.50185e-08 0 1.502e-08 0.0041358 1.50215e-08 0 1.52185e-08 0 1.522e-08 0.0041358 1.52215e-08 0 1.54185e-08 0 1.542e-08 0.0041358 1.54215e-08 0 1.56185e-08 0 1.562e-08 0.0041358 1.56215e-08 0 1.58185e-08 0 1.582e-08 0.0041358 1.58215e-08 0 1.60185e-08 0 1.602e-08 0.0041358 1.60215e-08 0 1.62185e-08 0 1.622e-08 0.0041358 1.62215e-08 0 1.64185e-08 0 1.642e-08 0.0041358 1.64215e-08 0 1.66185e-08 0 1.662e-08 0.0041358 1.66215e-08 0 1.68185e-08 0 1.682e-08 0.0041358 1.68215e-08 0 1.70185e-08 0 1.702e-08 0.0041358 1.70215e-08 0 1.72185e-08 0 1.722e-08 0.0041358 1.72215e-08 0 1.74185e-08 0 1.742e-08 0.0041358 1.74215e-08 0 1.76185e-08 0 1.762e-08 0.0041358 1.76215e-08 0 1.78185e-08 0 1.782e-08 0.0041358 1.78215e-08 0 1.80185e-08 0 1.802e-08 0.0041358 1.80215e-08 0 1.82185e-08 0 1.822e-08 0.0041358 1.82215e-08 0 1.84185e-08 0 1.842e-08 0.0041358 1.84215e-08 0 1.86185e-08 0 1.862e-08 0.0041358 1.86215e-08 0 1.88185e-08 0 1.882e-08 0.0041358 1.88215e-08 0 1.90185e-08 0 1.902e-08 0.0041358 1.90215e-08 0 1.92185e-08 0 1.922e-08 0.0041358 1.92215e-08 0 1.94185e-08 0 1.942e-08 0.0041358 1.94215e-08 0 1.96185e-08 0 1.962e-08 0.0041358 1.96215e-08 0 1.98185e-08 0 1.982e-08 0.0041358 1.98215e-08 0 2.00185e-08 0 2.002e-08 0.0041358 2.00215e-08 0 2.02185e-08 0 2.022e-08 0.0041358 2.02215e-08 0 2.04185e-08 0 2.042e-08 0.0041358 2.04215e-08 0 2.06185e-08 0 2.062e-08 0.0041358 2.06215e-08 0 2.08185e-08 0 2.082e-08 0.0041358 2.08215e-08 0 2.10185e-08 0 2.102e-08 0.0041358 2.10215e-08 0 2.12185e-08 0 2.122e-08 0.0041358 2.12215e-08 0 2.14185e-08 0 2.142e-08 0.0041358 2.14215e-08 0 2.16185e-08 0 2.162e-08 0.0041358 2.16215e-08 0 2.18185e-08 0 2.182e-08 0.0041358 2.18215e-08 0 2.20185e-08 0 2.202e-08 0.0041358 2.20215e-08 0 2.22185e-08 0 2.222e-08 0.0041358 2.22215e-08 0 2.24185e-08 0 2.242e-08 0.0041358 2.24215e-08 0 2.26185e-08 0 2.262e-08 0.0041358 2.26215e-08 0 2.28185e-08 0 2.282e-08 0.0041358 2.28215e-08 0 2.30185e-08 0 2.302e-08 0.0041358 2.30215e-08 0 2.32185e-08 0 2.322e-08 0.0041358 2.32215e-08 0 2.34185e-08 0 2.342e-08 0.0041358 2.34215e-08 0 2.36185e-08 0 2.362e-08 0.0041358 2.36215e-08 0 2.38185e-08 0 2.382e-08 0.0041358 2.38215e-08 0 2.40185e-08 0 2.402e-08 0.0041358 2.40215e-08 0 2.42185e-08 0 2.422e-08 0.0041358 2.42215e-08 0 2.44185e-08 0 2.442e-08 0.0041358 2.44215e-08 0 2.46185e-08 0 2.462e-08 0.0041358 2.46215e-08 0 2.48185e-08 0 2.482e-08 0.0041358 2.48215e-08 0 2.50185e-08 0 2.502e-08 0.0041358 2.50215e-08 0 2.52185e-08 0 2.522e-08 0.0041358 2.52215e-08 0 2.54185e-08 0 2.542e-08 0.0041358 2.54215e-08 0 2.56185e-08 0 2.562e-08 0.0041358 2.56215e-08 0 2.58185e-08 0 2.582e-08 0.0041358 2.58215e-08 0 2.60185e-08 0 2.602e-08 0.0041358 2.60215e-08 0 2.62185e-08 0 2.622e-08 0.0041358 2.62215e-08 0 2.64185e-08 0 2.642e-08 0.0041358 2.64215e-08 0 2.66185e-08 0 2.662e-08 0.0041358 2.66215e-08 0 2.68185e-08 0 2.682e-08 0.0041358 2.68215e-08 0 2.70185e-08 0 2.702e-08 0.0041358 2.70215e-08 0 2.72185e-08 0 2.722e-08 0.0041358 2.72215e-08 0 2.74185e-08 0 2.742e-08 0.0041358 2.74215e-08 0 2.76185e-08 0 2.762e-08 0.0041358 2.76215e-08 0 2.78185e-08 0 2.782e-08 0.0041358 2.78215e-08 0 2.80185e-08 0 2.802e-08 0.0041358 2.80215e-08 0 2.82185e-08 0 2.822e-08 0.0041358 2.82215e-08 0 2.84185e-08 0 2.842e-08 0.0041358 2.84215e-08 0 2.86185e-08 0 2.862e-08 0.0041358 2.86215e-08 0 2.88185e-08 0 2.882e-08 0.0041358 2.88215e-08 0 2.90185e-08 0 2.902e-08 0.0041358 2.90215e-08 0 2.92185e-08 0 2.922e-08 0.0041358 2.92215e-08 0 2.94185e-08 0 2.942e-08 0.0041358 2.94215e-08 0 2.96185e-08 0 2.962e-08 0.0041358 2.96215e-08 0 2.98185e-08 0 2.982e-08 0.0041358 2.98215e-08 0 3.00185e-08 0 3.002e-08 0.0041358 3.00215e-08 0 3.02185e-08 0 3.022e-08 0.0041358 3.02215e-08 0 3.04185e-08 0 3.042e-08 0.0041358 3.04215e-08 0 3.06185e-08 0 3.062e-08 0.0041358 3.06215e-08 0 3.08185e-08 0 3.082e-08 0.0041358 3.08215e-08 0 3.10185e-08 0 3.102e-08 0.0041358 3.10215e-08 0 3.12185e-08 0 3.122e-08 0.0041358 3.12215e-08 0 3.14185e-08 0 3.142e-08 0.0041358 3.14215e-08 0 3.16185e-08 0 3.162e-08 0.0041358 3.16215e-08 0 3.18185e-08 0 3.182e-08 0.0041358 3.18215e-08 0 3.20185e-08 0 3.202e-08 0.0041358 3.20215e-08 0 3.22185e-08 0 3.222e-08 0.0041358 3.22215e-08 0 3.24185e-08 0 3.242e-08 0.0041358 3.24215e-08 0 3.26185e-08 0 3.262e-08 0.0041358 3.26215e-08 0 3.28185e-08 0 3.282e-08 0.0041358 3.28215e-08 0 3.30185e-08 0 3.302e-08 0.0041358 3.30215e-08 0 3.32185e-08 0 3.322e-08 0.0041358 3.32215e-08 0 3.34185e-08 0 3.342e-08 0.0041358 3.34215e-08 0 3.36185e-08 0 3.362e-08 0.0041358 3.36215e-08 0 3.38185e-08 0 3.382e-08 0.0041358 3.38215e-08 0 3.40185e-08 0 3.402e-08 0.0041358 3.40215e-08 0 3.42185e-08 0 3.422e-08 0.0041358 3.42215e-08 0 3.44185e-08 0 3.442e-08 0.0041358 3.44215e-08 0 3.46185e-08 0 3.462e-08 0.0041358 3.46215e-08 0 3.48185e-08 0 3.482e-08 0.0041358 3.48215e-08 0 3.50185e-08 0 3.502e-08 0.0041358 3.50215e-08 0 3.52185e-08 0 3.522e-08 0.0041358 3.52215e-08 0 3.54185e-08 0 3.542e-08 0.0041358 3.54215e-08 0 3.56185e-08 0 3.562e-08 0.0041358 3.56215e-08 0 3.58185e-08 0 3.582e-08 0.0041358 3.58215e-08 0 3.60185e-08 0 3.602e-08 0.0041358 3.60215e-08 0 3.62185e-08 0 3.622e-08 0.0041358 3.62215e-08 0 3.64185e-08 0 3.642e-08 0.0041358 3.64215e-08 0 3.66185e-08 0 3.662e-08 0.0041358 3.66215e-08 0 3.68185e-08 0 3.682e-08 0.0041358 3.68215e-08 0 3.70185e-08 0 3.702e-08 0.0041358 3.70215e-08 0 3.72185e-08 0 3.722e-08 0.0041358 3.72215e-08 0 3.74185e-08 0 3.742e-08 0.0041358 3.74215e-08 0 3.76185e-08 0 3.762e-08 0.0041358 3.76215e-08 0 3.78185e-08 0 3.782e-08 0.0041358 3.78215e-08 0 3.80185e-08 0 3.802e-08 0.0041358 3.80215e-08 0 3.82185e-08 0 3.822e-08 0.0041358 3.82215e-08 0 3.84185e-08 0 3.842e-08 0.0041358 3.84215e-08 0 3.86185e-08 0 3.862e-08 0.0041358 3.86215e-08 0 3.88185e-08 0 3.882e-08 0.0041358 3.88215e-08 0 3.90185e-08 0 3.902e-08 0.0041358 3.90215e-08 0 3.92185e-08 0 3.922e-08 0.0041358 3.92215e-08 0 3.94185e-08 0 3.942e-08 0.0041358 3.94215e-08 0 3.96185e-08 0 3.962e-08 0.0041358 3.96215e-08 0 3.98185e-08 0 3.982e-08 0.0041358 3.98215e-08 0 4.00185e-08 0 4.002e-08 0.0041358 4.00215e-08 0 4.02185e-08 0 4.022e-08 0.0041358 4.02215e-08 0 4.04185e-08 0 4.042e-08 0.0041358 4.04215e-08 0 4.06185e-08 0 4.062e-08 0.0041358 4.06215e-08 0 4.08185e-08 0 4.082e-08 0.0041358 4.08215e-08 0 4.10185e-08 0 4.102e-08 0.0041358 4.10215e-08 0 4.12185e-08 0 4.122e-08 0.0041358 4.12215e-08 0 4.14185e-08 0 4.142e-08 0.0041358 4.14215e-08 0 4.16185e-08 0 4.162e-08 0.0041358 4.16215e-08 0 4.18185e-08 0 4.182e-08 0.0041358 4.18215e-08 0 4.20185e-08 0 4.202e-08 0.0041358 4.20215e-08 0 4.22185e-08 0 4.222e-08 0.0041358 4.22215e-08 0 4.24185e-08 0 4.242e-08 0.0041358 4.24215e-08 0 4.26185e-08 0 4.262e-08 0.0041358 4.26215e-08 0 4.28185e-08 0 4.282e-08 0.0041358 4.28215e-08 0 4.30185e-08 0 4.302e-08 0.0041358 4.30215e-08 0 4.32185e-08 0 4.322e-08 0.0041358 4.32215e-08 0 4.34185e-08 0 4.342e-08 0.0041358 4.34215e-08 0 4.36185e-08 0 4.362e-08 0.0041358 4.36215e-08 0 4.38185e-08 0 4.382e-08 0.0041358 4.38215e-08 0 4.40185e-08 0 4.402e-08 0.0041358 4.40215e-08 0 4.42185e-08 0 4.422e-08 0.0041358 4.42215e-08 0 4.44185e-08 0 4.442e-08 0.0041358 4.44215e-08 0 4.46185e-08 0 4.462e-08 0.0041358 4.46215e-08 0 4.48185e-08 0 4.482e-08 0.0041358 4.48215e-08 0 4.50185e-08 0 4.502e-08 0.0041358 4.50215e-08 0 4.52185e-08 0 4.522e-08 0.0041358 4.52215e-08 0 4.54185e-08 0 4.542e-08 0.0041358 4.54215e-08 0 4.56185e-08 0 4.562e-08 0.0041358 4.56215e-08 0 4.58185e-08 0 4.582e-08 0.0041358 4.58215e-08 0 4.60185e-08 0 4.602e-08 0.0041358 4.60215e-08 0 4.62185e-08 0 4.622e-08 0.0041358 4.62215e-08 0 4.64185e-08 0 4.642e-08 0.0041358 4.64215e-08 0 4.66185e-08 0 4.662e-08 0.0041358 4.66215e-08 0 4.68185e-08 0 4.682e-08 0.0041358 4.68215e-08 0 4.70185e-08 0 4.702e-08 0.0041358 4.70215e-08 0 4.72185e-08 0 4.722e-08 0.0041358 4.72215e-08 0 4.74185e-08 0 4.742e-08 0.0041358 4.74215e-08 0 4.76185e-08 0 4.762e-08 0.0041358 4.76215e-08 0 4.78185e-08 0 4.782e-08 0.0041358 4.78215e-08 0 4.80185e-08 0 4.802e-08 0.0041358 4.80215e-08 0 4.82185e-08 0 4.822e-08 0.0041358 4.82215e-08 0 4.84185e-08 0 4.842e-08 0.0041358 4.84215e-08 0 4.86185e-08 0 4.862e-08 0.0041358 4.86215e-08 0 4.88185e-08 0 4.882e-08 0.0041358 4.88215e-08 0 4.90185e-08 0 4.902e-08 0.0041358 4.90215e-08 0 4.92185e-08 0 4.922e-08 0.0041358 4.92215e-08 0 4.94185e-08 0 4.942e-08 0.0041358 4.94215e-08 0 4.96185e-08 0 4.962e-08 0.0041358 4.96215e-08 0 4.98185e-08 0 4.982e-08 0.0041358 4.98215e-08 0 5.00185e-08 0 5.002e-08 0.0041358 5.00215e-08 0 5.02185e-08 0 5.022e-08 0.0041358 5.02215e-08 0 5.04185e-08 0 5.042e-08 0.0041358 5.04215e-08 0 5.06185e-08 0 5.062e-08 0.0041358 5.06215e-08 0 5.08185e-08 0 5.082e-08 0.0041358 5.08215e-08 0 5.10185e-08 0 5.102e-08 0.0041358 5.10215e-08 0)
IT01_|T 0 T01_  PWL(0 0 1.85e-11 0 2e-11 0.0041358 2.15e-11 0 2.185e-10 0 2.2e-10 0.0041358 2.215e-10 0 4.185e-10 0 4.2e-10 0.0041358 4.215e-10 0 6.185e-10 0 6.2e-10 0.0041358 6.215e-10 0 8.185e-10 0 8.2e-10 0.0041358 8.215e-10 0 1.0185e-09 0 1.02e-09 0.0041358 1.0215e-09 0 1.2185e-09 0 1.22e-09 0.0041358 1.2215e-09 0 1.4185e-09 0 1.42e-09 0.0041358 1.4215e-09 0 1.6185e-09 0 1.62e-09 0.0041358 1.6215e-09 0 1.8185e-09 0 1.82e-09 0.0041358 1.8215e-09 0 2.0185e-09 0 2.02e-09 0.0041358 2.0215e-09 0 2.2185e-09 0 2.22e-09 0.0041358 2.2215e-09 0 2.4185e-09 0 2.42e-09 0.0041358 2.4215e-09 0 2.6185e-09 0 2.62e-09 0.0041358 2.6215e-09 0 2.8185e-09 0 2.82e-09 0.0041358 2.8215e-09 0 3.0185e-09 0 3.02e-09 0.0041358 3.0215e-09 0 3.2185e-09 0 3.22e-09 0.0041358 3.2215e-09 0 3.4185e-09 0 3.42e-09 0.0041358 3.4215e-09 0 3.6185e-09 0 3.62e-09 0.0041358 3.6215e-09 0 3.8185e-09 0 3.82e-09 0.0041358 3.8215e-09 0 4.0185e-09 0 4.02e-09 0.0041358 4.0215e-09 0 4.2185e-09 0 4.22e-09 0.0041358 4.2215e-09 0 4.4185e-09 0 4.42e-09 0.0041358 4.4215e-09 0 4.6185e-09 0 4.62e-09 0.0041358 4.6215e-09 0 4.8185e-09 0 4.82e-09 0.0041358 4.8215e-09 0 5.0185e-09 0 5.02e-09 0.0041358 5.0215e-09 0 5.2185e-09 0 5.22e-09 0.0041358 5.2215e-09 0 5.4185e-09 0 5.42e-09 0.0041358 5.4215e-09 0 5.6185e-09 0 5.62e-09 0.0041358 5.6215e-09 0 5.8185e-09 0 5.82e-09 0.0041358 5.8215e-09 0 6.0185e-09 0 6.02e-09 0.0041358 6.0215e-09 0 6.2185e-09 0 6.22e-09 0.0041358 6.2215e-09 0 6.4185e-09 0 6.42e-09 0.0041358 6.4215e-09 0 6.6185e-09 0 6.62e-09 0.0041358 6.6215e-09 0 6.8185e-09 0 6.82e-09 0.0041358 6.8215e-09 0 7.0185e-09 0 7.02e-09 0.0041358 7.0215e-09 0 7.2185e-09 0 7.22e-09 0.0041358 7.2215e-09 0 7.4185e-09 0 7.42e-09 0.0041358 7.4215e-09 0 7.6185e-09 0 7.62e-09 0.0041358 7.6215e-09 0 7.8185e-09 0 7.82e-09 0.0041358 7.8215e-09 0 8.0185e-09 0 8.02e-09 0.0041358 8.0215e-09 0 8.2185e-09 0 8.22e-09 0.0041358 8.2215e-09 0 8.4185e-09 0 8.42e-09 0.0041358 8.4215e-09 0 8.6185e-09 0 8.62e-09 0.0041358 8.6215e-09 0 8.8185e-09 0 8.82e-09 0.0041358 8.8215e-09 0 9.0185e-09 0 9.02e-09 0.0041358 9.0215e-09 0 9.2185e-09 0 9.22e-09 0.0041358 9.2215e-09 0 9.4185e-09 0 9.42e-09 0.0041358 9.4215e-09 0 9.6185e-09 0 9.62e-09 0.0041358 9.6215e-09 0 9.8185e-09 0 9.82e-09 0.0041358 9.8215e-09 0 1.00185e-08 0 1.002e-08 0.0041358 1.00215e-08 0 1.02185e-08 0 1.022e-08 0.0041358 1.02215e-08 0 1.04185e-08 0 1.042e-08 0.0041358 1.04215e-08 0 1.06185e-08 0 1.062e-08 0.0041358 1.06215e-08 0 1.08185e-08 0 1.082e-08 0.0041358 1.08215e-08 0 1.10185e-08 0 1.102e-08 0.0041358 1.10215e-08 0 1.12185e-08 0 1.122e-08 0.0041358 1.12215e-08 0 1.14185e-08 0 1.142e-08 0.0041358 1.14215e-08 0 1.16185e-08 0 1.162e-08 0.0041358 1.16215e-08 0 1.18185e-08 0 1.182e-08 0.0041358 1.18215e-08 0 1.20185e-08 0 1.202e-08 0.0041358 1.20215e-08 0 1.22185e-08 0 1.222e-08 0.0041358 1.22215e-08 0 1.24185e-08 0 1.242e-08 0.0041358 1.24215e-08 0 1.26185e-08 0 1.262e-08 0.0041358 1.26215e-08 0 1.28185e-08 0 1.282e-08 0.0041358 1.28215e-08 0 1.30185e-08 0 1.302e-08 0.0041358 1.30215e-08 0 1.32185e-08 0 1.322e-08 0.0041358 1.32215e-08 0 1.34185e-08 0 1.342e-08 0.0041358 1.34215e-08 0 1.36185e-08 0 1.362e-08 0.0041358 1.36215e-08 0 1.38185e-08 0 1.382e-08 0.0041358 1.38215e-08 0 1.40185e-08 0 1.402e-08 0.0041358 1.40215e-08 0 1.42185e-08 0 1.422e-08 0.0041358 1.42215e-08 0 1.44185e-08 0 1.442e-08 0.0041358 1.44215e-08 0 1.46185e-08 0 1.462e-08 0.0041358 1.46215e-08 0 1.48185e-08 0 1.482e-08 0.0041358 1.48215e-08 0 1.50185e-08 0 1.502e-08 0.0041358 1.50215e-08 0 1.52185e-08 0 1.522e-08 0.0041358 1.52215e-08 0 1.54185e-08 0 1.542e-08 0.0041358 1.54215e-08 0 1.56185e-08 0 1.562e-08 0.0041358 1.56215e-08 0 1.58185e-08 0 1.582e-08 0.0041358 1.58215e-08 0 1.60185e-08 0 1.602e-08 0.0041358 1.60215e-08 0 1.62185e-08 0 1.622e-08 0.0041358 1.62215e-08 0 1.64185e-08 0 1.642e-08 0.0041358 1.64215e-08 0 1.66185e-08 0 1.662e-08 0.0041358 1.66215e-08 0 1.68185e-08 0 1.682e-08 0.0041358 1.68215e-08 0 1.70185e-08 0 1.702e-08 0.0041358 1.70215e-08 0 1.72185e-08 0 1.722e-08 0.0041358 1.72215e-08 0 1.74185e-08 0 1.742e-08 0.0041358 1.74215e-08 0 1.76185e-08 0 1.762e-08 0.0041358 1.76215e-08 0 1.78185e-08 0 1.782e-08 0.0041358 1.78215e-08 0 1.80185e-08 0 1.802e-08 0.0041358 1.80215e-08 0 1.82185e-08 0 1.822e-08 0.0041358 1.82215e-08 0 1.84185e-08 0 1.842e-08 0.0041358 1.84215e-08 0 1.86185e-08 0 1.862e-08 0.0041358 1.86215e-08 0 1.88185e-08 0 1.882e-08 0.0041358 1.88215e-08 0 1.90185e-08 0 1.902e-08 0.0041358 1.90215e-08 0 1.92185e-08 0 1.922e-08 0.0041358 1.92215e-08 0 1.94185e-08 0 1.942e-08 0.0041358 1.94215e-08 0 1.96185e-08 0 1.962e-08 0.0041358 1.96215e-08 0 1.98185e-08 0 1.982e-08 0.0041358 1.98215e-08 0 2.00185e-08 0 2.002e-08 0.0041358 2.00215e-08 0 2.02185e-08 0 2.022e-08 0.0041358 2.02215e-08 0 2.04185e-08 0 2.042e-08 0.0041358 2.04215e-08 0 2.06185e-08 0 2.062e-08 0.0041358 2.06215e-08 0 2.08185e-08 0 2.082e-08 0.0041358 2.08215e-08 0 2.10185e-08 0 2.102e-08 0.0041358 2.10215e-08 0 2.12185e-08 0 2.122e-08 0.0041358 2.12215e-08 0 2.14185e-08 0 2.142e-08 0.0041358 2.14215e-08 0 2.16185e-08 0 2.162e-08 0.0041358 2.16215e-08 0 2.18185e-08 0 2.182e-08 0.0041358 2.18215e-08 0 2.20185e-08 0 2.202e-08 0.0041358 2.20215e-08 0 2.22185e-08 0 2.222e-08 0.0041358 2.22215e-08 0 2.24185e-08 0 2.242e-08 0.0041358 2.24215e-08 0 2.26185e-08 0 2.262e-08 0.0041358 2.26215e-08 0 2.28185e-08 0 2.282e-08 0.0041358 2.28215e-08 0 2.30185e-08 0 2.302e-08 0.0041358 2.30215e-08 0 2.32185e-08 0 2.322e-08 0.0041358 2.32215e-08 0 2.34185e-08 0 2.342e-08 0.0041358 2.34215e-08 0 2.36185e-08 0 2.362e-08 0.0041358 2.36215e-08 0 2.38185e-08 0 2.382e-08 0.0041358 2.38215e-08 0 2.40185e-08 0 2.402e-08 0.0041358 2.40215e-08 0 2.42185e-08 0 2.422e-08 0.0041358 2.42215e-08 0 2.44185e-08 0 2.442e-08 0.0041358 2.44215e-08 0 2.46185e-08 0 2.462e-08 0.0041358 2.46215e-08 0 2.48185e-08 0 2.482e-08 0.0041358 2.48215e-08 0 2.50185e-08 0 2.502e-08 0.0041358 2.50215e-08 0 2.52185e-08 0 2.522e-08 0.0041358 2.52215e-08 0 2.54185e-08 0 2.542e-08 0.0041358 2.54215e-08 0 2.56185e-08 0 2.562e-08 0.0041358 2.56215e-08 0 2.58185e-08 0 2.582e-08 0.0041358 2.58215e-08 0 2.60185e-08 0 2.602e-08 0.0041358 2.60215e-08 0 2.62185e-08 0 2.622e-08 0.0041358 2.62215e-08 0 2.64185e-08 0 2.642e-08 0.0041358 2.64215e-08 0 2.66185e-08 0 2.662e-08 0.0041358 2.66215e-08 0 2.68185e-08 0 2.682e-08 0.0041358 2.68215e-08 0 2.70185e-08 0 2.702e-08 0.0041358 2.70215e-08 0 2.72185e-08 0 2.722e-08 0.0041358 2.72215e-08 0 2.74185e-08 0 2.742e-08 0.0041358 2.74215e-08 0 2.76185e-08 0 2.762e-08 0.0041358 2.76215e-08 0 2.78185e-08 0 2.782e-08 0.0041358 2.78215e-08 0 2.80185e-08 0 2.802e-08 0.0041358 2.80215e-08 0 2.82185e-08 0 2.822e-08 0.0041358 2.82215e-08 0 2.84185e-08 0 2.842e-08 0.0041358 2.84215e-08 0 2.86185e-08 0 2.862e-08 0.0041358 2.86215e-08 0 2.88185e-08 0 2.882e-08 0.0041358 2.88215e-08 0 2.90185e-08 0 2.902e-08 0.0041358 2.90215e-08 0 2.92185e-08 0 2.922e-08 0.0041358 2.92215e-08 0 2.94185e-08 0 2.942e-08 0.0041358 2.94215e-08 0 2.96185e-08 0 2.962e-08 0.0041358 2.96215e-08 0 2.98185e-08 0 2.982e-08 0.0041358 2.98215e-08 0 3.00185e-08 0 3.002e-08 0.0041358 3.00215e-08 0 3.02185e-08 0 3.022e-08 0.0041358 3.02215e-08 0 3.04185e-08 0 3.042e-08 0.0041358 3.04215e-08 0 3.06185e-08 0 3.062e-08 0.0041358 3.06215e-08 0 3.08185e-08 0 3.082e-08 0.0041358 3.08215e-08 0 3.10185e-08 0 3.102e-08 0.0041358 3.10215e-08 0 3.12185e-08 0 3.122e-08 0.0041358 3.12215e-08 0 3.14185e-08 0 3.142e-08 0.0041358 3.14215e-08 0 3.16185e-08 0 3.162e-08 0.0041358 3.16215e-08 0 3.18185e-08 0 3.182e-08 0.0041358 3.18215e-08 0 3.20185e-08 0 3.202e-08 0.0041358 3.20215e-08 0 3.22185e-08 0 3.222e-08 0.0041358 3.22215e-08 0 3.24185e-08 0 3.242e-08 0.0041358 3.24215e-08 0 3.26185e-08 0 3.262e-08 0.0041358 3.26215e-08 0 3.28185e-08 0 3.282e-08 0.0041358 3.28215e-08 0 3.30185e-08 0 3.302e-08 0.0041358 3.30215e-08 0 3.32185e-08 0 3.322e-08 0.0041358 3.32215e-08 0 3.34185e-08 0 3.342e-08 0.0041358 3.34215e-08 0 3.36185e-08 0 3.362e-08 0.0041358 3.36215e-08 0 3.38185e-08 0 3.382e-08 0.0041358 3.38215e-08 0 3.40185e-08 0 3.402e-08 0.0041358 3.40215e-08 0 3.42185e-08 0 3.422e-08 0.0041358 3.42215e-08 0 3.44185e-08 0 3.442e-08 0.0041358 3.44215e-08 0 3.46185e-08 0 3.462e-08 0.0041358 3.46215e-08 0 3.48185e-08 0 3.482e-08 0.0041358 3.48215e-08 0 3.50185e-08 0 3.502e-08 0.0041358 3.50215e-08 0 3.52185e-08 0 3.522e-08 0.0041358 3.52215e-08 0 3.54185e-08 0 3.542e-08 0.0041358 3.54215e-08 0 3.56185e-08 0 3.562e-08 0.0041358 3.56215e-08 0 3.58185e-08 0 3.582e-08 0.0041358 3.58215e-08 0 3.60185e-08 0 3.602e-08 0.0041358 3.60215e-08 0 3.62185e-08 0 3.622e-08 0.0041358 3.62215e-08 0 3.64185e-08 0 3.642e-08 0.0041358 3.64215e-08 0 3.66185e-08 0 3.662e-08 0.0041358 3.66215e-08 0 3.68185e-08 0 3.682e-08 0.0041358 3.68215e-08 0 3.70185e-08 0 3.702e-08 0.0041358 3.70215e-08 0 3.72185e-08 0 3.722e-08 0.0041358 3.72215e-08 0 3.74185e-08 0 3.742e-08 0.0041358 3.74215e-08 0 3.76185e-08 0 3.762e-08 0.0041358 3.76215e-08 0 3.78185e-08 0 3.782e-08 0.0041358 3.78215e-08 0 3.80185e-08 0 3.802e-08 0.0041358 3.80215e-08 0 3.82185e-08 0 3.822e-08 0.0041358 3.82215e-08 0 3.84185e-08 0 3.842e-08 0.0041358 3.84215e-08 0 3.86185e-08 0 3.862e-08 0.0041358 3.86215e-08 0 3.88185e-08 0 3.882e-08 0.0041358 3.88215e-08 0 3.90185e-08 0 3.902e-08 0.0041358 3.90215e-08 0 3.92185e-08 0 3.922e-08 0.0041358 3.92215e-08 0 3.94185e-08 0 3.942e-08 0.0041358 3.94215e-08 0 3.96185e-08 0 3.962e-08 0.0041358 3.96215e-08 0 3.98185e-08 0 3.982e-08 0.0041358 3.98215e-08 0 4.00185e-08 0 4.002e-08 0.0041358 4.00215e-08 0 4.02185e-08 0 4.022e-08 0.0041358 4.02215e-08 0 4.04185e-08 0 4.042e-08 0.0041358 4.04215e-08 0 4.06185e-08 0 4.062e-08 0.0041358 4.06215e-08 0 4.08185e-08 0 4.082e-08 0.0041358 4.08215e-08 0 4.10185e-08 0 4.102e-08 0.0041358 4.10215e-08 0 4.12185e-08 0 4.122e-08 0.0041358 4.12215e-08 0 4.14185e-08 0 4.142e-08 0.0041358 4.14215e-08 0 4.16185e-08 0 4.162e-08 0.0041358 4.16215e-08 0 4.18185e-08 0 4.182e-08 0.0041358 4.18215e-08 0 4.20185e-08 0 4.202e-08 0.0041358 4.20215e-08 0 4.22185e-08 0 4.222e-08 0.0041358 4.22215e-08 0 4.24185e-08 0 4.242e-08 0.0041358 4.24215e-08 0 4.26185e-08 0 4.262e-08 0.0041358 4.26215e-08 0 4.28185e-08 0 4.282e-08 0.0041358 4.28215e-08 0 4.30185e-08 0 4.302e-08 0.0041358 4.30215e-08 0 4.32185e-08 0 4.322e-08 0.0041358 4.32215e-08 0 4.34185e-08 0 4.342e-08 0.0041358 4.34215e-08 0 4.36185e-08 0 4.362e-08 0.0041358 4.36215e-08 0 4.38185e-08 0 4.382e-08 0.0041358 4.38215e-08 0 4.40185e-08 0 4.402e-08 0.0041358 4.40215e-08 0 4.42185e-08 0 4.422e-08 0.0041358 4.42215e-08 0 4.44185e-08 0 4.442e-08 0.0041358 4.44215e-08 0 4.46185e-08 0 4.462e-08 0.0041358 4.46215e-08 0 4.48185e-08 0 4.482e-08 0.0041358 4.48215e-08 0 4.50185e-08 0 4.502e-08 0.0041358 4.50215e-08 0 4.52185e-08 0 4.522e-08 0.0041358 4.52215e-08 0 4.54185e-08 0 4.542e-08 0.0041358 4.54215e-08 0 4.56185e-08 0 4.562e-08 0.0041358 4.56215e-08 0 4.58185e-08 0 4.582e-08 0.0041358 4.58215e-08 0 4.60185e-08 0 4.602e-08 0.0041358 4.60215e-08 0 4.62185e-08 0 4.622e-08 0.0041358 4.62215e-08 0 4.64185e-08 0 4.642e-08 0.0041358 4.64215e-08 0 4.66185e-08 0 4.662e-08 0.0041358 4.66215e-08 0 4.68185e-08 0 4.682e-08 0.0041358 4.68215e-08 0 4.70185e-08 0 4.702e-08 0.0041358 4.70215e-08 0 4.72185e-08 0 4.722e-08 0.0041358 4.72215e-08 0 4.74185e-08 0 4.742e-08 0.0041358 4.74215e-08 0 4.76185e-08 0 4.762e-08 0.0041358 4.76215e-08 0 4.78185e-08 0 4.782e-08 0.0041358 4.78215e-08 0 4.80185e-08 0 4.802e-08 0.0041358 4.80215e-08 0 4.82185e-08 0 4.822e-08 0.0041358 4.82215e-08 0 4.84185e-08 0 4.842e-08 0.0041358 4.84215e-08 0 4.86185e-08 0 4.862e-08 0.0041358 4.86215e-08 0 4.88185e-08 0 4.882e-08 0.0041358 4.88215e-08 0 4.90185e-08 0 4.902e-08 0.0041358 4.90215e-08 0 4.92185e-08 0 4.922e-08 0.0041358 4.92215e-08 0 4.94185e-08 0 4.942e-08 0.0041358 4.94215e-08 0 4.96185e-08 0 4.962e-08 0.0041358 4.96215e-08 0 4.98185e-08 0 4.982e-08 0.0041358 4.98215e-08 0 5.00185e-08 0 5.002e-08 0.0041358 5.00215e-08 0 5.02185e-08 0 5.022e-08 0.0041358 5.02215e-08 0 5.04185e-08 0 5.042e-08 0.0041358 5.04215e-08 0 5.06185e-08 0 5.062e-08 0.0041358 5.06215e-08 0 5.08185e-08 0 5.082e-08 0.0041358 5.08215e-08 0 5.10185e-08 0 5.102e-08 0.0041358 5.10215e-08 0)
IT02_|T 0 T02_  PWL(0 0 1.85e-11 0 2e-11 0.0041358 2.15e-11 0 2.185e-10 0 2.2e-10 0.0041358 2.215e-10 0 4.185e-10 0 4.2e-10 0.0041358 4.215e-10 0 6.185e-10 0 6.2e-10 0.0041358 6.215e-10 0 8.185e-10 0 8.2e-10 0.0041358 8.215e-10 0 1.0185e-09 0 1.02e-09 0.0041358 1.0215e-09 0 1.2185e-09 0 1.22e-09 0.0041358 1.2215e-09 0 1.4185e-09 0 1.42e-09 0.0041358 1.4215e-09 0 1.6185e-09 0 1.62e-09 0.0041358 1.6215e-09 0 1.8185e-09 0 1.82e-09 0.0041358 1.8215e-09 0 2.0185e-09 0 2.02e-09 0.0041358 2.0215e-09 0 2.2185e-09 0 2.22e-09 0.0041358 2.2215e-09 0 2.4185e-09 0 2.42e-09 0.0041358 2.4215e-09 0 2.6185e-09 0 2.62e-09 0.0041358 2.6215e-09 0 2.8185e-09 0 2.82e-09 0.0041358 2.8215e-09 0 3.0185e-09 0 3.02e-09 0.0041358 3.0215e-09 0 3.2185e-09 0 3.22e-09 0.0041358 3.2215e-09 0 3.4185e-09 0 3.42e-09 0.0041358 3.4215e-09 0 3.6185e-09 0 3.62e-09 0.0041358 3.6215e-09 0 3.8185e-09 0 3.82e-09 0.0041358 3.8215e-09 0 4.0185e-09 0 4.02e-09 0.0041358 4.0215e-09 0 4.2185e-09 0 4.22e-09 0.0041358 4.2215e-09 0 4.4185e-09 0 4.42e-09 0.0041358 4.4215e-09 0 4.6185e-09 0 4.62e-09 0.0041358 4.6215e-09 0 4.8185e-09 0 4.82e-09 0.0041358 4.8215e-09 0 5.0185e-09 0 5.02e-09 0.0041358 5.0215e-09 0 5.2185e-09 0 5.22e-09 0.0041358 5.2215e-09 0 5.4185e-09 0 5.42e-09 0.0041358 5.4215e-09 0 5.6185e-09 0 5.62e-09 0.0041358 5.6215e-09 0 5.8185e-09 0 5.82e-09 0.0041358 5.8215e-09 0 6.0185e-09 0 6.02e-09 0.0041358 6.0215e-09 0 6.2185e-09 0 6.22e-09 0.0041358 6.2215e-09 0 6.4185e-09 0 6.42e-09 0.0041358 6.4215e-09 0 6.6185e-09 0 6.62e-09 0.0041358 6.6215e-09 0 6.8185e-09 0 6.82e-09 0.0041358 6.8215e-09 0 7.0185e-09 0 7.02e-09 0.0041358 7.0215e-09 0 7.2185e-09 0 7.22e-09 0.0041358 7.2215e-09 0 7.4185e-09 0 7.42e-09 0.0041358 7.4215e-09 0 7.6185e-09 0 7.62e-09 0.0041358 7.6215e-09 0 7.8185e-09 0 7.82e-09 0.0041358 7.8215e-09 0 8.0185e-09 0 8.02e-09 0.0041358 8.0215e-09 0 8.2185e-09 0 8.22e-09 0.0041358 8.2215e-09 0 8.4185e-09 0 8.42e-09 0.0041358 8.4215e-09 0 8.6185e-09 0 8.62e-09 0.0041358 8.6215e-09 0 8.8185e-09 0 8.82e-09 0.0041358 8.8215e-09 0 9.0185e-09 0 9.02e-09 0.0041358 9.0215e-09 0 9.2185e-09 0 9.22e-09 0.0041358 9.2215e-09 0 9.4185e-09 0 9.42e-09 0.0041358 9.4215e-09 0 9.6185e-09 0 9.62e-09 0.0041358 9.6215e-09 0 9.8185e-09 0 9.82e-09 0.0041358 9.8215e-09 0 1.00185e-08 0 1.002e-08 0.0041358 1.00215e-08 0 1.02185e-08 0 1.022e-08 0.0041358 1.02215e-08 0 1.04185e-08 0 1.042e-08 0.0041358 1.04215e-08 0 1.06185e-08 0 1.062e-08 0.0041358 1.06215e-08 0 1.08185e-08 0 1.082e-08 0.0041358 1.08215e-08 0 1.10185e-08 0 1.102e-08 0.0041358 1.10215e-08 0 1.12185e-08 0 1.122e-08 0.0041358 1.12215e-08 0 1.14185e-08 0 1.142e-08 0.0041358 1.14215e-08 0 1.16185e-08 0 1.162e-08 0.0041358 1.16215e-08 0 1.18185e-08 0 1.182e-08 0.0041358 1.18215e-08 0 1.20185e-08 0 1.202e-08 0.0041358 1.20215e-08 0 1.22185e-08 0 1.222e-08 0.0041358 1.22215e-08 0 1.24185e-08 0 1.242e-08 0.0041358 1.24215e-08 0 1.26185e-08 0 1.262e-08 0.0041358 1.26215e-08 0 1.28185e-08 0 1.282e-08 0.0041358 1.28215e-08 0 1.30185e-08 0 1.302e-08 0.0041358 1.30215e-08 0 1.32185e-08 0 1.322e-08 0.0041358 1.32215e-08 0 1.34185e-08 0 1.342e-08 0.0041358 1.34215e-08 0 1.36185e-08 0 1.362e-08 0.0041358 1.36215e-08 0 1.38185e-08 0 1.382e-08 0.0041358 1.38215e-08 0 1.40185e-08 0 1.402e-08 0.0041358 1.40215e-08 0 1.42185e-08 0 1.422e-08 0.0041358 1.42215e-08 0 1.44185e-08 0 1.442e-08 0.0041358 1.44215e-08 0 1.46185e-08 0 1.462e-08 0.0041358 1.46215e-08 0 1.48185e-08 0 1.482e-08 0.0041358 1.48215e-08 0 1.50185e-08 0 1.502e-08 0.0041358 1.50215e-08 0 1.52185e-08 0 1.522e-08 0.0041358 1.52215e-08 0 1.54185e-08 0 1.542e-08 0.0041358 1.54215e-08 0 1.56185e-08 0 1.562e-08 0.0041358 1.56215e-08 0 1.58185e-08 0 1.582e-08 0.0041358 1.58215e-08 0 1.60185e-08 0 1.602e-08 0.0041358 1.60215e-08 0 1.62185e-08 0 1.622e-08 0.0041358 1.62215e-08 0 1.64185e-08 0 1.642e-08 0.0041358 1.64215e-08 0 1.66185e-08 0 1.662e-08 0.0041358 1.66215e-08 0 1.68185e-08 0 1.682e-08 0.0041358 1.68215e-08 0 1.70185e-08 0 1.702e-08 0.0041358 1.70215e-08 0 1.72185e-08 0 1.722e-08 0.0041358 1.72215e-08 0 1.74185e-08 0 1.742e-08 0.0041358 1.74215e-08 0 1.76185e-08 0 1.762e-08 0.0041358 1.76215e-08 0 1.78185e-08 0 1.782e-08 0.0041358 1.78215e-08 0 1.80185e-08 0 1.802e-08 0.0041358 1.80215e-08 0 1.82185e-08 0 1.822e-08 0.0041358 1.82215e-08 0 1.84185e-08 0 1.842e-08 0.0041358 1.84215e-08 0 1.86185e-08 0 1.862e-08 0.0041358 1.86215e-08 0 1.88185e-08 0 1.882e-08 0.0041358 1.88215e-08 0 1.90185e-08 0 1.902e-08 0.0041358 1.90215e-08 0 1.92185e-08 0 1.922e-08 0.0041358 1.92215e-08 0 1.94185e-08 0 1.942e-08 0.0041358 1.94215e-08 0 1.96185e-08 0 1.962e-08 0.0041358 1.96215e-08 0 1.98185e-08 0 1.982e-08 0.0041358 1.98215e-08 0 2.00185e-08 0 2.002e-08 0.0041358 2.00215e-08 0 2.02185e-08 0 2.022e-08 0.0041358 2.02215e-08 0 2.04185e-08 0 2.042e-08 0.0041358 2.04215e-08 0 2.06185e-08 0 2.062e-08 0.0041358 2.06215e-08 0 2.08185e-08 0 2.082e-08 0.0041358 2.08215e-08 0 2.10185e-08 0 2.102e-08 0.0041358 2.10215e-08 0 2.12185e-08 0 2.122e-08 0.0041358 2.12215e-08 0 2.14185e-08 0 2.142e-08 0.0041358 2.14215e-08 0 2.16185e-08 0 2.162e-08 0.0041358 2.16215e-08 0 2.18185e-08 0 2.182e-08 0.0041358 2.18215e-08 0 2.20185e-08 0 2.202e-08 0.0041358 2.20215e-08 0 2.22185e-08 0 2.222e-08 0.0041358 2.22215e-08 0 2.24185e-08 0 2.242e-08 0.0041358 2.24215e-08 0 2.26185e-08 0 2.262e-08 0.0041358 2.26215e-08 0 2.28185e-08 0 2.282e-08 0.0041358 2.28215e-08 0 2.30185e-08 0 2.302e-08 0.0041358 2.30215e-08 0 2.32185e-08 0 2.322e-08 0.0041358 2.32215e-08 0 2.34185e-08 0 2.342e-08 0.0041358 2.34215e-08 0 2.36185e-08 0 2.362e-08 0.0041358 2.36215e-08 0 2.38185e-08 0 2.382e-08 0.0041358 2.38215e-08 0 2.40185e-08 0 2.402e-08 0.0041358 2.40215e-08 0 2.42185e-08 0 2.422e-08 0.0041358 2.42215e-08 0 2.44185e-08 0 2.442e-08 0.0041358 2.44215e-08 0 2.46185e-08 0 2.462e-08 0.0041358 2.46215e-08 0 2.48185e-08 0 2.482e-08 0.0041358 2.48215e-08 0 2.50185e-08 0 2.502e-08 0.0041358 2.50215e-08 0 2.52185e-08 0 2.522e-08 0.0041358 2.52215e-08 0 2.54185e-08 0 2.542e-08 0.0041358 2.54215e-08 0 2.56185e-08 0 2.562e-08 0.0041358 2.56215e-08 0 2.58185e-08 0 2.582e-08 0.0041358 2.58215e-08 0 2.60185e-08 0 2.602e-08 0.0041358 2.60215e-08 0 2.62185e-08 0 2.622e-08 0.0041358 2.62215e-08 0 2.64185e-08 0 2.642e-08 0.0041358 2.64215e-08 0 2.66185e-08 0 2.662e-08 0.0041358 2.66215e-08 0 2.68185e-08 0 2.682e-08 0.0041358 2.68215e-08 0 2.70185e-08 0 2.702e-08 0.0041358 2.70215e-08 0 2.72185e-08 0 2.722e-08 0.0041358 2.72215e-08 0 2.74185e-08 0 2.742e-08 0.0041358 2.74215e-08 0 2.76185e-08 0 2.762e-08 0.0041358 2.76215e-08 0 2.78185e-08 0 2.782e-08 0.0041358 2.78215e-08 0 2.80185e-08 0 2.802e-08 0.0041358 2.80215e-08 0 2.82185e-08 0 2.822e-08 0.0041358 2.82215e-08 0 2.84185e-08 0 2.842e-08 0.0041358 2.84215e-08 0 2.86185e-08 0 2.862e-08 0.0041358 2.86215e-08 0 2.88185e-08 0 2.882e-08 0.0041358 2.88215e-08 0 2.90185e-08 0 2.902e-08 0.0041358 2.90215e-08 0 2.92185e-08 0 2.922e-08 0.0041358 2.92215e-08 0 2.94185e-08 0 2.942e-08 0.0041358 2.94215e-08 0 2.96185e-08 0 2.962e-08 0.0041358 2.96215e-08 0 2.98185e-08 0 2.982e-08 0.0041358 2.98215e-08 0 3.00185e-08 0 3.002e-08 0.0041358 3.00215e-08 0 3.02185e-08 0 3.022e-08 0.0041358 3.02215e-08 0 3.04185e-08 0 3.042e-08 0.0041358 3.04215e-08 0 3.06185e-08 0 3.062e-08 0.0041358 3.06215e-08 0 3.08185e-08 0 3.082e-08 0.0041358 3.08215e-08 0 3.10185e-08 0 3.102e-08 0.0041358 3.10215e-08 0 3.12185e-08 0 3.122e-08 0.0041358 3.12215e-08 0 3.14185e-08 0 3.142e-08 0.0041358 3.14215e-08 0 3.16185e-08 0 3.162e-08 0.0041358 3.16215e-08 0 3.18185e-08 0 3.182e-08 0.0041358 3.18215e-08 0 3.20185e-08 0 3.202e-08 0.0041358 3.20215e-08 0 3.22185e-08 0 3.222e-08 0.0041358 3.22215e-08 0 3.24185e-08 0 3.242e-08 0.0041358 3.24215e-08 0 3.26185e-08 0 3.262e-08 0.0041358 3.26215e-08 0 3.28185e-08 0 3.282e-08 0.0041358 3.28215e-08 0 3.30185e-08 0 3.302e-08 0.0041358 3.30215e-08 0 3.32185e-08 0 3.322e-08 0.0041358 3.32215e-08 0 3.34185e-08 0 3.342e-08 0.0041358 3.34215e-08 0 3.36185e-08 0 3.362e-08 0.0041358 3.36215e-08 0 3.38185e-08 0 3.382e-08 0.0041358 3.38215e-08 0 3.40185e-08 0 3.402e-08 0.0041358 3.40215e-08 0 3.42185e-08 0 3.422e-08 0.0041358 3.42215e-08 0 3.44185e-08 0 3.442e-08 0.0041358 3.44215e-08 0 3.46185e-08 0 3.462e-08 0.0041358 3.46215e-08 0 3.48185e-08 0 3.482e-08 0.0041358 3.48215e-08 0 3.50185e-08 0 3.502e-08 0.0041358 3.50215e-08 0 3.52185e-08 0 3.522e-08 0.0041358 3.52215e-08 0 3.54185e-08 0 3.542e-08 0.0041358 3.54215e-08 0 3.56185e-08 0 3.562e-08 0.0041358 3.56215e-08 0 3.58185e-08 0 3.582e-08 0.0041358 3.58215e-08 0 3.60185e-08 0 3.602e-08 0.0041358 3.60215e-08 0 3.62185e-08 0 3.622e-08 0.0041358 3.62215e-08 0 3.64185e-08 0 3.642e-08 0.0041358 3.64215e-08 0 3.66185e-08 0 3.662e-08 0.0041358 3.66215e-08 0 3.68185e-08 0 3.682e-08 0.0041358 3.68215e-08 0 3.70185e-08 0 3.702e-08 0.0041358 3.70215e-08 0 3.72185e-08 0 3.722e-08 0.0041358 3.72215e-08 0 3.74185e-08 0 3.742e-08 0.0041358 3.74215e-08 0 3.76185e-08 0 3.762e-08 0.0041358 3.76215e-08 0 3.78185e-08 0 3.782e-08 0.0041358 3.78215e-08 0 3.80185e-08 0 3.802e-08 0.0041358 3.80215e-08 0 3.82185e-08 0 3.822e-08 0.0041358 3.82215e-08 0 3.84185e-08 0 3.842e-08 0.0041358 3.84215e-08 0 3.86185e-08 0 3.862e-08 0.0041358 3.86215e-08 0 3.88185e-08 0 3.882e-08 0.0041358 3.88215e-08 0 3.90185e-08 0 3.902e-08 0.0041358 3.90215e-08 0 3.92185e-08 0 3.922e-08 0.0041358 3.92215e-08 0 3.94185e-08 0 3.942e-08 0.0041358 3.94215e-08 0 3.96185e-08 0 3.962e-08 0.0041358 3.96215e-08 0 3.98185e-08 0 3.982e-08 0.0041358 3.98215e-08 0 4.00185e-08 0 4.002e-08 0.0041358 4.00215e-08 0 4.02185e-08 0 4.022e-08 0.0041358 4.02215e-08 0 4.04185e-08 0 4.042e-08 0.0041358 4.04215e-08 0 4.06185e-08 0 4.062e-08 0.0041358 4.06215e-08 0 4.08185e-08 0 4.082e-08 0.0041358 4.08215e-08 0 4.10185e-08 0 4.102e-08 0.0041358 4.10215e-08 0 4.12185e-08 0 4.122e-08 0.0041358 4.12215e-08 0 4.14185e-08 0 4.142e-08 0.0041358 4.14215e-08 0 4.16185e-08 0 4.162e-08 0.0041358 4.16215e-08 0 4.18185e-08 0 4.182e-08 0.0041358 4.18215e-08 0 4.20185e-08 0 4.202e-08 0.0041358 4.20215e-08 0 4.22185e-08 0 4.222e-08 0.0041358 4.22215e-08 0 4.24185e-08 0 4.242e-08 0.0041358 4.24215e-08 0 4.26185e-08 0 4.262e-08 0.0041358 4.26215e-08 0 4.28185e-08 0 4.282e-08 0.0041358 4.28215e-08 0 4.30185e-08 0 4.302e-08 0.0041358 4.30215e-08 0 4.32185e-08 0 4.322e-08 0.0041358 4.32215e-08 0 4.34185e-08 0 4.342e-08 0.0041358 4.34215e-08 0 4.36185e-08 0 4.362e-08 0.0041358 4.36215e-08 0 4.38185e-08 0 4.382e-08 0.0041358 4.38215e-08 0 4.40185e-08 0 4.402e-08 0.0041358 4.40215e-08 0 4.42185e-08 0 4.422e-08 0.0041358 4.42215e-08 0 4.44185e-08 0 4.442e-08 0.0041358 4.44215e-08 0 4.46185e-08 0 4.462e-08 0.0041358 4.46215e-08 0 4.48185e-08 0 4.482e-08 0.0041358 4.48215e-08 0 4.50185e-08 0 4.502e-08 0.0041358 4.50215e-08 0 4.52185e-08 0 4.522e-08 0.0041358 4.52215e-08 0 4.54185e-08 0 4.542e-08 0.0041358 4.54215e-08 0 4.56185e-08 0 4.562e-08 0.0041358 4.56215e-08 0 4.58185e-08 0 4.582e-08 0.0041358 4.58215e-08 0 4.60185e-08 0 4.602e-08 0.0041358 4.60215e-08 0 4.62185e-08 0 4.622e-08 0.0041358 4.62215e-08 0 4.64185e-08 0 4.642e-08 0.0041358 4.64215e-08 0 4.66185e-08 0 4.662e-08 0.0041358 4.66215e-08 0 4.68185e-08 0 4.682e-08 0.0041358 4.68215e-08 0 4.70185e-08 0 4.702e-08 0.0041358 4.70215e-08 0 4.72185e-08 0 4.722e-08 0.0041358 4.72215e-08 0 4.74185e-08 0 4.742e-08 0.0041358 4.74215e-08 0 4.76185e-08 0 4.762e-08 0.0041358 4.76215e-08 0 4.78185e-08 0 4.782e-08 0.0041358 4.78215e-08 0 4.80185e-08 0 4.802e-08 0.0041358 4.80215e-08 0 4.82185e-08 0 4.822e-08 0.0041358 4.82215e-08 0 4.84185e-08 0 4.842e-08 0.0041358 4.84215e-08 0 4.86185e-08 0 4.862e-08 0.0041358 4.86215e-08 0 4.88185e-08 0 4.882e-08 0.0041358 4.88215e-08 0 4.90185e-08 0 4.902e-08 0.0041358 4.90215e-08 0 4.92185e-08 0 4.922e-08 0.0041358 4.92215e-08 0 4.94185e-08 0 4.942e-08 0.0041358 4.94215e-08 0 4.96185e-08 0 4.962e-08 0.0041358 4.96215e-08 0 4.98185e-08 0 4.982e-08 0.0041358 4.98215e-08 0 5.00185e-08 0 5.002e-08 0.0041358 5.00215e-08 0 5.02185e-08 0 5.022e-08 0.0041358 5.02215e-08 0 5.04185e-08 0 5.042e-08 0.0041358 5.04215e-08 0 5.06185e-08 0 5.062e-08 0.0041358 5.06215e-08 0 5.08185e-08 0 5.082e-08 0.0041358 5.08215e-08 0 5.10185e-08 0 5.102e-08 0.0041358 5.10215e-08 0)
IT03_|T 0 T03_  PWL(0 0 1.85e-11 0 2e-11 0.0041358 2.15e-11 0 2.185e-10 0 2.2e-10 0.0041358 2.215e-10 0 4.185e-10 0 4.2e-10 0.0041358 4.215e-10 0 6.185e-10 0 6.2e-10 0.0041358 6.215e-10 0 8.185e-10 0 8.2e-10 0.0041358 8.215e-10 0 1.0185e-09 0 1.02e-09 0.0041358 1.0215e-09 0 1.2185e-09 0 1.22e-09 0.0041358 1.2215e-09 0 1.4185e-09 0 1.42e-09 0.0041358 1.4215e-09 0 1.6185e-09 0 1.62e-09 0.0041358 1.6215e-09 0 1.8185e-09 0 1.82e-09 0.0041358 1.8215e-09 0 2.0185e-09 0 2.02e-09 0.0041358 2.0215e-09 0 2.2185e-09 0 2.22e-09 0.0041358 2.2215e-09 0 2.4185e-09 0 2.42e-09 0.0041358 2.4215e-09 0 2.6185e-09 0 2.62e-09 0.0041358 2.6215e-09 0 2.8185e-09 0 2.82e-09 0.0041358 2.8215e-09 0 3.0185e-09 0 3.02e-09 0.0041358 3.0215e-09 0 3.2185e-09 0 3.22e-09 0.0041358 3.2215e-09 0 3.4185e-09 0 3.42e-09 0.0041358 3.4215e-09 0 3.6185e-09 0 3.62e-09 0.0041358 3.6215e-09 0 3.8185e-09 0 3.82e-09 0.0041358 3.8215e-09 0 4.0185e-09 0 4.02e-09 0.0041358 4.0215e-09 0 4.2185e-09 0 4.22e-09 0.0041358 4.2215e-09 0 4.4185e-09 0 4.42e-09 0.0041358 4.4215e-09 0 4.6185e-09 0 4.62e-09 0.0041358 4.6215e-09 0 4.8185e-09 0 4.82e-09 0.0041358 4.8215e-09 0 5.0185e-09 0 5.02e-09 0.0041358 5.0215e-09 0 5.2185e-09 0 5.22e-09 0.0041358 5.2215e-09 0 5.4185e-09 0 5.42e-09 0.0041358 5.4215e-09 0 5.6185e-09 0 5.62e-09 0.0041358 5.6215e-09 0 5.8185e-09 0 5.82e-09 0.0041358 5.8215e-09 0 6.0185e-09 0 6.02e-09 0.0041358 6.0215e-09 0 6.2185e-09 0 6.22e-09 0.0041358 6.2215e-09 0 6.4185e-09 0 6.42e-09 0.0041358 6.4215e-09 0 6.6185e-09 0 6.62e-09 0.0041358 6.6215e-09 0 6.8185e-09 0 6.82e-09 0.0041358 6.8215e-09 0 7.0185e-09 0 7.02e-09 0.0041358 7.0215e-09 0 7.2185e-09 0 7.22e-09 0.0041358 7.2215e-09 0 7.4185e-09 0 7.42e-09 0.0041358 7.4215e-09 0 7.6185e-09 0 7.62e-09 0.0041358 7.6215e-09 0 7.8185e-09 0 7.82e-09 0.0041358 7.8215e-09 0 8.0185e-09 0 8.02e-09 0.0041358 8.0215e-09 0 8.2185e-09 0 8.22e-09 0.0041358 8.2215e-09 0 8.4185e-09 0 8.42e-09 0.0041358 8.4215e-09 0 8.6185e-09 0 8.62e-09 0.0041358 8.6215e-09 0 8.8185e-09 0 8.82e-09 0.0041358 8.8215e-09 0 9.0185e-09 0 9.02e-09 0.0041358 9.0215e-09 0 9.2185e-09 0 9.22e-09 0.0041358 9.2215e-09 0 9.4185e-09 0 9.42e-09 0.0041358 9.4215e-09 0 9.6185e-09 0 9.62e-09 0.0041358 9.6215e-09 0 9.8185e-09 0 9.82e-09 0.0041358 9.8215e-09 0 1.00185e-08 0 1.002e-08 0.0041358 1.00215e-08 0 1.02185e-08 0 1.022e-08 0.0041358 1.02215e-08 0 1.04185e-08 0 1.042e-08 0.0041358 1.04215e-08 0 1.06185e-08 0 1.062e-08 0.0041358 1.06215e-08 0 1.08185e-08 0 1.082e-08 0.0041358 1.08215e-08 0 1.10185e-08 0 1.102e-08 0.0041358 1.10215e-08 0 1.12185e-08 0 1.122e-08 0.0041358 1.12215e-08 0 1.14185e-08 0 1.142e-08 0.0041358 1.14215e-08 0 1.16185e-08 0 1.162e-08 0.0041358 1.16215e-08 0 1.18185e-08 0 1.182e-08 0.0041358 1.18215e-08 0 1.20185e-08 0 1.202e-08 0.0041358 1.20215e-08 0 1.22185e-08 0 1.222e-08 0.0041358 1.22215e-08 0 1.24185e-08 0 1.242e-08 0.0041358 1.24215e-08 0 1.26185e-08 0 1.262e-08 0.0041358 1.26215e-08 0 1.28185e-08 0 1.282e-08 0.0041358 1.28215e-08 0 1.30185e-08 0 1.302e-08 0.0041358 1.30215e-08 0 1.32185e-08 0 1.322e-08 0.0041358 1.32215e-08 0 1.34185e-08 0 1.342e-08 0.0041358 1.34215e-08 0 1.36185e-08 0 1.362e-08 0.0041358 1.36215e-08 0 1.38185e-08 0 1.382e-08 0.0041358 1.38215e-08 0 1.40185e-08 0 1.402e-08 0.0041358 1.40215e-08 0 1.42185e-08 0 1.422e-08 0.0041358 1.42215e-08 0 1.44185e-08 0 1.442e-08 0.0041358 1.44215e-08 0 1.46185e-08 0 1.462e-08 0.0041358 1.46215e-08 0 1.48185e-08 0 1.482e-08 0.0041358 1.48215e-08 0 1.50185e-08 0 1.502e-08 0.0041358 1.50215e-08 0 1.52185e-08 0 1.522e-08 0.0041358 1.52215e-08 0 1.54185e-08 0 1.542e-08 0.0041358 1.54215e-08 0 1.56185e-08 0 1.562e-08 0.0041358 1.56215e-08 0 1.58185e-08 0 1.582e-08 0.0041358 1.58215e-08 0 1.60185e-08 0 1.602e-08 0.0041358 1.60215e-08 0 1.62185e-08 0 1.622e-08 0.0041358 1.62215e-08 0 1.64185e-08 0 1.642e-08 0.0041358 1.64215e-08 0 1.66185e-08 0 1.662e-08 0.0041358 1.66215e-08 0 1.68185e-08 0 1.682e-08 0.0041358 1.68215e-08 0 1.70185e-08 0 1.702e-08 0.0041358 1.70215e-08 0 1.72185e-08 0 1.722e-08 0.0041358 1.72215e-08 0 1.74185e-08 0 1.742e-08 0.0041358 1.74215e-08 0 1.76185e-08 0 1.762e-08 0.0041358 1.76215e-08 0 1.78185e-08 0 1.782e-08 0.0041358 1.78215e-08 0 1.80185e-08 0 1.802e-08 0.0041358 1.80215e-08 0 1.82185e-08 0 1.822e-08 0.0041358 1.82215e-08 0 1.84185e-08 0 1.842e-08 0.0041358 1.84215e-08 0 1.86185e-08 0 1.862e-08 0.0041358 1.86215e-08 0 1.88185e-08 0 1.882e-08 0.0041358 1.88215e-08 0 1.90185e-08 0 1.902e-08 0.0041358 1.90215e-08 0 1.92185e-08 0 1.922e-08 0.0041358 1.92215e-08 0 1.94185e-08 0 1.942e-08 0.0041358 1.94215e-08 0 1.96185e-08 0 1.962e-08 0.0041358 1.96215e-08 0 1.98185e-08 0 1.982e-08 0.0041358 1.98215e-08 0 2.00185e-08 0 2.002e-08 0.0041358 2.00215e-08 0 2.02185e-08 0 2.022e-08 0.0041358 2.02215e-08 0 2.04185e-08 0 2.042e-08 0.0041358 2.04215e-08 0 2.06185e-08 0 2.062e-08 0.0041358 2.06215e-08 0 2.08185e-08 0 2.082e-08 0.0041358 2.08215e-08 0 2.10185e-08 0 2.102e-08 0.0041358 2.10215e-08 0 2.12185e-08 0 2.122e-08 0.0041358 2.12215e-08 0 2.14185e-08 0 2.142e-08 0.0041358 2.14215e-08 0 2.16185e-08 0 2.162e-08 0.0041358 2.16215e-08 0 2.18185e-08 0 2.182e-08 0.0041358 2.18215e-08 0 2.20185e-08 0 2.202e-08 0.0041358 2.20215e-08 0 2.22185e-08 0 2.222e-08 0.0041358 2.22215e-08 0 2.24185e-08 0 2.242e-08 0.0041358 2.24215e-08 0 2.26185e-08 0 2.262e-08 0.0041358 2.26215e-08 0 2.28185e-08 0 2.282e-08 0.0041358 2.28215e-08 0 2.30185e-08 0 2.302e-08 0.0041358 2.30215e-08 0 2.32185e-08 0 2.322e-08 0.0041358 2.32215e-08 0 2.34185e-08 0 2.342e-08 0.0041358 2.34215e-08 0 2.36185e-08 0 2.362e-08 0.0041358 2.36215e-08 0 2.38185e-08 0 2.382e-08 0.0041358 2.38215e-08 0 2.40185e-08 0 2.402e-08 0.0041358 2.40215e-08 0 2.42185e-08 0 2.422e-08 0.0041358 2.42215e-08 0 2.44185e-08 0 2.442e-08 0.0041358 2.44215e-08 0 2.46185e-08 0 2.462e-08 0.0041358 2.46215e-08 0 2.48185e-08 0 2.482e-08 0.0041358 2.48215e-08 0 2.50185e-08 0 2.502e-08 0.0041358 2.50215e-08 0 2.52185e-08 0 2.522e-08 0.0041358 2.52215e-08 0 2.54185e-08 0 2.542e-08 0.0041358 2.54215e-08 0 2.56185e-08 0 2.562e-08 0.0041358 2.56215e-08 0 2.58185e-08 0 2.582e-08 0.0041358 2.58215e-08 0 2.60185e-08 0 2.602e-08 0.0041358 2.60215e-08 0 2.62185e-08 0 2.622e-08 0.0041358 2.62215e-08 0 2.64185e-08 0 2.642e-08 0.0041358 2.64215e-08 0 2.66185e-08 0 2.662e-08 0.0041358 2.66215e-08 0 2.68185e-08 0 2.682e-08 0.0041358 2.68215e-08 0 2.70185e-08 0 2.702e-08 0.0041358 2.70215e-08 0 2.72185e-08 0 2.722e-08 0.0041358 2.72215e-08 0 2.74185e-08 0 2.742e-08 0.0041358 2.74215e-08 0 2.76185e-08 0 2.762e-08 0.0041358 2.76215e-08 0 2.78185e-08 0 2.782e-08 0.0041358 2.78215e-08 0 2.80185e-08 0 2.802e-08 0.0041358 2.80215e-08 0 2.82185e-08 0 2.822e-08 0.0041358 2.82215e-08 0 2.84185e-08 0 2.842e-08 0.0041358 2.84215e-08 0 2.86185e-08 0 2.862e-08 0.0041358 2.86215e-08 0 2.88185e-08 0 2.882e-08 0.0041358 2.88215e-08 0 2.90185e-08 0 2.902e-08 0.0041358 2.90215e-08 0 2.92185e-08 0 2.922e-08 0.0041358 2.92215e-08 0 2.94185e-08 0 2.942e-08 0.0041358 2.94215e-08 0 2.96185e-08 0 2.962e-08 0.0041358 2.96215e-08 0 2.98185e-08 0 2.982e-08 0.0041358 2.98215e-08 0 3.00185e-08 0 3.002e-08 0.0041358 3.00215e-08 0 3.02185e-08 0 3.022e-08 0.0041358 3.02215e-08 0 3.04185e-08 0 3.042e-08 0.0041358 3.04215e-08 0 3.06185e-08 0 3.062e-08 0.0041358 3.06215e-08 0 3.08185e-08 0 3.082e-08 0.0041358 3.08215e-08 0 3.10185e-08 0 3.102e-08 0.0041358 3.10215e-08 0 3.12185e-08 0 3.122e-08 0.0041358 3.12215e-08 0 3.14185e-08 0 3.142e-08 0.0041358 3.14215e-08 0 3.16185e-08 0 3.162e-08 0.0041358 3.16215e-08 0 3.18185e-08 0 3.182e-08 0.0041358 3.18215e-08 0 3.20185e-08 0 3.202e-08 0.0041358 3.20215e-08 0 3.22185e-08 0 3.222e-08 0.0041358 3.22215e-08 0 3.24185e-08 0 3.242e-08 0.0041358 3.24215e-08 0 3.26185e-08 0 3.262e-08 0.0041358 3.26215e-08 0 3.28185e-08 0 3.282e-08 0.0041358 3.28215e-08 0 3.30185e-08 0 3.302e-08 0.0041358 3.30215e-08 0 3.32185e-08 0 3.322e-08 0.0041358 3.32215e-08 0 3.34185e-08 0 3.342e-08 0.0041358 3.34215e-08 0 3.36185e-08 0 3.362e-08 0.0041358 3.36215e-08 0 3.38185e-08 0 3.382e-08 0.0041358 3.38215e-08 0 3.40185e-08 0 3.402e-08 0.0041358 3.40215e-08 0 3.42185e-08 0 3.422e-08 0.0041358 3.42215e-08 0 3.44185e-08 0 3.442e-08 0.0041358 3.44215e-08 0 3.46185e-08 0 3.462e-08 0.0041358 3.46215e-08 0 3.48185e-08 0 3.482e-08 0.0041358 3.48215e-08 0 3.50185e-08 0 3.502e-08 0.0041358 3.50215e-08 0 3.52185e-08 0 3.522e-08 0.0041358 3.52215e-08 0 3.54185e-08 0 3.542e-08 0.0041358 3.54215e-08 0 3.56185e-08 0 3.562e-08 0.0041358 3.56215e-08 0 3.58185e-08 0 3.582e-08 0.0041358 3.58215e-08 0 3.60185e-08 0 3.602e-08 0.0041358 3.60215e-08 0 3.62185e-08 0 3.622e-08 0.0041358 3.62215e-08 0 3.64185e-08 0 3.642e-08 0.0041358 3.64215e-08 0 3.66185e-08 0 3.662e-08 0.0041358 3.66215e-08 0 3.68185e-08 0 3.682e-08 0.0041358 3.68215e-08 0 3.70185e-08 0 3.702e-08 0.0041358 3.70215e-08 0 3.72185e-08 0 3.722e-08 0.0041358 3.72215e-08 0 3.74185e-08 0 3.742e-08 0.0041358 3.74215e-08 0 3.76185e-08 0 3.762e-08 0.0041358 3.76215e-08 0 3.78185e-08 0 3.782e-08 0.0041358 3.78215e-08 0 3.80185e-08 0 3.802e-08 0.0041358 3.80215e-08 0 3.82185e-08 0 3.822e-08 0.0041358 3.82215e-08 0 3.84185e-08 0 3.842e-08 0.0041358 3.84215e-08 0 3.86185e-08 0 3.862e-08 0.0041358 3.86215e-08 0 3.88185e-08 0 3.882e-08 0.0041358 3.88215e-08 0 3.90185e-08 0 3.902e-08 0.0041358 3.90215e-08 0 3.92185e-08 0 3.922e-08 0.0041358 3.92215e-08 0 3.94185e-08 0 3.942e-08 0.0041358 3.94215e-08 0 3.96185e-08 0 3.962e-08 0.0041358 3.96215e-08 0 3.98185e-08 0 3.982e-08 0.0041358 3.98215e-08 0 4.00185e-08 0 4.002e-08 0.0041358 4.00215e-08 0 4.02185e-08 0 4.022e-08 0.0041358 4.02215e-08 0 4.04185e-08 0 4.042e-08 0.0041358 4.04215e-08 0 4.06185e-08 0 4.062e-08 0.0041358 4.06215e-08 0 4.08185e-08 0 4.082e-08 0.0041358 4.08215e-08 0 4.10185e-08 0 4.102e-08 0.0041358 4.10215e-08 0 4.12185e-08 0 4.122e-08 0.0041358 4.12215e-08 0 4.14185e-08 0 4.142e-08 0.0041358 4.14215e-08 0 4.16185e-08 0 4.162e-08 0.0041358 4.16215e-08 0 4.18185e-08 0 4.182e-08 0.0041358 4.18215e-08 0 4.20185e-08 0 4.202e-08 0.0041358 4.20215e-08 0 4.22185e-08 0 4.222e-08 0.0041358 4.22215e-08 0 4.24185e-08 0 4.242e-08 0.0041358 4.24215e-08 0 4.26185e-08 0 4.262e-08 0.0041358 4.26215e-08 0 4.28185e-08 0 4.282e-08 0.0041358 4.28215e-08 0 4.30185e-08 0 4.302e-08 0.0041358 4.30215e-08 0 4.32185e-08 0 4.322e-08 0.0041358 4.32215e-08 0 4.34185e-08 0 4.342e-08 0.0041358 4.34215e-08 0 4.36185e-08 0 4.362e-08 0.0041358 4.36215e-08 0 4.38185e-08 0 4.382e-08 0.0041358 4.38215e-08 0 4.40185e-08 0 4.402e-08 0.0041358 4.40215e-08 0 4.42185e-08 0 4.422e-08 0.0041358 4.42215e-08 0 4.44185e-08 0 4.442e-08 0.0041358 4.44215e-08 0 4.46185e-08 0 4.462e-08 0.0041358 4.46215e-08 0 4.48185e-08 0 4.482e-08 0.0041358 4.48215e-08 0 4.50185e-08 0 4.502e-08 0.0041358 4.50215e-08 0 4.52185e-08 0 4.522e-08 0.0041358 4.52215e-08 0 4.54185e-08 0 4.542e-08 0.0041358 4.54215e-08 0 4.56185e-08 0 4.562e-08 0.0041358 4.56215e-08 0 4.58185e-08 0 4.582e-08 0.0041358 4.58215e-08 0 4.60185e-08 0 4.602e-08 0.0041358 4.60215e-08 0 4.62185e-08 0 4.622e-08 0.0041358 4.62215e-08 0 4.64185e-08 0 4.642e-08 0.0041358 4.64215e-08 0 4.66185e-08 0 4.662e-08 0.0041358 4.66215e-08 0 4.68185e-08 0 4.682e-08 0.0041358 4.68215e-08 0 4.70185e-08 0 4.702e-08 0.0041358 4.70215e-08 0 4.72185e-08 0 4.722e-08 0.0041358 4.72215e-08 0 4.74185e-08 0 4.742e-08 0.0041358 4.74215e-08 0 4.76185e-08 0 4.762e-08 0.0041358 4.76215e-08 0 4.78185e-08 0 4.782e-08 0.0041358 4.78215e-08 0 4.80185e-08 0 4.802e-08 0.0041358 4.80215e-08 0 4.82185e-08 0 4.822e-08 0.0041358 4.82215e-08 0 4.84185e-08 0 4.842e-08 0.0041358 4.84215e-08 0 4.86185e-08 0 4.862e-08 0.0041358 4.86215e-08 0 4.88185e-08 0 4.882e-08 0.0041358 4.88215e-08 0 4.90185e-08 0 4.902e-08 0.0041358 4.90215e-08 0 4.92185e-08 0 4.922e-08 0.0041358 4.92215e-08 0 4.94185e-08 0 4.942e-08 0.0041358 4.94215e-08 0 4.96185e-08 0 4.962e-08 0.0041358 4.96215e-08 0 4.98185e-08 0 4.982e-08 0.0041358 4.98215e-08 0 5.00185e-08 0 5.002e-08 0.0041358 5.00215e-08 0 5.02185e-08 0 5.022e-08 0.0041358 5.02215e-08 0 5.04185e-08 0 5.042e-08 0.0041358 5.04215e-08 0 5.06185e-08 0 5.062e-08 0.0041358 5.06215e-08 0 5.08185e-08 0 5.082e-08 0.0041358 5.08215e-08 0 5.10185e-08 0 5.102e-08 0.0041358 5.10215e-08 0)
LSPL_IG0_0_|1 IG0_0_ SPL_IG0_0_|D1  2e-12
LSPL_IG0_0_|2 SPL_IG0_0_|D1 SPL_IG0_0_|D2  4.135667696e-12
LSPL_IG0_0_|3 SPL_IG0_0_|D2 SPL_IG0_0_|JCT  9.84682784761905e-13
LSPL_IG0_0_|4 SPL_IG0_0_|JCT SPL_IG0_0_|QA1  9.84682784761905e-13
LSPL_IG0_0_|5 SPL_IG0_0_|QA1 IG0_0_TO0_  2e-12
LSPL_IG0_0_|6 SPL_IG0_0_|JCT SPL_IG0_0_|QB1  9.84682784761905e-13
LSPL_IG0_0_|7 SPL_IG0_0_|QB1 IG0_0_TO1_  2e-12
LSPL_IP1_0_|1 IP1_0_ SPL_IP1_0_|D1  2e-12
LSPL_IP1_0_|2 SPL_IP1_0_|D1 SPL_IP1_0_|D2  4.135667696e-12
LSPL_IP1_0_|3 SPL_IP1_0_|D2 SPL_IP1_0_|JCT  9.84682784761905e-13
LSPL_IP1_0_|4 SPL_IP1_0_|JCT SPL_IP1_0_|QA1  9.84682784761905e-13
LSPL_IP1_0_|5 SPL_IP1_0_|QA1 IP1_0_TO1_  2e-12
LSPL_IP1_0_|6 SPL_IP1_0_|JCT SPL_IP1_0_|QB1  9.84682784761905e-13
LSPL_IP1_0_|7 SPL_IP1_0_|QB1 IP1_0_OUT_  2e-12
LSPL_IG2_0_|1 IG2_0_ SPL_IG2_0_|D1  2e-12
LSPL_IG2_0_|2 SPL_IG2_0_|D1 SPL_IG2_0_|D2  4.135667696e-12
LSPL_IG2_0_|3 SPL_IG2_0_|D2 SPL_IG2_0_|JCT  9.84682784761905e-13
LSPL_IG2_0_|4 SPL_IG2_0_|JCT SPL_IG2_0_|QA1  9.84682784761905e-13
LSPL_IG2_0_|5 SPL_IG2_0_|QA1 IG2_0_TO2_  2e-12
LSPL_IG2_0_|6 SPL_IG2_0_|JCT SPL_IG2_0_|QB1  9.84682784761905e-13
LSPL_IG2_0_|7 SPL_IG2_0_|QB1 IG2_0_TO3_  2e-12
LSPL_IP3_0_|1 IP3_0_ SPL_IP3_0_|D1  2e-12
LSPL_IP3_0_|2 SPL_IP3_0_|D1 SPL_IP3_0_|D2  4.135667696e-12
LSPL_IP3_0_|3 SPL_IP3_0_|D2 SPL_IP3_0_|JCT  9.84682784761905e-13
LSPL_IP3_0_|4 SPL_IP3_0_|JCT SPL_IP3_0_|QA1  9.84682784761905e-13
LSPL_IP3_0_|5 SPL_IP3_0_|QA1 IP3_0_TO1_  2e-12
LSPL_IP3_0_|6 SPL_IP3_0_|JCT SPL_IP3_0_|QB1  9.84682784761905e-13
LSPL_IP3_0_|7 SPL_IP3_0_|QB1 IP3_0_OUT_  2e-12
IT04_|T 0 T04_  PWL(0 0 1.35e-11 0 1.5e-11 0.0027572 1.65e-11 0 2.135e-10 0 2.15e-10 0.0027572 2.165e-10 0 4.135e-10 0 4.15e-10 0.0027572 4.165e-10 0 6.135e-10 0 6.15e-10 0.0027572 6.165e-10 0 8.135e-10 0 8.15e-10 0.0027572 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0027572 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0027572 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0027572 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0027572 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0027572 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0027572 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0027572 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0027572 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0027572 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0027572 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0027572 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0027572 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0027572 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0027572 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0027572 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0027572 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0027572 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0027572 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0027572 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0027572 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0027572 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0027572 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0027572 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0027572 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0027572 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0027572 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0027572 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0027572 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0027572 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0027572 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0027572 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0027572 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0027572 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0027572 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0027572 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0027572 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0027572 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0027572 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0027572 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0027572 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0027572 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0027572 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0027572 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0027572 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0027572 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0027572 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0027572 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0027572 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0027572 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0027572 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0027572 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0027572 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0027572 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0027572 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0027572 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0027572 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0027572 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0027572 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0027572 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0027572 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0027572 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0027572 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0027572 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0027572 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0027572 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0027572 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0027572 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0027572 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0027572 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0027572 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0027572 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0027572 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0027572 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0027572 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0027572 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0027572 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0027572 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0027572 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0027572 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0027572 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0027572 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0027572 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0027572 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0027572 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0027572 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0027572 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0027572 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0027572 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0027572 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0027572 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0027572 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0027572 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0027572 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0027572 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0027572 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0027572 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0027572 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0027572 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0027572 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0027572 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0027572 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0027572 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0027572 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0027572 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0027572 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0027572 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0027572 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0027572 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0027572 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0027572 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0027572 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0027572 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0027572 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0027572 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0027572 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0027572 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0027572 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0027572 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0027572 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0027572 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0027572 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0027572 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0027572 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0027572 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0027572 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0027572 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0027572 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0027572 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0027572 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0027572 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0027572 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0027572 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0027572 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0027572 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0027572 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0027572 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0027572 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0027572 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0027572 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0027572 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0027572 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0027572 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0027572 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0027572 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0027572 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0027572 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0027572 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0027572 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0027572 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0027572 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0027572 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0027572 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0027572 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0027572 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0027572 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0027572 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0027572 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0027572 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0027572 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0027572 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0027572 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0027572 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0027572 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0027572 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0027572 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0027572 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0027572 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0027572 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0027572 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0027572 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0027572 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0027572 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0027572 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0027572 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0027572 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0027572 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0027572 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0027572 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0027572 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0027572 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0027572 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0027572 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0027572 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0027572 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0027572 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0027572 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0027572 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0027572 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0027572 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0027572 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0027572 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0027572 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0027572 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0027572 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0027572 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0027572 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0027572 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0027572 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0027572 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0027572 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0027572 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0027572 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0027572 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0027572 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0027572 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0027572 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0027572 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0027572 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0027572 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0027572 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0027572 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0027572 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0027572 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0027572 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0027572 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0027572 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0027572 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0027572 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0027572 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0027572 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0027572 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0027572 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0027572 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0027572 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0027572 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0027572 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0027572 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0027572 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0027572 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0027572 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0027572 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0027572 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0027572 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0027572 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0027572 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0027572 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0027572 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0027572 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0027572 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0027572 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0027572 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0027572 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0027572 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0027572 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0027572 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0027572 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0027572 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0027572 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0027572 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0027572 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0027572 5.10165e-08 0)
IT05_|T 0 T05_  PWL(0 0 1.35e-11 0 1.5e-11 0.0027572 1.65e-11 0 2.135e-10 0 2.15e-10 0.0027572 2.165e-10 0 4.135e-10 0 4.15e-10 0.0027572 4.165e-10 0 6.135e-10 0 6.15e-10 0.0027572 6.165e-10 0 8.135e-10 0 8.15e-10 0.0027572 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0027572 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0027572 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0027572 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0027572 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0027572 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0027572 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0027572 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0027572 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0027572 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0027572 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0027572 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0027572 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0027572 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0027572 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0027572 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0027572 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0027572 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0027572 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0027572 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0027572 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0027572 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0027572 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0027572 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0027572 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0027572 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0027572 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0027572 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0027572 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0027572 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0027572 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0027572 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0027572 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0027572 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0027572 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0027572 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0027572 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0027572 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0027572 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0027572 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0027572 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0027572 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0027572 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0027572 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0027572 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0027572 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0027572 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0027572 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0027572 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0027572 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0027572 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0027572 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0027572 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0027572 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0027572 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0027572 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0027572 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0027572 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0027572 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0027572 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0027572 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0027572 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0027572 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0027572 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0027572 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0027572 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0027572 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0027572 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0027572 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0027572 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0027572 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0027572 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0027572 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0027572 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0027572 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0027572 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0027572 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0027572 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0027572 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0027572 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0027572 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0027572 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0027572 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0027572 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0027572 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0027572 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0027572 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0027572 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0027572 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0027572 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0027572 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0027572 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0027572 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0027572 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0027572 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0027572 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0027572 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0027572 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0027572 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0027572 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0027572 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0027572 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0027572 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0027572 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0027572 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0027572 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0027572 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0027572 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0027572 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0027572 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0027572 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0027572 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0027572 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0027572 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0027572 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0027572 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0027572 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0027572 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0027572 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0027572 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0027572 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0027572 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0027572 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0027572 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0027572 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0027572 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0027572 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0027572 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0027572 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0027572 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0027572 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0027572 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0027572 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0027572 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0027572 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0027572 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0027572 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0027572 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0027572 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0027572 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0027572 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0027572 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0027572 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0027572 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0027572 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0027572 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0027572 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0027572 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0027572 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0027572 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0027572 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0027572 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0027572 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0027572 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0027572 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0027572 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0027572 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0027572 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0027572 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0027572 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0027572 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0027572 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0027572 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0027572 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0027572 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0027572 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0027572 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0027572 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0027572 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0027572 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0027572 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0027572 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0027572 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0027572 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0027572 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0027572 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0027572 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0027572 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0027572 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0027572 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0027572 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0027572 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0027572 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0027572 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0027572 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0027572 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0027572 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0027572 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0027572 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0027572 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0027572 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0027572 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0027572 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0027572 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0027572 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0027572 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0027572 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0027572 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0027572 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0027572 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0027572 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0027572 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0027572 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0027572 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0027572 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0027572 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0027572 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0027572 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0027572 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0027572 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0027572 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0027572 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0027572 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0027572 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0027572 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0027572 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0027572 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0027572 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0027572 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0027572 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0027572 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0027572 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0027572 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0027572 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0027572 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0027572 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0027572 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0027572 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0027572 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0027572 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0027572 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0027572 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0027572 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0027572 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0027572 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0027572 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0027572 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0027572 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0027572 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0027572 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0027572 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0027572 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0027572 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0027572 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0027572 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0027572 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0027572 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0027572 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0027572 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0027572 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0027572 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0027572 5.10165e-08 0)
IT06_|T 0 T06_  PWL(0 0 1.35e-11 0 1.5e-11 0.0027572 1.65e-11 0 2.135e-10 0 2.15e-10 0.0027572 2.165e-10 0 4.135e-10 0 4.15e-10 0.0027572 4.165e-10 0 6.135e-10 0 6.15e-10 0.0027572 6.165e-10 0 8.135e-10 0 8.15e-10 0.0027572 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0027572 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0027572 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0027572 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0027572 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0027572 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0027572 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0027572 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0027572 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0027572 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0027572 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0027572 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0027572 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0027572 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0027572 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0027572 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0027572 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0027572 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0027572 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0027572 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0027572 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0027572 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0027572 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0027572 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0027572 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0027572 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0027572 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0027572 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0027572 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0027572 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0027572 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0027572 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0027572 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0027572 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0027572 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0027572 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0027572 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0027572 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0027572 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0027572 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0027572 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0027572 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0027572 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0027572 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0027572 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0027572 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0027572 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0027572 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0027572 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0027572 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0027572 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0027572 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0027572 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0027572 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0027572 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0027572 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0027572 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0027572 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0027572 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0027572 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0027572 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0027572 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0027572 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0027572 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0027572 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0027572 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0027572 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0027572 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0027572 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0027572 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0027572 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0027572 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0027572 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0027572 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0027572 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0027572 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0027572 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0027572 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0027572 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0027572 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0027572 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0027572 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0027572 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0027572 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0027572 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0027572 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0027572 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0027572 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0027572 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0027572 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0027572 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0027572 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0027572 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0027572 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0027572 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0027572 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0027572 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0027572 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0027572 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0027572 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0027572 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0027572 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0027572 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0027572 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0027572 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0027572 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0027572 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0027572 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0027572 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0027572 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0027572 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0027572 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0027572 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0027572 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0027572 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0027572 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0027572 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0027572 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0027572 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0027572 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0027572 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0027572 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0027572 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0027572 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0027572 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0027572 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0027572 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0027572 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0027572 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0027572 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0027572 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0027572 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0027572 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0027572 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0027572 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0027572 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0027572 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0027572 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0027572 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0027572 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0027572 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0027572 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0027572 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0027572 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0027572 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0027572 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0027572 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0027572 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0027572 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0027572 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0027572 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0027572 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0027572 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0027572 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0027572 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0027572 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0027572 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0027572 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0027572 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0027572 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0027572 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0027572 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0027572 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0027572 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0027572 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0027572 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0027572 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0027572 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0027572 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0027572 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0027572 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0027572 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0027572 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0027572 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0027572 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0027572 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0027572 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0027572 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0027572 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0027572 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0027572 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0027572 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0027572 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0027572 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0027572 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0027572 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0027572 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0027572 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0027572 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0027572 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0027572 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0027572 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0027572 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0027572 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0027572 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0027572 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0027572 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0027572 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0027572 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0027572 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0027572 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0027572 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0027572 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0027572 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0027572 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0027572 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0027572 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0027572 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0027572 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0027572 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0027572 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0027572 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0027572 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0027572 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0027572 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0027572 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0027572 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0027572 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0027572 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0027572 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0027572 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0027572 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0027572 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0027572 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0027572 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0027572 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0027572 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0027572 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0027572 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0027572 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0027572 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0027572 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0027572 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0027572 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0027572 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0027572 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0027572 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0027572 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0027572 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0027572 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0027572 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0027572 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0027572 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0027572 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0027572 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0027572 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0027572 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0027572 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0027572 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0027572 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0027572 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0027572 5.10165e-08 0)
IT07_|T 0 T07_  PWL(0 0 1.35e-11 0 1.5e-11 0.0055144 1.65e-11 0 2.135e-10 0 2.15e-10 0.0055144 2.165e-10 0 4.135e-10 0 4.15e-10 0.0055144 4.165e-10 0 6.135e-10 0 6.15e-10 0.0055144 6.165e-10 0 8.135e-10 0 8.15e-10 0.0055144 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0055144 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0055144 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0055144 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0055144 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0055144 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0055144 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0055144 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0055144 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0055144 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0055144 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0055144 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0055144 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0055144 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0055144 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0055144 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0055144 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0055144 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0055144 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0055144 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0055144 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0055144 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0055144 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0055144 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0055144 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0055144 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0055144 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0055144 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0055144 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0055144 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0055144 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0055144 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0055144 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0055144 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0055144 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0055144 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0055144 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0055144 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0055144 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0055144 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0055144 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0055144 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0055144 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0055144 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0055144 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0055144 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0055144 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0055144 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0055144 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0055144 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0055144 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0055144 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0055144 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0055144 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0055144 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0055144 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0055144 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0055144 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0055144 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0055144 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0055144 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0055144 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0055144 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0055144 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0055144 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0055144 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0055144 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0055144 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0055144 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0055144 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0055144 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0055144 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0055144 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0055144 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0055144 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0055144 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0055144 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0055144 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0055144 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0055144 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0055144 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0055144 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0055144 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0055144 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0055144 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0055144 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0055144 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0055144 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0055144 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0055144 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0055144 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0055144 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0055144 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0055144 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0055144 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0055144 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0055144 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0055144 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0055144 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0055144 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0055144 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0055144 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0055144 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0055144 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0055144 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0055144 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0055144 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0055144 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0055144 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0055144 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0055144 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0055144 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0055144 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0055144 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0055144 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0055144 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0055144 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0055144 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0055144 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0055144 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0055144 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0055144 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0055144 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0055144 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0055144 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0055144 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0055144 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0055144 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0055144 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0055144 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0055144 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0055144 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0055144 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0055144 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0055144 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0055144 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0055144 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0055144 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0055144 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0055144 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0055144 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0055144 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0055144 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0055144 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0055144 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0055144 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0055144 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0055144 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0055144 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0055144 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0055144 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0055144 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0055144 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0055144 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0055144 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0055144 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0055144 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0055144 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0055144 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0055144 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0055144 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0055144 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0055144 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0055144 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0055144 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0055144 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0055144 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0055144 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0055144 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0055144 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0055144 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0055144 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0055144 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0055144 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0055144 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0055144 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0055144 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0055144 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0055144 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0055144 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0055144 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0055144 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0055144 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0055144 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0055144 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0055144 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0055144 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0055144 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0055144 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0055144 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0055144 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0055144 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0055144 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0055144 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0055144 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0055144 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0055144 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0055144 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0055144 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0055144 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0055144 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0055144 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0055144 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0055144 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0055144 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0055144 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0055144 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0055144 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0055144 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0055144 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0055144 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0055144 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0055144 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0055144 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0055144 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0055144 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0055144 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0055144 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0055144 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0055144 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0055144 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0055144 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0055144 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0055144 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0055144 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0055144 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0055144 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0055144 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0055144 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0055144 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0055144 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0055144 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0055144 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0055144 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0055144 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0055144 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0055144 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0055144 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0055144 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0055144 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0055144 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0055144 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0055144 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0055144 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0055144 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0055144 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0055144 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0055144 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0055144 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0055144 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0055144 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0055144 5.10165e-08 0)
ID01_|T 0 D01_  PWL(0 0 1.35e-11 0 1.5e-11 0.0013786 1.65e-11 0 2.135e-10 0 2.15e-10 0.0013786 2.165e-10 0 4.135e-10 0 4.15e-10 0.0013786 4.165e-10 0 6.135e-10 0 6.15e-10 0.0013786 6.165e-10 0 8.135e-10 0 8.15e-10 0.0013786 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0013786 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0013786 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0013786 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0013786 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0013786 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0013786 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0013786 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0013786 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0013786 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0013786 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0013786 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0013786 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0013786 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0013786 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0013786 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0013786 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0013786 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0013786 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0013786 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0013786 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0013786 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0013786 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0013786 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0013786 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0013786 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0013786 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0013786 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0013786 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0013786 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0013786 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0013786 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0013786 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0013786 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0013786 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0013786 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0013786 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0013786 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0013786 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0013786 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0013786 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0013786 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0013786 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0013786 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0013786 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0013786 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0013786 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0013786 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0013786 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0013786 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0013786 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0013786 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0013786 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0013786 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0013786 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0013786 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0013786 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0013786 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0013786 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0013786 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0013786 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0013786 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0013786 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0013786 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0013786 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0013786 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0013786 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0013786 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0013786 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0013786 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0013786 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0013786 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0013786 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0013786 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0013786 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0013786 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0013786 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0013786 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0013786 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0013786 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0013786 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0013786 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0013786 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0013786 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0013786 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0013786 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0013786 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0013786 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0013786 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0013786 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0013786 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0013786 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0013786 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0013786 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0013786 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0013786 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0013786 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0013786 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0013786 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0013786 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0013786 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0013786 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0013786 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0013786 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0013786 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0013786 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0013786 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0013786 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0013786 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0013786 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0013786 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0013786 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0013786 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0013786 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0013786 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0013786 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0013786 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0013786 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0013786 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0013786 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0013786 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0013786 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0013786 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0013786 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0013786 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0013786 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0013786 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0013786 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0013786 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0013786 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0013786 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0013786 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0013786 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0013786 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0013786 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0013786 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0013786 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0013786 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0013786 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0013786 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0013786 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0013786 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0013786 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0013786 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0013786 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0013786 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0013786 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0013786 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0013786 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0013786 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0013786 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0013786 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0013786 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0013786 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0013786 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0013786 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0013786 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0013786 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0013786 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0013786 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0013786 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0013786 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0013786 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0013786 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0013786 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0013786 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0013786 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0013786 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0013786 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0013786 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0013786 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0013786 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0013786 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0013786 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0013786 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0013786 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0013786 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0013786 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0013786 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0013786 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0013786 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0013786 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0013786 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0013786 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0013786 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0013786 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0013786 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0013786 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0013786 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0013786 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0013786 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0013786 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0013786 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0013786 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0013786 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0013786 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0013786 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0013786 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0013786 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0013786 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0013786 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0013786 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0013786 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0013786 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0013786 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0013786 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0013786 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0013786 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0013786 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0013786 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0013786 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0013786 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0013786 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0013786 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0013786 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0013786 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0013786 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0013786 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0013786 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0013786 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0013786 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0013786 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0013786 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0013786 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0013786 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0013786 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0013786 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0013786 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0013786 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0013786 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0013786 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0013786 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0013786 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0013786 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0013786 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0013786 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0013786 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0013786 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0013786 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0013786 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0013786 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0013786 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0013786 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0013786 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0013786 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0013786 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0013786 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0013786 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0013786 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0013786 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0013786 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0013786 5.10165e-08 0)
L_DFF_IP1_01_|1 IP1_0_OUT_ _DFF_IP1_01_|A1  2.067833848e-12
L_DFF_IP1_01_|2 _DFF_IP1_01_|A1 _DFF_IP1_01_|A2  4.135667696e-12
L_DFF_IP1_01_|3 _DFF_IP1_01_|A3 _DFF_IP1_01_|A4  8.271335392e-12
L_DFF_IP1_01_|T D01_ _DFF_IP1_01_|T1  2.067833848e-12
L_DFF_IP1_01_|4 _DFF_IP1_01_|T1 _DFF_IP1_01_|T2  4.135667696e-12
L_DFF_IP1_01_|5 _DFF_IP1_01_|A4 _DFF_IP1_01_|Q1  4.135667696e-12
L_DFF_IP1_01_|6 _DFF_IP1_01_|Q1 IP1_1_OUT_  2.067833848e-12
ID02_|T 0 D02_  PWL(0 0 1.35e-11 0 1.5e-11 0.0013786 1.65e-11 0 2.135e-10 0 2.15e-10 0.0013786 2.165e-10 0 4.135e-10 0 4.15e-10 0.0013786 4.165e-10 0 6.135e-10 0 6.15e-10 0.0013786 6.165e-10 0 8.135e-10 0 8.15e-10 0.0013786 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0013786 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0013786 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0013786 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0013786 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0013786 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0013786 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0013786 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0013786 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0013786 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0013786 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0013786 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0013786 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0013786 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0013786 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0013786 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0013786 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0013786 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0013786 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0013786 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0013786 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0013786 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0013786 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0013786 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0013786 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0013786 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0013786 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0013786 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0013786 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0013786 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0013786 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0013786 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0013786 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0013786 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0013786 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0013786 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0013786 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0013786 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0013786 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0013786 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0013786 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0013786 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0013786 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0013786 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0013786 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0013786 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0013786 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0013786 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0013786 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0013786 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0013786 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0013786 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0013786 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0013786 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0013786 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0013786 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0013786 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0013786 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0013786 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0013786 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0013786 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0013786 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0013786 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0013786 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0013786 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0013786 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0013786 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0013786 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0013786 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0013786 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0013786 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0013786 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0013786 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0013786 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0013786 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0013786 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0013786 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0013786 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0013786 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0013786 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0013786 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0013786 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0013786 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0013786 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0013786 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0013786 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0013786 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0013786 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0013786 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0013786 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0013786 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0013786 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0013786 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0013786 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0013786 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0013786 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0013786 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0013786 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0013786 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0013786 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0013786 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0013786 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0013786 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0013786 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0013786 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0013786 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0013786 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0013786 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0013786 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0013786 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0013786 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0013786 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0013786 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0013786 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0013786 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0013786 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0013786 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0013786 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0013786 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0013786 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0013786 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0013786 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0013786 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0013786 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0013786 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0013786 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0013786 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0013786 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0013786 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0013786 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0013786 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0013786 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0013786 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0013786 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0013786 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0013786 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0013786 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0013786 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0013786 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0013786 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0013786 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0013786 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0013786 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0013786 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0013786 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0013786 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0013786 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0013786 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0013786 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0013786 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0013786 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0013786 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0013786 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0013786 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0013786 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0013786 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0013786 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0013786 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0013786 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0013786 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0013786 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0013786 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0013786 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0013786 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0013786 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0013786 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0013786 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0013786 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0013786 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0013786 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0013786 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0013786 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0013786 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0013786 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0013786 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0013786 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0013786 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0013786 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0013786 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0013786 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0013786 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0013786 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0013786 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0013786 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0013786 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0013786 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0013786 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0013786 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0013786 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0013786 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0013786 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0013786 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0013786 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0013786 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0013786 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0013786 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0013786 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0013786 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0013786 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0013786 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0013786 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0013786 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0013786 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0013786 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0013786 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0013786 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0013786 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0013786 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0013786 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0013786 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0013786 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0013786 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0013786 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0013786 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0013786 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0013786 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0013786 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0013786 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0013786 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0013786 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0013786 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0013786 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0013786 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0013786 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0013786 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0013786 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0013786 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0013786 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0013786 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0013786 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0013786 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0013786 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0013786 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0013786 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0013786 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0013786 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0013786 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0013786 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0013786 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0013786 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0013786 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0013786 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0013786 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0013786 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0013786 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0013786 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0013786 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0013786 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0013786 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0013786 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0013786 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0013786 5.10165e-08 0)
L_DFF_IP2_01_|1 IP2_0_OUT_ _DFF_IP2_01_|A1  2.067833848e-12
L_DFF_IP2_01_|2 _DFF_IP2_01_|A1 _DFF_IP2_01_|A2  4.135667696e-12
L_DFF_IP2_01_|3 _DFF_IP2_01_|A3 _DFF_IP2_01_|A4  8.271335392e-12
L_DFF_IP2_01_|T D02_ _DFF_IP2_01_|T1  2.067833848e-12
L_DFF_IP2_01_|4 _DFF_IP2_01_|T1 _DFF_IP2_01_|T2  4.135667696e-12
L_DFF_IP2_01_|5 _DFF_IP2_01_|A4 _DFF_IP2_01_|Q1  4.135667696e-12
L_DFF_IP2_01_|6 _DFF_IP2_01_|Q1 IP2_1_OUT_  2.067833848e-12
ID03_|T 0 D03_  PWL(0 0 1.35e-11 0 1.5e-11 0.0013786 1.65e-11 0 2.135e-10 0 2.15e-10 0.0013786 2.165e-10 0 4.135e-10 0 4.15e-10 0.0013786 4.165e-10 0 6.135e-10 0 6.15e-10 0.0013786 6.165e-10 0 8.135e-10 0 8.15e-10 0.0013786 8.165e-10 0 1.0135e-09 0 1.015e-09 0.0013786 1.0165e-09 0 1.2135e-09 0 1.215e-09 0.0013786 1.2165e-09 0 1.4135e-09 0 1.415e-09 0.0013786 1.4165e-09 0 1.6135e-09 0 1.615e-09 0.0013786 1.6165e-09 0 1.8135e-09 0 1.815e-09 0.0013786 1.8165e-09 0 2.0135e-09 0 2.015e-09 0.0013786 2.0165e-09 0 2.2135e-09 0 2.215e-09 0.0013786 2.2165e-09 0 2.4135e-09 0 2.415e-09 0.0013786 2.4165e-09 0 2.6135e-09 0 2.615e-09 0.0013786 2.6165e-09 0 2.8135e-09 0 2.815e-09 0.0013786 2.8165e-09 0 3.0135e-09 0 3.015e-09 0.0013786 3.0165e-09 0 3.2135e-09 0 3.215e-09 0.0013786 3.2165e-09 0 3.4135e-09 0 3.415e-09 0.0013786 3.4165e-09 0 3.6135e-09 0 3.615e-09 0.0013786 3.6165e-09 0 3.8135e-09 0 3.815e-09 0.0013786 3.8165e-09 0 4.0135e-09 0 4.015e-09 0.0013786 4.0165e-09 0 4.2135e-09 0 4.215e-09 0.0013786 4.2165e-09 0 4.4135e-09 0 4.415e-09 0.0013786 4.4165e-09 0 4.6135e-09 0 4.615e-09 0.0013786 4.6165e-09 0 4.8135e-09 0 4.815e-09 0.0013786 4.8165e-09 0 5.0135e-09 0 5.015e-09 0.0013786 5.0165e-09 0 5.2135e-09 0 5.215e-09 0.0013786 5.2165e-09 0 5.4135e-09 0 5.415e-09 0.0013786 5.4165e-09 0 5.6135e-09 0 5.615e-09 0.0013786 5.6165e-09 0 5.8135e-09 0 5.815e-09 0.0013786 5.8165e-09 0 6.0135e-09 0 6.015e-09 0.0013786 6.0165e-09 0 6.2135e-09 0 6.215e-09 0.0013786 6.2165e-09 0 6.4135e-09 0 6.415e-09 0.0013786 6.4165e-09 0 6.6135e-09 0 6.615e-09 0.0013786 6.6165e-09 0 6.8135e-09 0 6.815e-09 0.0013786 6.8165e-09 0 7.0135e-09 0 7.015e-09 0.0013786 7.0165e-09 0 7.2135e-09 0 7.215e-09 0.0013786 7.2165e-09 0 7.4135e-09 0 7.415e-09 0.0013786 7.4165e-09 0 7.6135e-09 0 7.615e-09 0.0013786 7.6165e-09 0 7.8135e-09 0 7.815e-09 0.0013786 7.8165e-09 0 8.0135e-09 0 8.015e-09 0.0013786 8.0165e-09 0 8.2135e-09 0 8.215e-09 0.0013786 8.2165e-09 0 8.4135e-09 0 8.415e-09 0.0013786 8.4165e-09 0 8.6135e-09 0 8.615e-09 0.0013786 8.6165e-09 0 8.8135e-09 0 8.815e-09 0.0013786 8.8165e-09 0 9.0135e-09 0 9.015e-09 0.0013786 9.0165e-09 0 9.2135e-09 0 9.215e-09 0.0013786 9.2165e-09 0 9.4135e-09 0 9.415e-09 0.0013786 9.4165e-09 0 9.6135e-09 0 9.615e-09 0.0013786 9.6165e-09 0 9.8135e-09 0 9.815e-09 0.0013786 9.8165e-09 0 1.00135e-08 0 1.0015e-08 0.0013786 1.00165e-08 0 1.02135e-08 0 1.0215e-08 0.0013786 1.02165e-08 0 1.04135e-08 0 1.0415e-08 0.0013786 1.04165e-08 0 1.06135e-08 0 1.0615e-08 0.0013786 1.06165e-08 0 1.08135e-08 0 1.0815e-08 0.0013786 1.08165e-08 0 1.10135e-08 0 1.1015e-08 0.0013786 1.10165e-08 0 1.12135e-08 0 1.1215e-08 0.0013786 1.12165e-08 0 1.14135e-08 0 1.1415e-08 0.0013786 1.14165e-08 0 1.16135e-08 0 1.1615e-08 0.0013786 1.16165e-08 0 1.18135e-08 0 1.1815e-08 0.0013786 1.18165e-08 0 1.20135e-08 0 1.2015e-08 0.0013786 1.20165e-08 0 1.22135e-08 0 1.2215e-08 0.0013786 1.22165e-08 0 1.24135e-08 0 1.2415e-08 0.0013786 1.24165e-08 0 1.26135e-08 0 1.2615e-08 0.0013786 1.26165e-08 0 1.28135e-08 0 1.2815e-08 0.0013786 1.28165e-08 0 1.30135e-08 0 1.3015e-08 0.0013786 1.30165e-08 0 1.32135e-08 0 1.3215e-08 0.0013786 1.32165e-08 0 1.34135e-08 0 1.3415e-08 0.0013786 1.34165e-08 0 1.36135e-08 0 1.3615e-08 0.0013786 1.36165e-08 0 1.38135e-08 0 1.3815e-08 0.0013786 1.38165e-08 0 1.40135e-08 0 1.4015e-08 0.0013786 1.40165e-08 0 1.42135e-08 0 1.4215e-08 0.0013786 1.42165e-08 0 1.44135e-08 0 1.4415e-08 0.0013786 1.44165e-08 0 1.46135e-08 0 1.4615e-08 0.0013786 1.46165e-08 0 1.48135e-08 0 1.4815e-08 0.0013786 1.48165e-08 0 1.50135e-08 0 1.5015e-08 0.0013786 1.50165e-08 0 1.52135e-08 0 1.5215e-08 0.0013786 1.52165e-08 0 1.54135e-08 0 1.5415e-08 0.0013786 1.54165e-08 0 1.56135e-08 0 1.5615e-08 0.0013786 1.56165e-08 0 1.58135e-08 0 1.5815e-08 0.0013786 1.58165e-08 0 1.60135e-08 0 1.6015e-08 0.0013786 1.60165e-08 0 1.62135e-08 0 1.6215e-08 0.0013786 1.62165e-08 0 1.64135e-08 0 1.6415e-08 0.0013786 1.64165e-08 0 1.66135e-08 0 1.6615e-08 0.0013786 1.66165e-08 0 1.68135e-08 0 1.6815e-08 0.0013786 1.68165e-08 0 1.70135e-08 0 1.7015e-08 0.0013786 1.70165e-08 0 1.72135e-08 0 1.7215e-08 0.0013786 1.72165e-08 0 1.74135e-08 0 1.7415e-08 0.0013786 1.74165e-08 0 1.76135e-08 0 1.7615e-08 0.0013786 1.76165e-08 0 1.78135e-08 0 1.7815e-08 0.0013786 1.78165e-08 0 1.80135e-08 0 1.8015e-08 0.0013786 1.80165e-08 0 1.82135e-08 0 1.8215e-08 0.0013786 1.82165e-08 0 1.84135e-08 0 1.8415e-08 0.0013786 1.84165e-08 0 1.86135e-08 0 1.8615e-08 0.0013786 1.86165e-08 0 1.88135e-08 0 1.8815e-08 0.0013786 1.88165e-08 0 1.90135e-08 0 1.9015e-08 0.0013786 1.90165e-08 0 1.92135e-08 0 1.9215e-08 0.0013786 1.92165e-08 0 1.94135e-08 0 1.9415e-08 0.0013786 1.94165e-08 0 1.96135e-08 0 1.9615e-08 0.0013786 1.96165e-08 0 1.98135e-08 0 1.9815e-08 0.0013786 1.98165e-08 0 2.00135e-08 0 2.0015e-08 0.0013786 2.00165e-08 0 2.02135e-08 0 2.0215e-08 0.0013786 2.02165e-08 0 2.04135e-08 0 2.0415e-08 0.0013786 2.04165e-08 0 2.06135e-08 0 2.0615e-08 0.0013786 2.06165e-08 0 2.08135e-08 0 2.0815e-08 0.0013786 2.08165e-08 0 2.10135e-08 0 2.1015e-08 0.0013786 2.10165e-08 0 2.12135e-08 0 2.1215e-08 0.0013786 2.12165e-08 0 2.14135e-08 0 2.1415e-08 0.0013786 2.14165e-08 0 2.16135e-08 0 2.1615e-08 0.0013786 2.16165e-08 0 2.18135e-08 0 2.1815e-08 0.0013786 2.18165e-08 0 2.20135e-08 0 2.2015e-08 0.0013786 2.20165e-08 0 2.22135e-08 0 2.2215e-08 0.0013786 2.22165e-08 0 2.24135e-08 0 2.2415e-08 0.0013786 2.24165e-08 0 2.26135e-08 0 2.2615e-08 0.0013786 2.26165e-08 0 2.28135e-08 0 2.2815e-08 0.0013786 2.28165e-08 0 2.30135e-08 0 2.3015e-08 0.0013786 2.30165e-08 0 2.32135e-08 0 2.3215e-08 0.0013786 2.32165e-08 0 2.34135e-08 0 2.3415e-08 0.0013786 2.34165e-08 0 2.36135e-08 0 2.3615e-08 0.0013786 2.36165e-08 0 2.38135e-08 0 2.3815e-08 0.0013786 2.38165e-08 0 2.40135e-08 0 2.4015e-08 0.0013786 2.40165e-08 0 2.42135e-08 0 2.4215e-08 0.0013786 2.42165e-08 0 2.44135e-08 0 2.4415e-08 0.0013786 2.44165e-08 0 2.46135e-08 0 2.4615e-08 0.0013786 2.46165e-08 0 2.48135e-08 0 2.4815e-08 0.0013786 2.48165e-08 0 2.50135e-08 0 2.5015e-08 0.0013786 2.50165e-08 0 2.52135e-08 0 2.5215e-08 0.0013786 2.52165e-08 0 2.54135e-08 0 2.5415e-08 0.0013786 2.54165e-08 0 2.56135e-08 0 2.5615e-08 0.0013786 2.56165e-08 0 2.58135e-08 0 2.5815e-08 0.0013786 2.58165e-08 0 2.60135e-08 0 2.6015e-08 0.0013786 2.60165e-08 0 2.62135e-08 0 2.6215e-08 0.0013786 2.62165e-08 0 2.64135e-08 0 2.6415e-08 0.0013786 2.64165e-08 0 2.66135e-08 0 2.6615e-08 0.0013786 2.66165e-08 0 2.68135e-08 0 2.6815e-08 0.0013786 2.68165e-08 0 2.70135e-08 0 2.7015e-08 0.0013786 2.70165e-08 0 2.72135e-08 0 2.7215e-08 0.0013786 2.72165e-08 0 2.74135e-08 0 2.7415e-08 0.0013786 2.74165e-08 0 2.76135e-08 0 2.7615e-08 0.0013786 2.76165e-08 0 2.78135e-08 0 2.7815e-08 0.0013786 2.78165e-08 0 2.80135e-08 0 2.8015e-08 0.0013786 2.80165e-08 0 2.82135e-08 0 2.8215e-08 0.0013786 2.82165e-08 0 2.84135e-08 0 2.8415e-08 0.0013786 2.84165e-08 0 2.86135e-08 0 2.8615e-08 0.0013786 2.86165e-08 0 2.88135e-08 0 2.8815e-08 0.0013786 2.88165e-08 0 2.90135e-08 0 2.9015e-08 0.0013786 2.90165e-08 0 2.92135e-08 0 2.9215e-08 0.0013786 2.92165e-08 0 2.94135e-08 0 2.9415e-08 0.0013786 2.94165e-08 0 2.96135e-08 0 2.9615e-08 0.0013786 2.96165e-08 0 2.98135e-08 0 2.9815e-08 0.0013786 2.98165e-08 0 3.00135e-08 0 3.0015e-08 0.0013786 3.00165e-08 0 3.02135e-08 0 3.0215e-08 0.0013786 3.02165e-08 0 3.04135e-08 0 3.0415e-08 0.0013786 3.04165e-08 0 3.06135e-08 0 3.0615e-08 0.0013786 3.06165e-08 0 3.08135e-08 0 3.0815e-08 0.0013786 3.08165e-08 0 3.10135e-08 0 3.1015e-08 0.0013786 3.10165e-08 0 3.12135e-08 0 3.1215e-08 0.0013786 3.12165e-08 0 3.14135e-08 0 3.1415e-08 0.0013786 3.14165e-08 0 3.16135e-08 0 3.1615e-08 0.0013786 3.16165e-08 0 3.18135e-08 0 3.1815e-08 0.0013786 3.18165e-08 0 3.20135e-08 0 3.2015e-08 0.0013786 3.20165e-08 0 3.22135e-08 0 3.2215e-08 0.0013786 3.22165e-08 0 3.24135e-08 0 3.2415e-08 0.0013786 3.24165e-08 0 3.26135e-08 0 3.2615e-08 0.0013786 3.26165e-08 0 3.28135e-08 0 3.2815e-08 0.0013786 3.28165e-08 0 3.30135e-08 0 3.3015e-08 0.0013786 3.30165e-08 0 3.32135e-08 0 3.3215e-08 0.0013786 3.32165e-08 0 3.34135e-08 0 3.3415e-08 0.0013786 3.34165e-08 0 3.36135e-08 0 3.3615e-08 0.0013786 3.36165e-08 0 3.38135e-08 0 3.3815e-08 0.0013786 3.38165e-08 0 3.40135e-08 0 3.4015e-08 0.0013786 3.40165e-08 0 3.42135e-08 0 3.4215e-08 0.0013786 3.42165e-08 0 3.44135e-08 0 3.4415e-08 0.0013786 3.44165e-08 0 3.46135e-08 0 3.4615e-08 0.0013786 3.46165e-08 0 3.48135e-08 0 3.4815e-08 0.0013786 3.48165e-08 0 3.50135e-08 0 3.5015e-08 0.0013786 3.50165e-08 0 3.52135e-08 0 3.5215e-08 0.0013786 3.52165e-08 0 3.54135e-08 0 3.5415e-08 0.0013786 3.54165e-08 0 3.56135e-08 0 3.5615e-08 0.0013786 3.56165e-08 0 3.58135e-08 0 3.5815e-08 0.0013786 3.58165e-08 0 3.60135e-08 0 3.6015e-08 0.0013786 3.60165e-08 0 3.62135e-08 0 3.6215e-08 0.0013786 3.62165e-08 0 3.64135e-08 0 3.6415e-08 0.0013786 3.64165e-08 0 3.66135e-08 0 3.6615e-08 0.0013786 3.66165e-08 0 3.68135e-08 0 3.6815e-08 0.0013786 3.68165e-08 0 3.70135e-08 0 3.7015e-08 0.0013786 3.70165e-08 0 3.72135e-08 0 3.7215e-08 0.0013786 3.72165e-08 0 3.74135e-08 0 3.7415e-08 0.0013786 3.74165e-08 0 3.76135e-08 0 3.7615e-08 0.0013786 3.76165e-08 0 3.78135e-08 0 3.7815e-08 0.0013786 3.78165e-08 0 3.80135e-08 0 3.8015e-08 0.0013786 3.80165e-08 0 3.82135e-08 0 3.8215e-08 0.0013786 3.82165e-08 0 3.84135e-08 0 3.8415e-08 0.0013786 3.84165e-08 0 3.86135e-08 0 3.8615e-08 0.0013786 3.86165e-08 0 3.88135e-08 0 3.8815e-08 0.0013786 3.88165e-08 0 3.90135e-08 0 3.9015e-08 0.0013786 3.90165e-08 0 3.92135e-08 0 3.9215e-08 0.0013786 3.92165e-08 0 3.94135e-08 0 3.9415e-08 0.0013786 3.94165e-08 0 3.96135e-08 0 3.9615e-08 0.0013786 3.96165e-08 0 3.98135e-08 0 3.9815e-08 0.0013786 3.98165e-08 0 4.00135e-08 0 4.0015e-08 0.0013786 4.00165e-08 0 4.02135e-08 0 4.0215e-08 0.0013786 4.02165e-08 0 4.04135e-08 0 4.0415e-08 0.0013786 4.04165e-08 0 4.06135e-08 0 4.0615e-08 0.0013786 4.06165e-08 0 4.08135e-08 0 4.0815e-08 0.0013786 4.08165e-08 0 4.10135e-08 0 4.1015e-08 0.0013786 4.10165e-08 0 4.12135e-08 0 4.1215e-08 0.0013786 4.12165e-08 0 4.14135e-08 0 4.1415e-08 0.0013786 4.14165e-08 0 4.16135e-08 0 4.1615e-08 0.0013786 4.16165e-08 0 4.18135e-08 0 4.1815e-08 0.0013786 4.18165e-08 0 4.20135e-08 0 4.2015e-08 0.0013786 4.20165e-08 0 4.22135e-08 0 4.2215e-08 0.0013786 4.22165e-08 0 4.24135e-08 0 4.2415e-08 0.0013786 4.24165e-08 0 4.26135e-08 0 4.2615e-08 0.0013786 4.26165e-08 0 4.28135e-08 0 4.2815e-08 0.0013786 4.28165e-08 0 4.30135e-08 0 4.3015e-08 0.0013786 4.30165e-08 0 4.32135e-08 0 4.3215e-08 0.0013786 4.32165e-08 0 4.34135e-08 0 4.3415e-08 0.0013786 4.34165e-08 0 4.36135e-08 0 4.3615e-08 0.0013786 4.36165e-08 0 4.38135e-08 0 4.3815e-08 0.0013786 4.38165e-08 0 4.40135e-08 0 4.4015e-08 0.0013786 4.40165e-08 0 4.42135e-08 0 4.4215e-08 0.0013786 4.42165e-08 0 4.44135e-08 0 4.4415e-08 0.0013786 4.44165e-08 0 4.46135e-08 0 4.4615e-08 0.0013786 4.46165e-08 0 4.48135e-08 0 4.4815e-08 0.0013786 4.48165e-08 0 4.50135e-08 0 4.5015e-08 0.0013786 4.50165e-08 0 4.52135e-08 0 4.5215e-08 0.0013786 4.52165e-08 0 4.54135e-08 0 4.5415e-08 0.0013786 4.54165e-08 0 4.56135e-08 0 4.5615e-08 0.0013786 4.56165e-08 0 4.58135e-08 0 4.5815e-08 0.0013786 4.58165e-08 0 4.60135e-08 0 4.6015e-08 0.0013786 4.60165e-08 0 4.62135e-08 0 4.6215e-08 0.0013786 4.62165e-08 0 4.64135e-08 0 4.6415e-08 0.0013786 4.64165e-08 0 4.66135e-08 0 4.6615e-08 0.0013786 4.66165e-08 0 4.68135e-08 0 4.6815e-08 0.0013786 4.68165e-08 0 4.70135e-08 0 4.7015e-08 0.0013786 4.70165e-08 0 4.72135e-08 0 4.7215e-08 0.0013786 4.72165e-08 0 4.74135e-08 0 4.7415e-08 0.0013786 4.74165e-08 0 4.76135e-08 0 4.7615e-08 0.0013786 4.76165e-08 0 4.78135e-08 0 4.7815e-08 0.0013786 4.78165e-08 0 4.80135e-08 0 4.8015e-08 0.0013786 4.80165e-08 0 4.82135e-08 0 4.8215e-08 0.0013786 4.82165e-08 0 4.84135e-08 0 4.8415e-08 0.0013786 4.84165e-08 0 4.86135e-08 0 4.8615e-08 0.0013786 4.86165e-08 0 4.88135e-08 0 4.8815e-08 0.0013786 4.88165e-08 0 4.90135e-08 0 4.9015e-08 0.0013786 4.90165e-08 0 4.92135e-08 0 4.9215e-08 0.0013786 4.92165e-08 0 4.94135e-08 0 4.9415e-08 0.0013786 4.94165e-08 0 4.96135e-08 0 4.9615e-08 0.0013786 4.96165e-08 0 4.98135e-08 0 4.9815e-08 0.0013786 4.98165e-08 0 5.00135e-08 0 5.0015e-08 0.0013786 5.00165e-08 0 5.02135e-08 0 5.0215e-08 0.0013786 5.02165e-08 0 5.04135e-08 0 5.0415e-08 0.0013786 5.04165e-08 0 5.06135e-08 0 5.0615e-08 0.0013786 5.06165e-08 0 5.08135e-08 0 5.0815e-08 0.0013786 5.08165e-08 0 5.10135e-08 0 5.1015e-08 0.0013786 5.10165e-08 0)
L_DFF_IP3_01_|1 IP3_0_OUT_ _DFF_IP3_01_|A1  2.067833848e-12
L_DFF_IP3_01_|2 _DFF_IP3_01_|A1 _DFF_IP3_01_|A2  4.135667696e-12
L_DFF_IP3_01_|3 _DFF_IP3_01_|A3 _DFF_IP3_01_|A4  8.271335392e-12
L_DFF_IP3_01_|T D03_ _DFF_IP3_01_|T1  2.067833848e-12
L_DFF_IP3_01_|4 _DFF_IP3_01_|T1 _DFF_IP3_01_|T2  4.135667696e-12
L_DFF_IP3_01_|5 _DFF_IP3_01_|A4 _DFF_IP3_01_|Q1  4.135667696e-12
L_DFF_IP3_01_|6 _DFF_IP3_01_|Q1 IP3_1_OUT_  2.067833848e-12
LI0_|_SPL_A|1 A0_ I0_|_SPL_A|D1  2e-12
LI0_|_SPL_A|2 I0_|_SPL_A|D1 I0_|_SPL_A|D2  4.135667696e-12
LI0_|_SPL_A|3 I0_|_SPL_A|D2 I0_|_SPL_A|JCT  9.84682784761905e-13
LI0_|_SPL_A|4 I0_|_SPL_A|JCT I0_|_SPL_A|QA1  9.84682784761905e-13
LI0_|_SPL_A|5 I0_|_SPL_A|QA1 I0_|A1  2e-12
LI0_|_SPL_A|6 I0_|_SPL_A|JCT I0_|_SPL_A|QB1  9.84682784761905e-13
LI0_|_SPL_A|7 I0_|_SPL_A|QB1 I0_|A2  2e-12
LI0_|_SPL_B|1 B0_ I0_|_SPL_B|D1  2e-12
LI0_|_SPL_B|2 I0_|_SPL_B|D1 I0_|_SPL_B|D2  4.135667696e-12
LI0_|_SPL_B|3 I0_|_SPL_B|D2 I0_|_SPL_B|JCT  9.84682784761905e-13
LI0_|_SPL_B|4 I0_|_SPL_B|JCT I0_|_SPL_B|QA1  9.84682784761905e-13
LI0_|_SPL_B|5 I0_|_SPL_B|QA1 I0_|B1  2e-12
LI0_|_SPL_B|6 I0_|_SPL_B|JCT I0_|_SPL_B|QB1  9.84682784761905e-13
LI0_|_SPL_B|7 I0_|_SPL_B|QB1 I0_|B2  2e-12
LI0_|_DFF_A|1 I0_|A1 I0_|_DFF_A|A1  2.067833848e-12
LI0_|_DFF_A|2 I0_|_DFF_A|A1 I0_|_DFF_A|A2  4.135667696e-12
LI0_|_DFF_A|3 I0_|_DFF_A|A3 I0_|_DFF_A|A4  8.271335392e-12
LI0_|_DFF_A|T T00_ I0_|_DFF_A|T1  2.067833848e-12
LI0_|_DFF_A|4 I0_|_DFF_A|T1 I0_|_DFF_A|T2  4.135667696e-12
LI0_|_DFF_A|5 I0_|_DFF_A|A4 I0_|_DFF_A|Q1  4.135667696e-12
LI0_|_DFF_A|6 I0_|_DFF_A|Q1 I0_|A1_SYNC  2.067833848e-12
LI0_|_DFF_B|1 I0_|B1 I0_|_DFF_B|A1  2.067833848e-12
LI0_|_DFF_B|2 I0_|_DFF_B|A1 I0_|_DFF_B|A2  4.135667696e-12
LI0_|_DFF_B|3 I0_|_DFF_B|A3 I0_|_DFF_B|A4  8.271335392e-12
LI0_|_DFF_B|T T00_ I0_|_DFF_B|T1  2.067833848e-12
LI0_|_DFF_B|4 I0_|_DFF_B|T1 I0_|_DFF_B|T2  4.135667696e-12
LI0_|_DFF_B|5 I0_|_DFF_B|A4 I0_|_DFF_B|Q1  4.135667696e-12
LI0_|_DFF_B|6 I0_|_DFF_B|Q1 I0_|B1_SYNC  2.067833848e-12
LI0_|_XOR|A1 I0_|A2 I0_|_XOR|A1  2.067833848e-12
LI0_|_XOR|A2 I0_|_XOR|A1 I0_|_XOR|A2  4.135667696e-12
LI0_|_XOR|A3 I0_|_XOR|A3 I0_|_XOR|AB  8.271335392e-12
LI0_|_XOR|B1 I0_|B2 I0_|_XOR|B1  2.067833848e-12
LI0_|_XOR|B2 I0_|_XOR|B1 I0_|_XOR|B2  4.135667696e-12
LI0_|_XOR|B3 I0_|_XOR|B3 I0_|_XOR|AB  8.271335392e-12
LI0_|_XOR|T1 T00_ I0_|_XOR|T1  2.067833848e-12
LI0_|_XOR|T2 I0_|_XOR|T1 I0_|_XOR|T2  4.135667696e-12
LI0_|_XOR|Q2 I0_|_XOR|ABTQ I0_|_XOR|Q1  4.135667696e-12
LI0_|_XOR|Q1 I0_|_XOR|Q1 IP0_0_  2.067833848e-12
LI0_|_AND|A1 I0_|A1_SYNC I0_|_AND|A1  2.067833848e-12
LI0_|_AND|A2 I0_|_AND|A1 I0_|_AND|A2  4.135667696e-12
LI0_|_AND|A3 I0_|_AND|A3 I0_|_AND|Q3  1.2e-12
LI0_|_AND|B1 I0_|B1_SYNC I0_|_AND|B1  2.067833848e-12
LI0_|_AND|B2 I0_|_AND|B1 I0_|_AND|B2  4.135667696e-12
LI0_|_AND|B3 I0_|_AND|B3 I0_|_AND|Q3  1.2e-12
LI0_|_AND|Q3 I0_|_AND|Q3 I0_|_AND|Q2  4.135667696e-12
LI0_|_AND|Q2 I0_|_AND|Q2 I0_|_AND|Q1  4.135667696e-12
LI0_|_AND|Q1 I0_|_AND|Q1 IG0_0_  2.067833848e-12
LI1_|_SPL_A|1 A1_ I1_|_SPL_A|D1  2e-12
LI1_|_SPL_A|2 I1_|_SPL_A|D1 I1_|_SPL_A|D2  4.135667696e-12
LI1_|_SPL_A|3 I1_|_SPL_A|D2 I1_|_SPL_A|JCT  9.84682784761905e-13
LI1_|_SPL_A|4 I1_|_SPL_A|JCT I1_|_SPL_A|QA1  9.84682784761905e-13
LI1_|_SPL_A|5 I1_|_SPL_A|QA1 I1_|A1  2e-12
LI1_|_SPL_A|6 I1_|_SPL_A|JCT I1_|_SPL_A|QB1  9.84682784761905e-13
LI1_|_SPL_A|7 I1_|_SPL_A|QB1 I1_|A2  2e-12
LI1_|_SPL_B|1 B1_ I1_|_SPL_B|D1  2e-12
LI1_|_SPL_B|2 I1_|_SPL_B|D1 I1_|_SPL_B|D2  4.135667696e-12
LI1_|_SPL_B|3 I1_|_SPL_B|D2 I1_|_SPL_B|JCT  9.84682784761905e-13
LI1_|_SPL_B|4 I1_|_SPL_B|JCT I1_|_SPL_B|QA1  9.84682784761905e-13
LI1_|_SPL_B|5 I1_|_SPL_B|QA1 I1_|B1  2e-12
LI1_|_SPL_B|6 I1_|_SPL_B|JCT I1_|_SPL_B|QB1  9.84682784761905e-13
LI1_|_SPL_B|7 I1_|_SPL_B|QB1 I1_|B2  2e-12
LI1_|_DFF_A|1 I1_|A1 I1_|_DFF_A|A1  2.067833848e-12
LI1_|_DFF_A|2 I1_|_DFF_A|A1 I1_|_DFF_A|A2  4.135667696e-12
LI1_|_DFF_A|3 I1_|_DFF_A|A3 I1_|_DFF_A|A4  8.271335392e-12
LI1_|_DFF_A|T T01_ I1_|_DFF_A|T1  2.067833848e-12
LI1_|_DFF_A|4 I1_|_DFF_A|T1 I1_|_DFF_A|T2  4.135667696e-12
LI1_|_DFF_A|5 I1_|_DFF_A|A4 I1_|_DFF_A|Q1  4.135667696e-12
LI1_|_DFF_A|6 I1_|_DFF_A|Q1 I1_|A1_SYNC  2.067833848e-12
LI1_|_DFF_B|1 I1_|B1 I1_|_DFF_B|A1  2.067833848e-12
LI1_|_DFF_B|2 I1_|_DFF_B|A1 I1_|_DFF_B|A2  4.135667696e-12
LI1_|_DFF_B|3 I1_|_DFF_B|A3 I1_|_DFF_B|A4  8.271335392e-12
LI1_|_DFF_B|T T01_ I1_|_DFF_B|T1  2.067833848e-12
LI1_|_DFF_B|4 I1_|_DFF_B|T1 I1_|_DFF_B|T2  4.135667696e-12
LI1_|_DFF_B|5 I1_|_DFF_B|A4 I1_|_DFF_B|Q1  4.135667696e-12
LI1_|_DFF_B|6 I1_|_DFF_B|Q1 I1_|B1_SYNC  2.067833848e-12
LI1_|_XOR|A1 I1_|A2 I1_|_XOR|A1  2.067833848e-12
LI1_|_XOR|A2 I1_|_XOR|A1 I1_|_XOR|A2  4.135667696e-12
LI1_|_XOR|A3 I1_|_XOR|A3 I1_|_XOR|AB  8.271335392e-12
LI1_|_XOR|B1 I1_|B2 I1_|_XOR|B1  2.067833848e-12
LI1_|_XOR|B2 I1_|_XOR|B1 I1_|_XOR|B2  4.135667696e-12
LI1_|_XOR|B3 I1_|_XOR|B3 I1_|_XOR|AB  8.271335392e-12
LI1_|_XOR|T1 T01_ I1_|_XOR|T1  2.067833848e-12
LI1_|_XOR|T2 I1_|_XOR|T1 I1_|_XOR|T2  4.135667696e-12
LI1_|_XOR|Q2 I1_|_XOR|ABTQ I1_|_XOR|Q1  4.135667696e-12
LI1_|_XOR|Q1 I1_|_XOR|Q1 IP1_0_  2.067833848e-12
LI1_|_AND|A1 I1_|A1_SYNC I1_|_AND|A1  2.067833848e-12
LI1_|_AND|A2 I1_|_AND|A1 I1_|_AND|A2  4.135667696e-12
LI1_|_AND|A3 I1_|_AND|A3 I1_|_AND|Q3  1.2e-12
LI1_|_AND|B1 I1_|B1_SYNC I1_|_AND|B1  2.067833848e-12
LI1_|_AND|B2 I1_|_AND|B1 I1_|_AND|B2  4.135667696e-12
LI1_|_AND|B3 I1_|_AND|B3 I1_|_AND|Q3  1.2e-12
LI1_|_AND|Q3 I1_|_AND|Q3 I1_|_AND|Q2  4.135667696e-12
LI1_|_AND|Q2 I1_|_AND|Q2 I1_|_AND|Q1  4.135667696e-12
LI1_|_AND|Q1 I1_|_AND|Q1 IG1_0_  2.067833848e-12
LI2_|_SPL_A|1 A2_ I2_|_SPL_A|D1  2e-12
LI2_|_SPL_A|2 I2_|_SPL_A|D1 I2_|_SPL_A|D2  4.135667696e-12
LI2_|_SPL_A|3 I2_|_SPL_A|D2 I2_|_SPL_A|JCT  9.84682784761905e-13
LI2_|_SPL_A|4 I2_|_SPL_A|JCT I2_|_SPL_A|QA1  9.84682784761905e-13
LI2_|_SPL_A|5 I2_|_SPL_A|QA1 I2_|A1  2e-12
LI2_|_SPL_A|6 I2_|_SPL_A|JCT I2_|_SPL_A|QB1  9.84682784761905e-13
LI2_|_SPL_A|7 I2_|_SPL_A|QB1 I2_|A2  2e-12
LI2_|_SPL_B|1 B2_ I2_|_SPL_B|D1  2e-12
LI2_|_SPL_B|2 I2_|_SPL_B|D1 I2_|_SPL_B|D2  4.135667696e-12
LI2_|_SPL_B|3 I2_|_SPL_B|D2 I2_|_SPL_B|JCT  9.84682784761905e-13
LI2_|_SPL_B|4 I2_|_SPL_B|JCT I2_|_SPL_B|QA1  9.84682784761905e-13
LI2_|_SPL_B|5 I2_|_SPL_B|QA1 I2_|B1  2e-12
LI2_|_SPL_B|6 I2_|_SPL_B|JCT I2_|_SPL_B|QB1  9.84682784761905e-13
LI2_|_SPL_B|7 I2_|_SPL_B|QB1 I2_|B2  2e-12
LI2_|_DFF_A|1 I2_|A1 I2_|_DFF_A|A1  2.067833848e-12
LI2_|_DFF_A|2 I2_|_DFF_A|A1 I2_|_DFF_A|A2  4.135667696e-12
LI2_|_DFF_A|3 I2_|_DFF_A|A3 I2_|_DFF_A|A4  8.271335392e-12
LI2_|_DFF_A|T T02_ I2_|_DFF_A|T1  2.067833848e-12
LI2_|_DFF_A|4 I2_|_DFF_A|T1 I2_|_DFF_A|T2  4.135667696e-12
LI2_|_DFF_A|5 I2_|_DFF_A|A4 I2_|_DFF_A|Q1  4.135667696e-12
LI2_|_DFF_A|6 I2_|_DFF_A|Q1 I2_|A1_SYNC  2.067833848e-12
LI2_|_DFF_B|1 I2_|B1 I2_|_DFF_B|A1  2.067833848e-12
LI2_|_DFF_B|2 I2_|_DFF_B|A1 I2_|_DFF_B|A2  4.135667696e-12
LI2_|_DFF_B|3 I2_|_DFF_B|A3 I2_|_DFF_B|A4  8.271335392e-12
LI2_|_DFF_B|T T02_ I2_|_DFF_B|T1  2.067833848e-12
LI2_|_DFF_B|4 I2_|_DFF_B|T1 I2_|_DFF_B|T2  4.135667696e-12
LI2_|_DFF_B|5 I2_|_DFF_B|A4 I2_|_DFF_B|Q1  4.135667696e-12
LI2_|_DFF_B|6 I2_|_DFF_B|Q1 I2_|B1_SYNC  2.067833848e-12
LI2_|_XOR|A1 I2_|A2 I2_|_XOR|A1  2.067833848e-12
LI2_|_XOR|A2 I2_|_XOR|A1 I2_|_XOR|A2  4.135667696e-12
LI2_|_XOR|A3 I2_|_XOR|A3 I2_|_XOR|AB  8.271335392e-12
LI2_|_XOR|B1 I2_|B2 I2_|_XOR|B1  2.067833848e-12
LI2_|_XOR|B2 I2_|_XOR|B1 I2_|_XOR|B2  4.135667696e-12
LI2_|_XOR|B3 I2_|_XOR|B3 I2_|_XOR|AB  8.271335392e-12
LI2_|_XOR|T1 T02_ I2_|_XOR|T1  2.067833848e-12
LI2_|_XOR|T2 I2_|_XOR|T1 I2_|_XOR|T2  4.135667696e-12
LI2_|_XOR|Q2 I2_|_XOR|ABTQ I2_|_XOR|Q1  4.135667696e-12
LI2_|_XOR|Q1 I2_|_XOR|Q1 IP2_0_  2.067833848e-12
LI2_|_AND|A1 I2_|A1_SYNC I2_|_AND|A1  2.067833848e-12
LI2_|_AND|A2 I2_|_AND|A1 I2_|_AND|A2  4.135667696e-12
LI2_|_AND|A3 I2_|_AND|A3 I2_|_AND|Q3  1.2e-12
LI2_|_AND|B1 I2_|B1_SYNC I2_|_AND|B1  2.067833848e-12
LI2_|_AND|B2 I2_|_AND|B1 I2_|_AND|B2  4.135667696e-12
LI2_|_AND|B3 I2_|_AND|B3 I2_|_AND|Q3  1.2e-12
LI2_|_AND|Q3 I2_|_AND|Q3 I2_|_AND|Q2  4.135667696e-12
LI2_|_AND|Q2 I2_|_AND|Q2 I2_|_AND|Q1  4.135667696e-12
LI2_|_AND|Q1 I2_|_AND|Q1 IG2_0_  2.067833848e-12
LI3_|_SPL_A|1 A3_ I3_|_SPL_A|D1  2e-12
LI3_|_SPL_A|2 I3_|_SPL_A|D1 I3_|_SPL_A|D2  4.135667696e-12
LI3_|_SPL_A|3 I3_|_SPL_A|D2 I3_|_SPL_A|JCT  9.84682784761905e-13
LI3_|_SPL_A|4 I3_|_SPL_A|JCT I3_|_SPL_A|QA1  9.84682784761905e-13
LI3_|_SPL_A|5 I3_|_SPL_A|QA1 I3_|A1  2e-12
LI3_|_SPL_A|6 I3_|_SPL_A|JCT I3_|_SPL_A|QB1  9.84682784761905e-13
LI3_|_SPL_A|7 I3_|_SPL_A|QB1 I3_|A2  2e-12
LI3_|_SPL_B|1 B3_ I3_|_SPL_B|D1  2e-12
LI3_|_SPL_B|2 I3_|_SPL_B|D1 I3_|_SPL_B|D2  4.135667696e-12
LI3_|_SPL_B|3 I3_|_SPL_B|D2 I3_|_SPL_B|JCT  9.84682784761905e-13
LI3_|_SPL_B|4 I3_|_SPL_B|JCT I3_|_SPL_B|QA1  9.84682784761905e-13
LI3_|_SPL_B|5 I3_|_SPL_B|QA1 I3_|B1  2e-12
LI3_|_SPL_B|6 I3_|_SPL_B|JCT I3_|_SPL_B|QB1  9.84682784761905e-13
LI3_|_SPL_B|7 I3_|_SPL_B|QB1 I3_|B2  2e-12
LI3_|_DFF_A|1 I3_|A1 I3_|_DFF_A|A1  2.067833848e-12
LI3_|_DFF_A|2 I3_|_DFF_A|A1 I3_|_DFF_A|A2  4.135667696e-12
LI3_|_DFF_A|3 I3_|_DFF_A|A3 I3_|_DFF_A|A4  8.271335392e-12
LI3_|_DFF_A|T T03_ I3_|_DFF_A|T1  2.067833848e-12
LI3_|_DFF_A|4 I3_|_DFF_A|T1 I3_|_DFF_A|T2  4.135667696e-12
LI3_|_DFF_A|5 I3_|_DFF_A|A4 I3_|_DFF_A|Q1  4.135667696e-12
LI3_|_DFF_A|6 I3_|_DFF_A|Q1 I3_|A1_SYNC  2.067833848e-12
LI3_|_DFF_B|1 I3_|B1 I3_|_DFF_B|A1  2.067833848e-12
LI3_|_DFF_B|2 I3_|_DFF_B|A1 I3_|_DFF_B|A2  4.135667696e-12
LI3_|_DFF_B|3 I3_|_DFF_B|A3 I3_|_DFF_B|A4  8.271335392e-12
LI3_|_DFF_B|T T03_ I3_|_DFF_B|T1  2.067833848e-12
LI3_|_DFF_B|4 I3_|_DFF_B|T1 I3_|_DFF_B|T2  4.135667696e-12
LI3_|_DFF_B|5 I3_|_DFF_B|A4 I3_|_DFF_B|Q1  4.135667696e-12
LI3_|_DFF_B|6 I3_|_DFF_B|Q1 I3_|B1_SYNC  2.067833848e-12
LI3_|_XOR|A1 I3_|A2 I3_|_XOR|A1  2.067833848e-12
LI3_|_XOR|A2 I3_|_XOR|A1 I3_|_XOR|A2  4.135667696e-12
LI3_|_XOR|A3 I3_|_XOR|A3 I3_|_XOR|AB  8.271335392e-12
LI3_|_XOR|B1 I3_|B2 I3_|_XOR|B1  2.067833848e-12
LI3_|_XOR|B2 I3_|_XOR|B1 I3_|_XOR|B2  4.135667696e-12
LI3_|_XOR|B3 I3_|_XOR|B3 I3_|_XOR|AB  8.271335392e-12
LI3_|_XOR|T1 T03_ I3_|_XOR|T1  2.067833848e-12
LI3_|_XOR|T2 I3_|_XOR|T1 I3_|_XOR|T2  4.135667696e-12
LI3_|_XOR|Q2 I3_|_XOR|ABTQ I3_|_XOR|Q1  4.135667696e-12
LI3_|_XOR|Q1 I3_|_XOR|Q1 IP3_0_  2.067833848e-12
LI3_|_AND|A1 I3_|A1_SYNC I3_|_AND|A1  2.067833848e-12
LI3_|_AND|A2 I3_|_AND|A1 I3_|_AND|A2  4.135667696e-12
LI3_|_AND|A3 I3_|_AND|A3 I3_|_AND|Q3  1.2e-12
LI3_|_AND|B1 I3_|B1_SYNC I3_|_AND|B1  2.067833848e-12
LI3_|_AND|B2 I3_|_AND|B1 I3_|_AND|B2  4.135667696e-12
LI3_|_AND|B3 I3_|_AND|B3 I3_|_AND|Q3  1.2e-12
LI3_|_AND|Q3 I3_|_AND|Q3 I3_|_AND|Q2  4.135667696e-12
LI3_|_AND|Q2 I3_|_AND|Q2 I3_|_AND|Q1  4.135667696e-12
LI3_|_AND|Q1 I3_|_AND|Q1 IG3_0_  2.067833848e-12
LSPL_IG0_0_|I_D1|B SPL_IG0_0_|D1 SPL_IG0_0_|I_D1|MID  2e-12
ISPL_IG0_0_|I_D1|B 0 SPL_IG0_0_|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IG0_0_|I_D2|B SPL_IG0_0_|D2 SPL_IG0_0_|I_D2|MID  2e-12
ISPL_IG0_0_|I_D2|B 0 SPL_IG0_0_|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IG0_0_|I_Q1|B SPL_IG0_0_|QA1 SPL_IG0_0_|I_Q1|MID  2e-12
ISPL_IG0_0_|I_Q1|B 0 SPL_IG0_0_|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IG0_0_|I_Q2|B SPL_IG0_0_|QB1 SPL_IG0_0_|I_Q2|MID  2e-12
ISPL_IG0_0_|I_Q2|B 0 SPL_IG0_0_|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IG0_0_|1|1 SPL_IG0_0_|D1 SPL_IG0_0_|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0_|1|P SPL_IG0_0_|1|MID_SERIES 0  2e-13
RSPL_IG0_0_|1|B SPL_IG0_0_|D1 SPL_IG0_0_|1|MID_SHUNT  2.7439617672
LSPL_IG0_0_|1|RB SPL_IG0_0_|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0_|2|1 SPL_IG0_0_|D2 SPL_IG0_0_|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0_|2|P SPL_IG0_0_|2|MID_SERIES 0  2e-13
RSPL_IG0_0_|2|B SPL_IG0_0_|D2 SPL_IG0_0_|2|MID_SHUNT  2.7439617672
LSPL_IG0_0_|2|RB SPL_IG0_0_|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0_|A|1 SPL_IG0_0_|QA1 SPL_IG0_0_|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0_|A|P SPL_IG0_0_|A|MID_SERIES 0  2e-13
RSPL_IG0_0_|A|B SPL_IG0_0_|QA1 SPL_IG0_0_|A|MID_SHUNT  2.7439617672
LSPL_IG0_0_|A|RB SPL_IG0_0_|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0_|B|1 SPL_IG0_0_|QB1 SPL_IG0_0_|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0_|B|P SPL_IG0_0_|B|MID_SERIES 0  2e-13
RSPL_IG0_0_|B|B SPL_IG0_0_|QB1 SPL_IG0_0_|B|MID_SHUNT  2.7439617672
LSPL_IG0_0_|B|RB SPL_IG0_0_|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP1_0_|I_D1|B SPL_IP1_0_|D1 SPL_IP1_0_|I_D1|MID  2e-12
ISPL_IP1_0_|I_D1|B 0 SPL_IP1_0_|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP1_0_|I_D2|B SPL_IP1_0_|D2 SPL_IP1_0_|I_D2|MID  2e-12
ISPL_IP1_0_|I_D2|B 0 SPL_IP1_0_|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IP1_0_|I_Q1|B SPL_IP1_0_|QA1 SPL_IP1_0_|I_Q1|MID  2e-12
ISPL_IP1_0_|I_Q1|B 0 SPL_IP1_0_|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP1_0_|I_Q2|B SPL_IP1_0_|QB1 SPL_IP1_0_|I_Q2|MID  2e-12
ISPL_IP1_0_|I_Q2|B 0 SPL_IP1_0_|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IP1_0_|1|1 SPL_IP1_0_|D1 SPL_IP1_0_|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0_|1|P SPL_IP1_0_|1|MID_SERIES 0  2e-13
RSPL_IP1_0_|1|B SPL_IP1_0_|D1 SPL_IP1_0_|1|MID_SHUNT  2.7439617672
LSPL_IP1_0_|1|RB SPL_IP1_0_|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0_|2|1 SPL_IP1_0_|D2 SPL_IP1_0_|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0_|2|P SPL_IP1_0_|2|MID_SERIES 0  2e-13
RSPL_IP1_0_|2|B SPL_IP1_0_|D2 SPL_IP1_0_|2|MID_SHUNT  2.7439617672
LSPL_IP1_0_|2|RB SPL_IP1_0_|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0_|A|1 SPL_IP1_0_|QA1 SPL_IP1_0_|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0_|A|P SPL_IP1_0_|A|MID_SERIES 0  2e-13
RSPL_IP1_0_|A|B SPL_IP1_0_|QA1 SPL_IP1_0_|A|MID_SHUNT  2.7439617672
LSPL_IP1_0_|A|RB SPL_IP1_0_|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0_|B|1 SPL_IP1_0_|QB1 SPL_IP1_0_|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0_|B|P SPL_IP1_0_|B|MID_SERIES 0  2e-13
RSPL_IP1_0_|B|B SPL_IP1_0_|QB1 SPL_IP1_0_|B|MID_SHUNT  2.7439617672
LSPL_IP1_0_|B|RB SPL_IP1_0_|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0_|SPL1|1 IP2_0_ SPL_IP2_0_|SPL1|D1  2e-12
LSPL_IP2_0_|SPL1|2 SPL_IP2_0_|SPL1|D1 SPL_IP2_0_|SPL1|D2  4.135667696e-12
LSPL_IP2_0_|SPL1|3 SPL_IP2_0_|SPL1|D2 SPL_IP2_0_|SPL1|JCT  9.84682784761905e-13
LSPL_IP2_0_|SPL1|4 SPL_IP2_0_|SPL1|JCT SPL_IP2_0_|SPL1|QA1  9.84682784761905e-13
LSPL_IP2_0_|SPL1|5 SPL_IP2_0_|SPL1|QA1 IP2_0_TO2_  2e-12
LSPL_IP2_0_|SPL1|6 SPL_IP2_0_|SPL1|JCT SPL_IP2_0_|SPL1|QB1  9.84682784761905e-13
LSPL_IP2_0_|SPL1|7 SPL_IP2_0_|SPL1|QB1 SPL_IP2_0_|QTMP  2e-12
LSPL_IP2_0_|SPL2|1 SPL_IP2_0_|QTMP SPL_IP2_0_|SPL2|D1  2e-12
LSPL_IP2_0_|SPL2|2 SPL_IP2_0_|SPL2|D1 SPL_IP2_0_|SPL2|D2  4.135667696e-12
LSPL_IP2_0_|SPL2|3 SPL_IP2_0_|SPL2|D2 SPL_IP2_0_|SPL2|JCT  9.84682784761905e-13
LSPL_IP2_0_|SPL2|4 SPL_IP2_0_|SPL2|JCT SPL_IP2_0_|SPL2|QA1  9.84682784761905e-13
LSPL_IP2_0_|SPL2|5 SPL_IP2_0_|SPL2|QA1 IP2_0_TO3_  2e-12
LSPL_IP2_0_|SPL2|6 SPL_IP2_0_|SPL2|JCT SPL_IP2_0_|SPL2|QB1  9.84682784761905e-13
LSPL_IP2_0_|SPL2|7 SPL_IP2_0_|SPL2|QB1 IP2_0_OUT_  2e-12
LSPL_IG2_0_|I_D1|B SPL_IG2_0_|D1 SPL_IG2_0_|I_D1|MID  2e-12
ISPL_IG2_0_|I_D1|B 0 SPL_IG2_0_|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IG2_0_|I_D2|B SPL_IG2_0_|D2 SPL_IG2_0_|I_D2|MID  2e-12
ISPL_IG2_0_|I_D2|B 0 SPL_IG2_0_|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IG2_0_|I_Q1|B SPL_IG2_0_|QA1 SPL_IG2_0_|I_Q1|MID  2e-12
ISPL_IG2_0_|I_Q1|B 0 SPL_IG2_0_|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IG2_0_|I_Q2|B SPL_IG2_0_|QB1 SPL_IG2_0_|I_Q2|MID  2e-12
ISPL_IG2_0_|I_Q2|B 0 SPL_IG2_0_|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IG2_0_|1|1 SPL_IG2_0_|D1 SPL_IG2_0_|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0_|1|P SPL_IG2_0_|1|MID_SERIES 0  2e-13
RSPL_IG2_0_|1|B SPL_IG2_0_|D1 SPL_IG2_0_|1|MID_SHUNT  2.7439617672
LSPL_IG2_0_|1|RB SPL_IG2_0_|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0_|2|1 SPL_IG2_0_|D2 SPL_IG2_0_|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0_|2|P SPL_IG2_0_|2|MID_SERIES 0  2e-13
RSPL_IG2_0_|2|B SPL_IG2_0_|D2 SPL_IG2_0_|2|MID_SHUNT  2.7439617672
LSPL_IG2_0_|2|RB SPL_IG2_0_|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0_|A|1 SPL_IG2_0_|QA1 SPL_IG2_0_|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0_|A|P SPL_IG2_0_|A|MID_SERIES 0  2e-13
RSPL_IG2_0_|A|B SPL_IG2_0_|QA1 SPL_IG2_0_|A|MID_SHUNT  2.7439617672
LSPL_IG2_0_|A|RB SPL_IG2_0_|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0_|B|1 SPL_IG2_0_|QB1 SPL_IG2_0_|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0_|B|P SPL_IG2_0_|B|MID_SERIES 0  2e-13
RSPL_IG2_0_|B|B SPL_IG2_0_|QB1 SPL_IG2_0_|B|MID_SHUNT  2.7439617672
LSPL_IG2_0_|B|RB SPL_IG2_0_|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP3_0_|I_D1|B SPL_IP3_0_|D1 SPL_IP3_0_|I_D1|MID  2e-12
ISPL_IP3_0_|I_D1|B 0 SPL_IP3_0_|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP3_0_|I_D2|B SPL_IP3_0_|D2 SPL_IP3_0_|I_D2|MID  2e-12
ISPL_IP3_0_|I_D2|B 0 SPL_IP3_0_|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IP3_0_|I_Q1|B SPL_IP3_0_|QA1 SPL_IP3_0_|I_Q1|MID  2e-12
ISPL_IP3_0_|I_Q1|B 0 SPL_IP3_0_|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP3_0_|I_Q2|B SPL_IP3_0_|QB1 SPL_IP3_0_|I_Q2|MID  2e-12
ISPL_IP3_0_|I_Q2|B 0 SPL_IP3_0_|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IP3_0_|1|1 SPL_IP3_0_|D1 SPL_IP3_0_|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0_|1|P SPL_IP3_0_|1|MID_SERIES 0  2e-13
RSPL_IP3_0_|1|B SPL_IP3_0_|D1 SPL_IP3_0_|1|MID_SHUNT  2.7439617672
LSPL_IP3_0_|1|RB SPL_IP3_0_|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0_|2|1 SPL_IP3_0_|D2 SPL_IP3_0_|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0_|2|P SPL_IP3_0_|2|MID_SERIES 0  2e-13
RSPL_IP3_0_|2|B SPL_IP3_0_|D2 SPL_IP3_0_|2|MID_SHUNT  2.7439617672
LSPL_IP3_0_|2|RB SPL_IP3_0_|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0_|A|1 SPL_IP3_0_|QA1 SPL_IP3_0_|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0_|A|P SPL_IP3_0_|A|MID_SERIES 0  2e-13
RSPL_IP3_0_|A|B SPL_IP3_0_|QA1 SPL_IP3_0_|A|MID_SHUNT  2.7439617672
LSPL_IP3_0_|A|RB SPL_IP3_0_|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0_|B|1 SPL_IP3_0_|QB1 SPL_IP3_0_|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0_|B|P SPL_IP3_0_|B|MID_SERIES 0  2e-13
RSPL_IP3_0_|B|B SPL_IP3_0_|QB1 SPL_IP3_0_|B|MID_SHUNT  2.7439617672
LSPL_IP3_0_|B|RB SPL_IP3_0_|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01_|P|1 IP0_0_ _PG0_01_|P|A1  2.067833848e-12
L_PG0_01_|P|2 _PG0_01_|P|A1 _PG0_01_|P|A2  4.135667696e-12
L_PG0_01_|P|3 _PG0_01_|P|A3 _PG0_01_|P|A4  8.271335392e-12
L_PG0_01_|P|T T04_ _PG0_01_|P|T1  2.067833848e-12
L_PG0_01_|P|4 _PG0_01_|P|T1 _PG0_01_|P|T2  4.135667696e-12
L_PG0_01_|P|5 _PG0_01_|P|A4 _PG0_01_|P|Q1  4.135667696e-12
L_PG0_01_|P|6 _PG0_01_|P|Q1 P0_1_  2.067833848e-12
L_PG0_01_|G|1 IG0_0_TO0_ _PG0_01_|G|A1  2.067833848e-12
L_PG0_01_|G|2 _PG0_01_|G|A1 _PG0_01_|G|A2  4.135667696e-12
L_PG0_01_|G|3 _PG0_01_|G|A3 _PG0_01_|G|A4  8.271335392e-12
L_PG0_01_|G|T T04_ _PG0_01_|G|T1  2.067833848e-12
L_PG0_01_|G|4 _PG0_01_|G|T1 _PG0_01_|G|T2  4.135667696e-12
L_PG0_01_|G|5 _PG0_01_|G|A4 _PG0_01_|G|Q1  4.135667696e-12
L_PG0_01_|G|6 _PG0_01_|G|Q1 G0_1_  2.067833848e-12
L_PG1_01_|_SPL_G1|1 IG1_0_ _PG1_01_|_SPL_G1|D1  2e-12
L_PG1_01_|_SPL_G1|2 _PG1_01_|_SPL_G1|D1 _PG1_01_|_SPL_G1|D2  4.135667696e-12
L_PG1_01_|_SPL_G1|3 _PG1_01_|_SPL_G1|D2 _PG1_01_|_SPL_G1|JCT  9.84682784761905e-13
L_PG1_01_|_SPL_G1|4 _PG1_01_|_SPL_G1|JCT _PG1_01_|_SPL_G1|QA1  9.84682784761905e-13
L_PG1_01_|_SPL_G1|5 _PG1_01_|_SPL_G1|QA1 _PG1_01_|G1_COPY_1  2e-12
L_PG1_01_|_SPL_G1|6 _PG1_01_|_SPL_G1|JCT _PG1_01_|_SPL_G1|QB1  9.84682784761905e-13
L_PG1_01_|_SPL_G1|7 _PG1_01_|_SPL_G1|QB1 _PG1_01_|G1_COPY_2  2e-12
L_PG1_01_|_PG|A1 IP1_0_TO1_ _PG1_01_|_PG|A1  2.067833848e-12
L_PG1_01_|_PG|A2 _PG1_01_|_PG|A1 _PG1_01_|_PG|A2  4.135667696e-12
L_PG1_01_|_PG|A3 _PG1_01_|_PG|A3 _PG1_01_|_PG|Q3  1.2e-12
L_PG1_01_|_PG|B1 _PG1_01_|G1_COPY_1 _PG1_01_|_PG|B1  2.067833848e-12
L_PG1_01_|_PG|B2 _PG1_01_|_PG|B1 _PG1_01_|_PG|B2  4.135667696e-12
L_PG1_01_|_PG|B3 _PG1_01_|_PG|B3 _PG1_01_|_PG|Q3  1.2e-12
L_PG1_01_|_PG|Q3 _PG1_01_|_PG|Q3 _PG1_01_|_PG|Q2  4.135667696e-12
L_PG1_01_|_PG|Q2 _PG1_01_|_PG|Q2 _PG1_01_|_PG|Q1  4.135667696e-12
L_PG1_01_|_PG|Q1 _PG1_01_|_PG|Q1 _PG1_01_|PG  2.067833848e-12
L_PG1_01_|_GG|A1 IG0_0_TO1_ _PG1_01_|_GG|A1  2.067833848e-12
L_PG1_01_|_GG|A2 _PG1_01_|_GG|A1 _PG1_01_|_GG|A2  4.135667696e-12
L_PG1_01_|_GG|A3 _PG1_01_|_GG|A3 _PG1_01_|_GG|Q3  1.2e-12
L_PG1_01_|_GG|B1 _PG1_01_|G1_COPY_2 _PG1_01_|_GG|B1  2.067833848e-12
L_PG1_01_|_GG|B2 _PG1_01_|_GG|B1 _PG1_01_|_GG|B2  4.135667696e-12
L_PG1_01_|_GG|B3 _PG1_01_|_GG|B3 _PG1_01_|_GG|Q3  1.2e-12
L_PG1_01_|_GG|Q3 _PG1_01_|_GG|Q3 _PG1_01_|_GG|Q2  4.135667696e-12
L_PG1_01_|_GG|Q2 _PG1_01_|_GG|Q2 _PG1_01_|_GG|Q1  4.135667696e-12
L_PG1_01_|_GG|Q1 _PG1_01_|_GG|Q1 _PG1_01_|GG  2.067833848e-12
L_PG1_01_|_DFF_PG|1 _PG1_01_|PG _PG1_01_|_DFF_PG|A1  2.067833848e-12
L_PG1_01_|_DFF_PG|2 _PG1_01_|_DFF_PG|A1 _PG1_01_|_DFF_PG|A2  4.135667696e-12
L_PG1_01_|_DFF_PG|3 _PG1_01_|_DFF_PG|A3 _PG1_01_|_DFF_PG|A4  8.271335392e-12
L_PG1_01_|_DFF_PG|T T05_ _PG1_01_|_DFF_PG|T1  2.067833848e-12
L_PG1_01_|_DFF_PG|4 _PG1_01_|_DFF_PG|T1 _PG1_01_|_DFF_PG|T2  4.135667696e-12
L_PG1_01_|_DFF_PG|5 _PG1_01_|_DFF_PG|A4 _PG1_01_|_DFF_PG|Q1  4.135667696e-12
L_PG1_01_|_DFF_PG|6 _PG1_01_|_DFF_PG|Q1 _PG1_01_|PG_SYNC  2.067833848e-12
L_PG1_01_|_DFF_GG|1 _PG1_01_|GG _PG1_01_|_DFF_GG|A1  2.067833848e-12
L_PG1_01_|_DFF_GG|2 _PG1_01_|_DFF_GG|A1 _PG1_01_|_DFF_GG|A2  4.135667696e-12
L_PG1_01_|_DFF_GG|3 _PG1_01_|_DFF_GG|A3 _PG1_01_|_DFF_GG|A4  8.271335392e-12
L_PG1_01_|_DFF_GG|T T05_ _PG1_01_|_DFF_GG|T1  2.067833848e-12
L_PG1_01_|_DFF_GG|4 _PG1_01_|_DFF_GG|T1 _PG1_01_|_DFF_GG|T2  4.135667696e-12
L_PG1_01_|_DFF_GG|5 _PG1_01_|_DFF_GG|A4 _PG1_01_|_DFF_GG|Q1  4.135667696e-12
L_PG1_01_|_DFF_GG|6 _PG1_01_|_DFF_GG|Q1 _PG1_01_|GG_SYNC  2.067833848e-12
L_PG1_01_|_AND_G|A1 _PG1_01_|PG_SYNC _PG1_01_|_AND_G|A1  2.067833848e-12
L_PG1_01_|_AND_G|A2 _PG1_01_|_AND_G|A1 _PG1_01_|_AND_G|A2  4.135667696e-12
L_PG1_01_|_AND_G|A3 _PG1_01_|_AND_G|A3 _PG1_01_|_AND_G|Q3  1.2e-12
L_PG1_01_|_AND_G|B1 _PG1_01_|GG_SYNC _PG1_01_|_AND_G|B1  2.067833848e-12
L_PG1_01_|_AND_G|B2 _PG1_01_|_AND_G|B1 _PG1_01_|_AND_G|B2  4.135667696e-12
L_PG1_01_|_AND_G|B3 _PG1_01_|_AND_G|B3 _PG1_01_|_AND_G|Q3  1.2e-12
L_PG1_01_|_AND_G|Q3 _PG1_01_|_AND_G|Q3 _PG1_01_|_AND_G|Q2  4.135667696e-12
L_PG1_01_|_AND_G|Q2 _PG1_01_|_AND_G|Q2 _PG1_01_|_AND_G|Q1  4.135667696e-12
L_PG1_01_|_AND_G|Q1 _PG1_01_|_AND_G|Q1 G1_1_  2.067833848e-12
L_PG2_01_|P|1 IP2_0_TO2_ _PG2_01_|P|A1  2.067833848e-12
L_PG2_01_|P|2 _PG2_01_|P|A1 _PG2_01_|P|A2  4.135667696e-12
L_PG2_01_|P|3 _PG2_01_|P|A3 _PG2_01_|P|A4  8.271335392e-12
L_PG2_01_|P|T T06_ _PG2_01_|P|T1  2.067833848e-12
L_PG2_01_|P|4 _PG2_01_|P|T1 _PG2_01_|P|T2  4.135667696e-12
L_PG2_01_|P|5 _PG2_01_|P|A4 _PG2_01_|P|Q1  4.135667696e-12
L_PG2_01_|P|6 _PG2_01_|P|Q1 P2_1_  2.067833848e-12
L_PG2_01_|G|1 IG2_0_TO2_ _PG2_01_|G|A1  2.067833848e-12
L_PG2_01_|G|2 _PG2_01_|G|A1 _PG2_01_|G|A2  4.135667696e-12
L_PG2_01_|G|3 _PG2_01_|G|A3 _PG2_01_|G|A4  8.271335392e-12
L_PG2_01_|G|T T06_ _PG2_01_|G|T1  2.067833848e-12
L_PG2_01_|G|4 _PG2_01_|G|T1 _PG2_01_|G|T2  4.135667696e-12
L_PG2_01_|G|5 _PG2_01_|G|A4 _PG2_01_|G|Q1  4.135667696e-12
L_PG2_01_|G|6 _PG2_01_|G|Q1 G2_1_  2.067833848e-12
L_PG3_01_|_SPL_G1|1 IG3_0_ _PG3_01_|_SPL_G1|D1  2e-12
L_PG3_01_|_SPL_G1|2 _PG3_01_|_SPL_G1|D1 _PG3_01_|_SPL_G1|D2  4.135667696e-12
L_PG3_01_|_SPL_G1|3 _PG3_01_|_SPL_G1|D2 _PG3_01_|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_01_|_SPL_G1|4 _PG3_01_|_SPL_G1|JCT _PG3_01_|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_01_|_SPL_G1|5 _PG3_01_|_SPL_G1|QA1 _PG3_01_|G1_COPY_1  2e-12
L_PG3_01_|_SPL_G1|6 _PG3_01_|_SPL_G1|JCT _PG3_01_|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_01_|_SPL_G1|7 _PG3_01_|_SPL_G1|QB1 _PG3_01_|G1_COPY_2  2e-12
L_PG3_01_|_SPL_P1|1 IP3_0_TO1_ _PG3_01_|_SPL_P1|D1  2e-12
L_PG3_01_|_SPL_P1|2 _PG3_01_|_SPL_P1|D1 _PG3_01_|_SPL_P1|D2  4.135667696e-12
L_PG3_01_|_SPL_P1|3 _PG3_01_|_SPL_P1|D2 _PG3_01_|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_01_|_SPL_P1|4 _PG3_01_|_SPL_P1|JCT _PG3_01_|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_01_|_SPL_P1|5 _PG3_01_|_SPL_P1|QA1 _PG3_01_|P1_COPY_1  2e-12
L_PG3_01_|_SPL_P1|6 _PG3_01_|_SPL_P1|JCT _PG3_01_|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_01_|_SPL_P1|7 _PG3_01_|_SPL_P1|QB1 _PG3_01_|P1_COPY_2  2e-12
L_PG3_01_|_PG|A1 _PG3_01_|P1_COPY_1 _PG3_01_|_PG|A1  2.067833848e-12
L_PG3_01_|_PG|A2 _PG3_01_|_PG|A1 _PG3_01_|_PG|A2  4.135667696e-12
L_PG3_01_|_PG|A3 _PG3_01_|_PG|A3 _PG3_01_|_PG|Q3  1.2e-12
L_PG3_01_|_PG|B1 _PG3_01_|G1_COPY_1 _PG3_01_|_PG|B1  2.067833848e-12
L_PG3_01_|_PG|B2 _PG3_01_|_PG|B1 _PG3_01_|_PG|B2  4.135667696e-12
L_PG3_01_|_PG|B3 _PG3_01_|_PG|B3 _PG3_01_|_PG|Q3  1.2e-12
L_PG3_01_|_PG|Q3 _PG3_01_|_PG|Q3 _PG3_01_|_PG|Q2  4.135667696e-12
L_PG3_01_|_PG|Q2 _PG3_01_|_PG|Q2 _PG3_01_|_PG|Q1  4.135667696e-12
L_PG3_01_|_PG|Q1 _PG3_01_|_PG|Q1 _PG3_01_|PG  2.067833848e-12
L_PG3_01_|_GG|A1 IG2_0_TO3_ _PG3_01_|_GG|A1  2.067833848e-12
L_PG3_01_|_GG|A2 _PG3_01_|_GG|A1 _PG3_01_|_GG|A2  4.135667696e-12
L_PG3_01_|_GG|A3 _PG3_01_|_GG|A3 _PG3_01_|_GG|Q3  1.2e-12
L_PG3_01_|_GG|B1 _PG3_01_|G1_COPY_2 _PG3_01_|_GG|B1  2.067833848e-12
L_PG3_01_|_GG|B2 _PG3_01_|_GG|B1 _PG3_01_|_GG|B2  4.135667696e-12
L_PG3_01_|_GG|B3 _PG3_01_|_GG|B3 _PG3_01_|_GG|Q3  1.2e-12
L_PG3_01_|_GG|Q3 _PG3_01_|_GG|Q3 _PG3_01_|_GG|Q2  4.135667696e-12
L_PG3_01_|_GG|Q2 _PG3_01_|_GG|Q2 _PG3_01_|_GG|Q1  4.135667696e-12
L_PG3_01_|_GG|Q1 _PG3_01_|_GG|Q1 _PG3_01_|GG  2.067833848e-12
L_PG3_01_|_DFF_P0|1 IP2_0_TO3_ _PG3_01_|_DFF_P0|A1  2.067833848e-12
L_PG3_01_|_DFF_P0|2 _PG3_01_|_DFF_P0|A1 _PG3_01_|_DFF_P0|A2  4.135667696e-12
L_PG3_01_|_DFF_P0|3 _PG3_01_|_DFF_P0|A3 _PG3_01_|_DFF_P0|A4  8.271335392e-12
L_PG3_01_|_DFF_P0|T T07_ _PG3_01_|_DFF_P0|T1  2.067833848e-12
L_PG3_01_|_DFF_P0|4 _PG3_01_|_DFF_P0|T1 _PG3_01_|_DFF_P0|T2  4.135667696e-12
L_PG3_01_|_DFF_P0|5 _PG3_01_|_DFF_P0|A4 _PG3_01_|_DFF_P0|Q1  4.135667696e-12
L_PG3_01_|_DFF_P0|6 _PG3_01_|_DFF_P0|Q1 _PG3_01_|P0_SYNC  2.067833848e-12
L_PG3_01_|_DFF_P1|1 _PG3_01_|P1_COPY_2 _PG3_01_|_DFF_P1|A1  2.067833848e-12
L_PG3_01_|_DFF_P1|2 _PG3_01_|_DFF_P1|A1 _PG3_01_|_DFF_P1|A2  4.135667696e-12
L_PG3_01_|_DFF_P1|3 _PG3_01_|_DFF_P1|A3 _PG3_01_|_DFF_P1|A4  8.271335392e-12
L_PG3_01_|_DFF_P1|T T07_ _PG3_01_|_DFF_P1|T1  2.067833848e-12
L_PG3_01_|_DFF_P1|4 _PG3_01_|_DFF_P1|T1 _PG3_01_|_DFF_P1|T2  4.135667696e-12
L_PG3_01_|_DFF_P1|5 _PG3_01_|_DFF_P1|A4 _PG3_01_|_DFF_P1|Q1  4.135667696e-12
L_PG3_01_|_DFF_P1|6 _PG3_01_|_DFF_P1|Q1 _PG3_01_|P1_SYNC  2.067833848e-12
L_PG3_01_|_DFF_PG|1 _PG3_01_|PG _PG3_01_|_DFF_PG|A1  2.067833848e-12
L_PG3_01_|_DFF_PG|2 _PG3_01_|_DFF_PG|A1 _PG3_01_|_DFF_PG|A2  4.135667696e-12
L_PG3_01_|_DFF_PG|3 _PG3_01_|_DFF_PG|A3 _PG3_01_|_DFF_PG|A4  8.271335392e-12
L_PG3_01_|_DFF_PG|T T07_ _PG3_01_|_DFF_PG|T1  2.067833848e-12
L_PG3_01_|_DFF_PG|4 _PG3_01_|_DFF_PG|T1 _PG3_01_|_DFF_PG|T2  4.135667696e-12
L_PG3_01_|_DFF_PG|5 _PG3_01_|_DFF_PG|A4 _PG3_01_|_DFF_PG|Q1  4.135667696e-12
L_PG3_01_|_DFF_PG|6 _PG3_01_|_DFF_PG|Q1 _PG3_01_|PG_SYNC  2.067833848e-12
L_PG3_01_|_DFF_GG|1 _PG3_01_|GG _PG3_01_|_DFF_GG|A1  2.067833848e-12
L_PG3_01_|_DFF_GG|2 _PG3_01_|_DFF_GG|A1 _PG3_01_|_DFF_GG|A2  4.135667696e-12
L_PG3_01_|_DFF_GG|3 _PG3_01_|_DFF_GG|A3 _PG3_01_|_DFF_GG|A4  8.271335392e-12
L_PG3_01_|_DFF_GG|T T07_ _PG3_01_|_DFF_GG|T1  2.067833848e-12
L_PG3_01_|_DFF_GG|4 _PG3_01_|_DFF_GG|T1 _PG3_01_|_DFF_GG|T2  4.135667696e-12
L_PG3_01_|_DFF_GG|5 _PG3_01_|_DFF_GG|A4 _PG3_01_|_DFF_GG|Q1  4.135667696e-12
L_PG3_01_|_DFF_GG|6 _PG3_01_|_DFF_GG|Q1 _PG3_01_|GG_SYNC  2.067833848e-12
L_PG3_01_|_AND_G|A1 _PG3_01_|PG_SYNC _PG3_01_|_AND_G|A1  2.067833848e-12
L_PG3_01_|_AND_G|A2 _PG3_01_|_AND_G|A1 _PG3_01_|_AND_G|A2  4.135667696e-12
L_PG3_01_|_AND_G|A3 _PG3_01_|_AND_G|A3 _PG3_01_|_AND_G|Q3  1.2e-12
L_PG3_01_|_AND_G|B1 _PG3_01_|GG_SYNC _PG3_01_|_AND_G|B1  2.067833848e-12
L_PG3_01_|_AND_G|B2 _PG3_01_|_AND_G|B1 _PG3_01_|_AND_G|B2  4.135667696e-12
L_PG3_01_|_AND_G|B3 _PG3_01_|_AND_G|B3 _PG3_01_|_AND_G|Q3  1.2e-12
L_PG3_01_|_AND_G|Q3 _PG3_01_|_AND_G|Q3 _PG3_01_|_AND_G|Q2  4.135667696e-12
L_PG3_01_|_AND_G|Q2 _PG3_01_|_AND_G|Q2 _PG3_01_|_AND_G|Q1  4.135667696e-12
L_PG3_01_|_AND_G|Q1 _PG3_01_|_AND_G|Q1 G3_1_  2.067833848e-12
L_PG3_01_|_AND_P|A1 _PG3_01_|P0_SYNC _PG3_01_|_AND_P|A1  2.067833848e-12
L_PG3_01_|_AND_P|A2 _PG3_01_|_AND_P|A1 _PG3_01_|_AND_P|A2  4.135667696e-12
L_PG3_01_|_AND_P|A3 _PG3_01_|_AND_P|A3 _PG3_01_|_AND_P|Q3  1.2e-12
L_PG3_01_|_AND_P|B1 _PG3_01_|P1_SYNC _PG3_01_|_AND_P|B1  2.067833848e-12
L_PG3_01_|_AND_P|B2 _PG3_01_|_AND_P|B1 _PG3_01_|_AND_P|B2  4.135667696e-12
L_PG3_01_|_AND_P|B3 _PG3_01_|_AND_P|B3 _PG3_01_|_AND_P|Q3  1.2e-12
L_PG3_01_|_AND_P|Q3 _PG3_01_|_AND_P|Q3 _PG3_01_|_AND_P|Q2  4.135667696e-12
L_PG3_01_|_AND_P|Q2 _PG3_01_|_AND_P|Q2 _PG3_01_|_AND_P|Q1  4.135667696e-12
L_PG3_01_|_AND_P|Q1 _PG3_01_|_AND_P|Q1 P3_1_  2.067833848e-12
L_DFF_IP1_01_|I_1|B _DFF_IP1_01_|A1 _DFF_IP1_01_|I_1|MID  2e-12
I_DFF_IP1_01_|I_1|B 0 _DFF_IP1_01_|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01_|I_3|B _DFF_IP1_01_|A3 _DFF_IP1_01_|I_3|MID  2e-12
I_DFF_IP1_01_|I_3|B 0 _DFF_IP1_01_|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_01_|I_T|B _DFF_IP1_01_|T1 _DFF_IP1_01_|I_T|MID  2e-12
I_DFF_IP1_01_|I_T|B 0 _DFF_IP1_01_|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01_|I_6|B _DFF_IP1_01_|Q1 _DFF_IP1_01_|I_6|MID  2e-12
I_DFF_IP1_01_|I_6|B 0 _DFF_IP1_01_|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_01_|1|1 _DFF_IP1_01_|A1 _DFF_IP1_01_|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01_|1|P _DFF_IP1_01_|1|MID_SERIES 0  2e-13
R_DFF_IP1_01_|1|B _DFF_IP1_01_|A1 _DFF_IP1_01_|1|MID_SHUNT  2.7439617672
L_DFF_IP1_01_|1|RB _DFF_IP1_01_|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01_|23|1 _DFF_IP1_01_|A2 _DFF_IP1_01_|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01_|23|B _DFF_IP1_01_|A2 _DFF_IP1_01_|23|MID_SHUNT  3.84154647408
L_DFF_IP1_01_|23|RB _DFF_IP1_01_|23|MID_SHUNT _DFF_IP1_01_|A3  2.1704737578552e-12
B_DFF_IP1_01_|3|1 _DFF_IP1_01_|A3 _DFF_IP1_01_|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01_|3|P _DFF_IP1_01_|3|MID_SERIES 0  2e-13
R_DFF_IP1_01_|3|B _DFF_IP1_01_|A3 _DFF_IP1_01_|3|MID_SHUNT  2.7439617672
L_DFF_IP1_01_|3|RB _DFF_IP1_01_|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01_|4|1 _DFF_IP1_01_|A4 _DFF_IP1_01_|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01_|4|P _DFF_IP1_01_|4|MID_SERIES 0  2e-13
R_DFF_IP1_01_|4|B _DFF_IP1_01_|A4 _DFF_IP1_01_|4|MID_SHUNT  2.7439617672
L_DFF_IP1_01_|4|RB _DFF_IP1_01_|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01_|T|1 _DFF_IP1_01_|T1 _DFF_IP1_01_|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01_|T|P _DFF_IP1_01_|T|MID_SERIES 0  2e-13
R_DFF_IP1_01_|T|B _DFF_IP1_01_|T1 _DFF_IP1_01_|T|MID_SHUNT  2.7439617672
L_DFF_IP1_01_|T|RB _DFF_IP1_01_|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01_|45|1 _DFF_IP1_01_|T2 _DFF_IP1_01_|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01_|45|B _DFF_IP1_01_|T2 _DFF_IP1_01_|45|MID_SHUNT  3.84154647408
L_DFF_IP1_01_|45|RB _DFF_IP1_01_|45|MID_SHUNT _DFF_IP1_01_|A4  2.1704737578552e-12
B_DFF_IP1_01_|6|1 _DFF_IP1_01_|Q1 _DFF_IP1_01_|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01_|6|P _DFF_IP1_01_|6|MID_SERIES 0  2e-13
R_DFF_IP1_01_|6|B _DFF_IP1_01_|Q1 _DFF_IP1_01_|6|MID_SHUNT  2.7439617672
L_DFF_IP1_01_|6|RB _DFF_IP1_01_|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_01_|I_1|B _DFF_IP2_01_|A1 _DFF_IP2_01_|I_1|MID  2e-12
I_DFF_IP2_01_|I_1|B 0 _DFF_IP2_01_|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01_|I_3|B _DFF_IP2_01_|A3 _DFF_IP2_01_|I_3|MID  2e-12
I_DFF_IP2_01_|I_3|B 0 _DFF_IP2_01_|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_01_|I_T|B _DFF_IP2_01_|T1 _DFF_IP2_01_|I_T|MID  2e-12
I_DFF_IP2_01_|I_T|B 0 _DFF_IP2_01_|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01_|I_6|B _DFF_IP2_01_|Q1 _DFF_IP2_01_|I_6|MID  2e-12
I_DFF_IP2_01_|I_6|B 0 _DFF_IP2_01_|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_01_|1|1 _DFF_IP2_01_|A1 _DFF_IP2_01_|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01_|1|P _DFF_IP2_01_|1|MID_SERIES 0  2e-13
R_DFF_IP2_01_|1|B _DFF_IP2_01_|A1 _DFF_IP2_01_|1|MID_SHUNT  2.7439617672
L_DFF_IP2_01_|1|RB _DFF_IP2_01_|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01_|23|1 _DFF_IP2_01_|A2 _DFF_IP2_01_|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01_|23|B _DFF_IP2_01_|A2 _DFF_IP2_01_|23|MID_SHUNT  3.84154647408
L_DFF_IP2_01_|23|RB _DFF_IP2_01_|23|MID_SHUNT _DFF_IP2_01_|A3  2.1704737578552e-12
B_DFF_IP2_01_|3|1 _DFF_IP2_01_|A3 _DFF_IP2_01_|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01_|3|P _DFF_IP2_01_|3|MID_SERIES 0  2e-13
R_DFF_IP2_01_|3|B _DFF_IP2_01_|A3 _DFF_IP2_01_|3|MID_SHUNT  2.7439617672
L_DFF_IP2_01_|3|RB _DFF_IP2_01_|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01_|4|1 _DFF_IP2_01_|A4 _DFF_IP2_01_|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01_|4|P _DFF_IP2_01_|4|MID_SERIES 0  2e-13
R_DFF_IP2_01_|4|B _DFF_IP2_01_|A4 _DFF_IP2_01_|4|MID_SHUNT  2.7439617672
L_DFF_IP2_01_|4|RB _DFF_IP2_01_|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01_|T|1 _DFF_IP2_01_|T1 _DFF_IP2_01_|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01_|T|P _DFF_IP2_01_|T|MID_SERIES 0  2e-13
R_DFF_IP2_01_|T|B _DFF_IP2_01_|T1 _DFF_IP2_01_|T|MID_SHUNT  2.7439617672
L_DFF_IP2_01_|T|RB _DFF_IP2_01_|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01_|45|1 _DFF_IP2_01_|T2 _DFF_IP2_01_|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01_|45|B _DFF_IP2_01_|T2 _DFF_IP2_01_|45|MID_SHUNT  3.84154647408
L_DFF_IP2_01_|45|RB _DFF_IP2_01_|45|MID_SHUNT _DFF_IP2_01_|A4  2.1704737578552e-12
B_DFF_IP2_01_|6|1 _DFF_IP2_01_|Q1 _DFF_IP2_01_|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01_|6|P _DFF_IP2_01_|6|MID_SERIES 0  2e-13
R_DFF_IP2_01_|6|B _DFF_IP2_01_|Q1 _DFF_IP2_01_|6|MID_SHUNT  2.7439617672
L_DFF_IP2_01_|6|RB _DFF_IP2_01_|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_01_|I_1|B _DFF_IP3_01_|A1 _DFF_IP3_01_|I_1|MID  2e-12
I_DFF_IP3_01_|I_1|B 0 _DFF_IP3_01_|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01_|I_3|B _DFF_IP3_01_|A3 _DFF_IP3_01_|I_3|MID  2e-12
I_DFF_IP3_01_|I_3|B 0 _DFF_IP3_01_|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_01_|I_T|B _DFF_IP3_01_|T1 _DFF_IP3_01_|I_T|MID  2e-12
I_DFF_IP3_01_|I_T|B 0 _DFF_IP3_01_|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01_|I_6|B _DFF_IP3_01_|Q1 _DFF_IP3_01_|I_6|MID  2e-12
I_DFF_IP3_01_|I_6|B 0 _DFF_IP3_01_|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_01_|1|1 _DFF_IP3_01_|A1 _DFF_IP3_01_|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01_|1|P _DFF_IP3_01_|1|MID_SERIES 0  2e-13
R_DFF_IP3_01_|1|B _DFF_IP3_01_|A1 _DFF_IP3_01_|1|MID_SHUNT  2.7439617672
L_DFF_IP3_01_|1|RB _DFF_IP3_01_|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01_|23|1 _DFF_IP3_01_|A2 _DFF_IP3_01_|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01_|23|B _DFF_IP3_01_|A2 _DFF_IP3_01_|23|MID_SHUNT  3.84154647408
L_DFF_IP3_01_|23|RB _DFF_IP3_01_|23|MID_SHUNT _DFF_IP3_01_|A3  2.1704737578552e-12
B_DFF_IP3_01_|3|1 _DFF_IP3_01_|A3 _DFF_IP3_01_|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01_|3|P _DFF_IP3_01_|3|MID_SERIES 0  2e-13
R_DFF_IP3_01_|3|B _DFF_IP3_01_|A3 _DFF_IP3_01_|3|MID_SHUNT  2.7439617672
L_DFF_IP3_01_|3|RB _DFF_IP3_01_|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01_|4|1 _DFF_IP3_01_|A4 _DFF_IP3_01_|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01_|4|P _DFF_IP3_01_|4|MID_SERIES 0  2e-13
R_DFF_IP3_01_|4|B _DFF_IP3_01_|A4 _DFF_IP3_01_|4|MID_SHUNT  2.7439617672
L_DFF_IP3_01_|4|RB _DFF_IP3_01_|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01_|T|1 _DFF_IP3_01_|T1 _DFF_IP3_01_|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01_|T|P _DFF_IP3_01_|T|MID_SERIES 0  2e-13
R_DFF_IP3_01_|T|B _DFF_IP3_01_|T1 _DFF_IP3_01_|T|MID_SHUNT  2.7439617672
L_DFF_IP3_01_|T|RB _DFF_IP3_01_|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01_|45|1 _DFF_IP3_01_|T2 _DFF_IP3_01_|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01_|45|B _DFF_IP3_01_|T2 _DFF_IP3_01_|45|MID_SHUNT  3.84154647408
L_DFF_IP3_01_|45|RB _DFF_IP3_01_|45|MID_SHUNT _DFF_IP3_01_|A4  2.1704737578552e-12
B_DFF_IP3_01_|6|1 _DFF_IP3_01_|Q1 _DFF_IP3_01_|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01_|6|P _DFF_IP3_01_|6|MID_SERIES 0  2e-13
R_DFF_IP3_01_|6|B _DFF_IP3_01_|Q1 _DFF_IP3_01_|6|MID_SHUNT  2.7439617672
L_DFF_IP3_01_|6|RB _DFF_IP3_01_|6|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1_|SPL1|1 G1_1_ SPL_G1_1_|SPL1|D1  2e-12
LSPL_G1_1_|SPL1|2 SPL_G1_1_|SPL1|D1 SPL_G1_1_|SPL1|D2  4.135667696e-12
LSPL_G1_1_|SPL1|3 SPL_G1_1_|SPL1|D2 SPL_G1_1_|SPL1|JCT  9.84682784761905e-13
LSPL_G1_1_|SPL1|4 SPL_G1_1_|SPL1|JCT SPL_G1_1_|SPL1|QA1  9.84682784761905e-13
LSPL_G1_1_|SPL1|5 SPL_G1_1_|SPL1|QA1 G1_1_TO1_  2e-12
LSPL_G1_1_|SPL1|6 SPL_G1_1_|SPL1|JCT SPL_G1_1_|SPL1|QB1  9.84682784761905e-13
LSPL_G1_1_|SPL1|7 SPL_G1_1_|SPL1|QB1 SPL_G1_1_|QTMP  2e-12
LSPL_G1_1_|SPL2|1 SPL_G1_1_|QTMP SPL_G1_1_|SPL2|D1  2e-12
LSPL_G1_1_|SPL2|2 SPL_G1_1_|SPL2|D1 SPL_G1_1_|SPL2|D2  4.135667696e-12
LSPL_G1_1_|SPL2|3 SPL_G1_1_|SPL2|D2 SPL_G1_1_|SPL2|JCT  9.84682784761905e-13
LSPL_G1_1_|SPL2|4 SPL_G1_1_|SPL2|JCT SPL_G1_1_|SPL2|QA1  9.84682784761905e-13
LSPL_G1_1_|SPL2|5 SPL_G1_1_|SPL2|QA1 G1_1_TO2_  2e-12
LSPL_G1_1_|SPL2|6 SPL_G1_1_|SPL2|JCT SPL_G1_1_|SPL2|QB1  9.84682784761905e-13
LSPL_G1_1_|SPL2|7 SPL_G1_1_|SPL2|QB1 G1_1_TO3_  2e-12
LI0_|_SPL_A|I_D1|B I0_|_SPL_A|D1 I0_|_SPL_A|I_D1|MID  2e-12
II0_|_SPL_A|I_D1|B 0 I0_|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_SPL_A|I_D2|B I0_|_SPL_A|D2 I0_|_SPL_A|I_D2|MID  2e-12
II0_|_SPL_A|I_D2|B 0 I0_|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI0_|_SPL_A|I_Q1|B I0_|_SPL_A|QA1 I0_|_SPL_A|I_Q1|MID  2e-12
II0_|_SPL_A|I_Q1|B 0 I0_|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_SPL_A|I_Q2|B I0_|_SPL_A|QB1 I0_|_SPL_A|I_Q2|MID  2e-12
II0_|_SPL_A|I_Q2|B 0 I0_|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI0_|_SPL_A|1|1 I0_|_SPL_A|D1 I0_|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_A|1|P I0_|_SPL_A|1|MID_SERIES 0  2e-13
RI0_|_SPL_A|1|B I0_|_SPL_A|D1 I0_|_SPL_A|1|MID_SHUNT  2.7439617672
LI0_|_SPL_A|1|RB I0_|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI0_|_SPL_A|2|1 I0_|_SPL_A|D2 I0_|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_A|2|P I0_|_SPL_A|2|MID_SERIES 0  2e-13
RI0_|_SPL_A|2|B I0_|_SPL_A|D2 I0_|_SPL_A|2|MID_SHUNT  2.7439617672
LI0_|_SPL_A|2|RB I0_|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI0_|_SPL_A|A|1 I0_|_SPL_A|QA1 I0_|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_A|A|P I0_|_SPL_A|A|MID_SERIES 0  2e-13
RI0_|_SPL_A|A|B I0_|_SPL_A|QA1 I0_|_SPL_A|A|MID_SHUNT  2.7439617672
LI0_|_SPL_A|A|RB I0_|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI0_|_SPL_A|B|1 I0_|_SPL_A|QB1 I0_|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_A|B|P I0_|_SPL_A|B|MID_SERIES 0  2e-13
RI0_|_SPL_A|B|B I0_|_SPL_A|QB1 I0_|_SPL_A|B|MID_SHUNT  2.7439617672
LI0_|_SPL_A|B|RB I0_|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI0_|_SPL_B|I_D1|B I0_|_SPL_B|D1 I0_|_SPL_B|I_D1|MID  2e-12
II0_|_SPL_B|I_D1|B 0 I0_|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_SPL_B|I_D2|B I0_|_SPL_B|D2 I0_|_SPL_B|I_D2|MID  2e-12
II0_|_SPL_B|I_D2|B 0 I0_|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI0_|_SPL_B|I_Q1|B I0_|_SPL_B|QA1 I0_|_SPL_B|I_Q1|MID  2e-12
II0_|_SPL_B|I_Q1|B 0 I0_|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_SPL_B|I_Q2|B I0_|_SPL_B|QB1 I0_|_SPL_B|I_Q2|MID  2e-12
II0_|_SPL_B|I_Q2|B 0 I0_|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI0_|_SPL_B|1|1 I0_|_SPL_B|D1 I0_|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_B|1|P I0_|_SPL_B|1|MID_SERIES 0  2e-13
RI0_|_SPL_B|1|B I0_|_SPL_B|D1 I0_|_SPL_B|1|MID_SHUNT  2.7439617672
LI0_|_SPL_B|1|RB I0_|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI0_|_SPL_B|2|1 I0_|_SPL_B|D2 I0_|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_B|2|P I0_|_SPL_B|2|MID_SERIES 0  2e-13
RI0_|_SPL_B|2|B I0_|_SPL_B|D2 I0_|_SPL_B|2|MID_SHUNT  2.7439617672
LI0_|_SPL_B|2|RB I0_|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI0_|_SPL_B|A|1 I0_|_SPL_B|QA1 I0_|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_B|A|P I0_|_SPL_B|A|MID_SERIES 0  2e-13
RI0_|_SPL_B|A|B I0_|_SPL_B|QA1 I0_|_SPL_B|A|MID_SHUNT  2.7439617672
LI0_|_SPL_B|A|RB I0_|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI0_|_SPL_B|B|1 I0_|_SPL_B|QB1 I0_|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI0_|_SPL_B|B|P I0_|_SPL_B|B|MID_SERIES 0  2e-13
RI0_|_SPL_B|B|B I0_|_SPL_B|QB1 I0_|_SPL_B|B|MID_SHUNT  2.7439617672
LI0_|_SPL_B|B|RB I0_|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI0_|_DFF_A|I_1|B I0_|_DFF_A|A1 I0_|_DFF_A|I_1|MID  2e-12
II0_|_DFF_A|I_1|B 0 I0_|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_DFF_A|I_3|B I0_|_DFF_A|A3 I0_|_DFF_A|I_3|MID  2e-12
II0_|_DFF_A|I_3|B 0 I0_|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0_|_DFF_A|I_T|B I0_|_DFF_A|T1 I0_|_DFF_A|I_T|MID  2e-12
II0_|_DFF_A|I_T|B 0 I0_|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0_|_DFF_A|I_6|B I0_|_DFF_A|Q1 I0_|_DFF_A|I_6|MID  2e-12
II0_|_DFF_A|I_6|B 0 I0_|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0_|_DFF_A|1|1 I0_|_DFF_A|A1 I0_|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_A|1|P I0_|_DFF_A|1|MID_SERIES 0  2e-13
RI0_|_DFF_A|1|B I0_|_DFF_A|A1 I0_|_DFF_A|1|MID_SHUNT  2.7439617672
LI0_|_DFF_A|1|RB I0_|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_A|23|1 I0_|_DFF_A|A2 I0_|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI0_|_DFF_A|23|B I0_|_DFF_A|A2 I0_|_DFF_A|23|MID_SHUNT  3.84154647408
LI0_|_DFF_A|23|RB I0_|_DFF_A|23|MID_SHUNT I0_|_DFF_A|A3  2.1704737578552e-12
BI0_|_DFF_A|3|1 I0_|_DFF_A|A3 I0_|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_A|3|P I0_|_DFF_A|3|MID_SERIES 0  2e-13
RI0_|_DFF_A|3|B I0_|_DFF_A|A3 I0_|_DFF_A|3|MID_SHUNT  2.7439617672
LI0_|_DFF_A|3|RB I0_|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_A|4|1 I0_|_DFF_A|A4 I0_|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_A|4|P I0_|_DFF_A|4|MID_SERIES 0  2e-13
RI0_|_DFF_A|4|B I0_|_DFF_A|A4 I0_|_DFF_A|4|MID_SHUNT  2.7439617672
LI0_|_DFF_A|4|RB I0_|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_A|T|1 I0_|_DFF_A|T1 I0_|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_A|T|P I0_|_DFF_A|T|MID_SERIES 0  2e-13
RI0_|_DFF_A|T|B I0_|_DFF_A|T1 I0_|_DFF_A|T|MID_SHUNT  2.7439617672
LI0_|_DFF_A|T|RB I0_|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_A|45|1 I0_|_DFF_A|T2 I0_|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI0_|_DFF_A|45|B I0_|_DFF_A|T2 I0_|_DFF_A|45|MID_SHUNT  3.84154647408
LI0_|_DFF_A|45|RB I0_|_DFF_A|45|MID_SHUNT I0_|_DFF_A|A4  2.1704737578552e-12
BI0_|_DFF_A|6|1 I0_|_DFF_A|Q1 I0_|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_A|6|P I0_|_DFF_A|6|MID_SERIES 0  2e-13
RI0_|_DFF_A|6|B I0_|_DFF_A|Q1 I0_|_DFF_A|6|MID_SHUNT  2.7439617672
LI0_|_DFF_A|6|RB I0_|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI0_|_DFF_B|I_1|B I0_|_DFF_B|A1 I0_|_DFF_B|I_1|MID  2e-12
II0_|_DFF_B|I_1|B 0 I0_|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_DFF_B|I_3|B I0_|_DFF_B|A3 I0_|_DFF_B|I_3|MID  2e-12
II0_|_DFF_B|I_3|B 0 I0_|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0_|_DFF_B|I_T|B I0_|_DFF_B|T1 I0_|_DFF_B|I_T|MID  2e-12
II0_|_DFF_B|I_T|B 0 I0_|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0_|_DFF_B|I_6|B I0_|_DFF_B|Q1 I0_|_DFF_B|I_6|MID  2e-12
II0_|_DFF_B|I_6|B 0 I0_|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0_|_DFF_B|1|1 I0_|_DFF_B|A1 I0_|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_B|1|P I0_|_DFF_B|1|MID_SERIES 0  2e-13
RI0_|_DFF_B|1|B I0_|_DFF_B|A1 I0_|_DFF_B|1|MID_SHUNT  2.7439617672
LI0_|_DFF_B|1|RB I0_|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_B|23|1 I0_|_DFF_B|A2 I0_|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI0_|_DFF_B|23|B I0_|_DFF_B|A2 I0_|_DFF_B|23|MID_SHUNT  3.84154647408
LI0_|_DFF_B|23|RB I0_|_DFF_B|23|MID_SHUNT I0_|_DFF_B|A3  2.1704737578552e-12
BI0_|_DFF_B|3|1 I0_|_DFF_B|A3 I0_|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_B|3|P I0_|_DFF_B|3|MID_SERIES 0  2e-13
RI0_|_DFF_B|3|B I0_|_DFF_B|A3 I0_|_DFF_B|3|MID_SHUNT  2.7439617672
LI0_|_DFF_B|3|RB I0_|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_B|4|1 I0_|_DFF_B|A4 I0_|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_B|4|P I0_|_DFF_B|4|MID_SERIES 0  2e-13
RI0_|_DFF_B|4|B I0_|_DFF_B|A4 I0_|_DFF_B|4|MID_SHUNT  2.7439617672
LI0_|_DFF_B|4|RB I0_|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_B|T|1 I0_|_DFF_B|T1 I0_|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_B|T|P I0_|_DFF_B|T|MID_SERIES 0  2e-13
RI0_|_DFF_B|T|B I0_|_DFF_B|T1 I0_|_DFF_B|T|MID_SHUNT  2.7439617672
LI0_|_DFF_B|T|RB I0_|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI0_|_DFF_B|45|1 I0_|_DFF_B|T2 I0_|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI0_|_DFF_B|45|B I0_|_DFF_B|T2 I0_|_DFF_B|45|MID_SHUNT  3.84154647408
LI0_|_DFF_B|45|RB I0_|_DFF_B|45|MID_SHUNT I0_|_DFF_B|A4  2.1704737578552e-12
BI0_|_DFF_B|6|1 I0_|_DFF_B|Q1 I0_|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI0_|_DFF_B|6|P I0_|_DFF_B|6|MID_SERIES 0  2e-13
RI0_|_DFF_B|6|B I0_|_DFF_B|Q1 I0_|_DFF_B|6|MID_SHUNT  2.7439617672
LI0_|_DFF_B|6|RB I0_|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI0_|_XOR|I_A1|B I0_|_XOR|A1 I0_|_XOR|I_A1|MID  2e-12
II0_|_XOR|I_A1|B 0 I0_|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_XOR|I_A3|B I0_|_XOR|A3 I0_|_XOR|I_A3|MID  2e-12
II0_|_XOR|I_A3|B 0 I0_|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI0_|_XOR|I_B1|B I0_|_XOR|B1 I0_|_XOR|I_B1|MID  2e-12
II0_|_XOR|I_B1|B 0 I0_|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_XOR|I_B3|B I0_|_XOR|B3 I0_|_XOR|I_B3|MID  2e-12
II0_|_XOR|I_B3|B 0 I0_|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI0_|_XOR|I_Q1|B I0_|_XOR|Q1 I0_|_XOR|I_Q1|MID  2e-12
II0_|_XOR|I_Q1|B 0 I0_|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0_|_XOR|A1|1 I0_|_XOR|A1 I0_|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|A1|P I0_|_XOR|A1|MID_SERIES 0  5e-13
RI0_|_XOR|A1|B I0_|_XOR|A1 I0_|_XOR|A1|MID_SHUNT  2.7439617672
LI0_|_XOR|A1|RB I0_|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI0_|_XOR|A2|1 I0_|_XOR|A2 I0_|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|A2|P I0_|_XOR|A2|MID_SERIES 0  5e-13
RI0_|_XOR|A2|B I0_|_XOR|A2 I0_|_XOR|A2|MID_SHUNT  2.7439617672
LI0_|_XOR|A2|RB I0_|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI0_|_XOR|A3|1 I0_|_XOR|A2 I0_|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|A3|P I0_|_XOR|A3|MID_SERIES I0_|_XOR|A3  1.2e-12
RI0_|_XOR|A3|B I0_|_XOR|A2 I0_|_XOR|A3|MID_SHUNT  2.7439617672
LI0_|_XOR|A3|RB I0_|_XOR|A3|MID_SHUNT I0_|_XOR|A3  2.050338398468e-12
BI0_|_XOR|B1|1 I0_|_XOR|B1 I0_|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|B1|P I0_|_XOR|B1|MID_SERIES 0  5e-13
RI0_|_XOR|B1|B I0_|_XOR|B1 I0_|_XOR|B1|MID_SHUNT  2.7439617672
LI0_|_XOR|B1|RB I0_|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI0_|_XOR|B2|1 I0_|_XOR|B2 I0_|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|B2|P I0_|_XOR|B2|MID_SERIES 0  5e-13
RI0_|_XOR|B2|B I0_|_XOR|B2 I0_|_XOR|B2|MID_SHUNT  2.7439617672
LI0_|_XOR|B2|RB I0_|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI0_|_XOR|B3|1 I0_|_XOR|B2 I0_|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|B3|P I0_|_XOR|B3|MID_SERIES I0_|_XOR|B3  1.2e-12
RI0_|_XOR|B3|B I0_|_XOR|B2 I0_|_XOR|B3|MID_SHUNT  2.7439617672
LI0_|_XOR|B3|RB I0_|_XOR|B3|MID_SHUNT I0_|_XOR|B3  2.050338398468e-12
BI0_|_XOR|T1|1 I0_|_XOR|T1 I0_|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|T1|P I0_|_XOR|T1|MID_SERIES 0  5e-13
RI0_|_XOR|T1|B I0_|_XOR|T1 I0_|_XOR|T1|MID_SHUNT  2.7439617672
LI0_|_XOR|T1|RB I0_|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI0_|_XOR|T2|1 I0_|_XOR|T2 I0_|_XOR|ABTQ JJMIT AREA=2.0
RI0_|_XOR|T2|B I0_|_XOR|T2 I0_|_XOR|T2|MID_SHUNT  3.429952209
LI0_|_XOR|T2|RB I0_|_XOR|T2|MID_SHUNT I0_|_XOR|ABTQ  2.437922998085e-12
BI0_|_XOR|AB|1 I0_|_XOR|AB I0_|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI0_|_XOR|AB|P I0_|_XOR|AB|MID_SERIES I0_|_XOR|ABTQ  1.2e-12
RI0_|_XOR|AB|B I0_|_XOR|AB I0_|_XOR|AB|MID_SHUNT  3.429952209
LI0_|_XOR|AB|RB I0_|_XOR|AB|MID_SHUNT I0_|_XOR|ABTQ  2.437922998085e-12
BI0_|_XOR|ABTQ|1 I0_|_XOR|ABTQ I0_|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|ABTQ|P I0_|_XOR|ABTQ|MID_SERIES 0  5e-13
RI0_|_XOR|ABTQ|B I0_|_XOR|ABTQ I0_|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI0_|_XOR|ABTQ|RB I0_|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI0_|_XOR|Q1|1 I0_|_XOR|Q1 I0_|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI0_|_XOR|Q1|P I0_|_XOR|Q1|MID_SERIES 0  5e-13
RI0_|_XOR|Q1|B I0_|_XOR|Q1 I0_|_XOR|Q1|MID_SHUNT  2.7439617672
LI0_|_XOR|Q1|RB I0_|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI0_|_AND|I_A1|B I0_|_AND|A1 I0_|_AND|I_A1|MID  2e-12
II0_|_AND|I_A1|B 0 I0_|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_AND|I_B1|B I0_|_AND|B1 I0_|_AND|I_B1|MID  2e-12
II0_|_AND|I_B1|B 0 I0_|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0_|_AND|I_Q3|B I0_|_AND|Q3 I0_|_AND|I_Q3|MID  2e-12
II0_|_AND|I_Q3|B 0 I0_|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0_|_AND|I_Q2|B I0_|_AND|Q2 I0_|_AND|I_Q2|MID  2e-12
II0_|_AND|I_Q2|B 0 I0_|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0_|_AND|I_Q1|B I0_|_AND|Q1 I0_|_AND|I_Q1|MID  2e-12
II0_|_AND|I_Q1|B 0 I0_|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0_|_AND|A1|1 I0_|_AND|A1 I0_|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0_|_AND|A1|P I0_|_AND|A1|MID_SERIES 0  2e-13
RI0_|_AND|A1|B I0_|_AND|A1 I0_|_AND|A1|MID_SHUNT  2.7439617672
LI0_|_AND|A1|RB I0_|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0_|_AND|A2|1 I0_|_AND|A2 I0_|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0_|_AND|A2|P I0_|_AND|A2|MID_SERIES 0  2e-13
RI0_|_AND|A2|B I0_|_AND|A2 I0_|_AND|A2|MID_SHUNT  2.7439617672
LI0_|_AND|A2|RB I0_|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0_|_AND|A12|1 I0_|_AND|A2 I0_|_AND|A3 JJMIT AREA=1.7857142857142858
RI0_|_AND|A12|B I0_|_AND|A2 I0_|_AND|A12|MID_SHUNT  3.84154647408
LI0_|_AND|A12|RB I0_|_AND|A12|MID_SHUNT I0_|_AND|A3  2.1704737578552e-12
BI0_|_AND|B1|1 I0_|_AND|B1 I0_|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0_|_AND|B1|P I0_|_AND|B1|MID_SERIES 0  2e-13
RI0_|_AND|B1|B I0_|_AND|B1 I0_|_AND|B1|MID_SHUNT  2.7439617672
LI0_|_AND|B1|RB I0_|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0_|_AND|B2|1 I0_|_AND|B2 I0_|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0_|_AND|B2|P I0_|_AND|B2|MID_SERIES 0  2e-13
RI0_|_AND|B2|B I0_|_AND|B2 I0_|_AND|B2|MID_SHUNT  2.7439617672
LI0_|_AND|B2|RB I0_|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0_|_AND|B12|1 I0_|_AND|B2 I0_|_AND|B3 JJMIT AREA=1.7857142857142858
RI0_|_AND|B12|B I0_|_AND|B2 I0_|_AND|B12|MID_SHUNT  3.84154647408
LI0_|_AND|B12|RB I0_|_AND|B12|MID_SHUNT I0_|_AND|B3  2.1704737578552e-12
BI0_|_AND|Q2|1 I0_|_AND|Q2 I0_|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0_|_AND|Q2|P I0_|_AND|Q2|MID_SERIES 0  2e-13
RI0_|_AND|Q2|B I0_|_AND|Q2 I0_|_AND|Q2|MID_SHUNT  2.7439617672
LI0_|_AND|Q2|RB I0_|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0_|_AND|Q1|1 I0_|_AND|Q1 I0_|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0_|_AND|Q1|P I0_|_AND|Q1|MID_SERIES 0  2e-13
RI0_|_AND|Q1|B I0_|_AND|Q1 I0_|_AND|Q1|MID_SHUNT  2.7439617672
LI0_|_AND|Q1|RB I0_|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1_|_SPL_A|I_D1|B I1_|_SPL_A|D1 I1_|_SPL_A|I_D1|MID  2e-12
II1_|_SPL_A|I_D1|B 0 I1_|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_SPL_A|I_D2|B I1_|_SPL_A|D2 I1_|_SPL_A|I_D2|MID  2e-12
II1_|_SPL_A|I_D2|B 0 I1_|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI1_|_SPL_A|I_Q1|B I1_|_SPL_A|QA1 I1_|_SPL_A|I_Q1|MID  2e-12
II1_|_SPL_A|I_Q1|B 0 I1_|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_SPL_A|I_Q2|B I1_|_SPL_A|QB1 I1_|_SPL_A|I_Q2|MID  2e-12
II1_|_SPL_A|I_Q2|B 0 I1_|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI1_|_SPL_A|1|1 I1_|_SPL_A|D1 I1_|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_A|1|P I1_|_SPL_A|1|MID_SERIES 0  2e-13
RI1_|_SPL_A|1|B I1_|_SPL_A|D1 I1_|_SPL_A|1|MID_SHUNT  2.7439617672
LI1_|_SPL_A|1|RB I1_|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI1_|_SPL_A|2|1 I1_|_SPL_A|D2 I1_|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_A|2|P I1_|_SPL_A|2|MID_SERIES 0  2e-13
RI1_|_SPL_A|2|B I1_|_SPL_A|D2 I1_|_SPL_A|2|MID_SHUNT  2.7439617672
LI1_|_SPL_A|2|RB I1_|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI1_|_SPL_A|A|1 I1_|_SPL_A|QA1 I1_|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_A|A|P I1_|_SPL_A|A|MID_SERIES 0  2e-13
RI1_|_SPL_A|A|B I1_|_SPL_A|QA1 I1_|_SPL_A|A|MID_SHUNT  2.7439617672
LI1_|_SPL_A|A|RB I1_|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI1_|_SPL_A|B|1 I1_|_SPL_A|QB1 I1_|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_A|B|P I1_|_SPL_A|B|MID_SERIES 0  2e-13
RI1_|_SPL_A|B|B I1_|_SPL_A|QB1 I1_|_SPL_A|B|MID_SHUNT  2.7439617672
LI1_|_SPL_A|B|RB I1_|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI1_|_SPL_B|I_D1|B I1_|_SPL_B|D1 I1_|_SPL_B|I_D1|MID  2e-12
II1_|_SPL_B|I_D1|B 0 I1_|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_SPL_B|I_D2|B I1_|_SPL_B|D2 I1_|_SPL_B|I_D2|MID  2e-12
II1_|_SPL_B|I_D2|B 0 I1_|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI1_|_SPL_B|I_Q1|B I1_|_SPL_B|QA1 I1_|_SPL_B|I_Q1|MID  2e-12
II1_|_SPL_B|I_Q1|B 0 I1_|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_SPL_B|I_Q2|B I1_|_SPL_B|QB1 I1_|_SPL_B|I_Q2|MID  2e-12
II1_|_SPL_B|I_Q2|B 0 I1_|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI1_|_SPL_B|1|1 I1_|_SPL_B|D1 I1_|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_B|1|P I1_|_SPL_B|1|MID_SERIES 0  2e-13
RI1_|_SPL_B|1|B I1_|_SPL_B|D1 I1_|_SPL_B|1|MID_SHUNT  2.7439617672
LI1_|_SPL_B|1|RB I1_|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI1_|_SPL_B|2|1 I1_|_SPL_B|D2 I1_|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_B|2|P I1_|_SPL_B|2|MID_SERIES 0  2e-13
RI1_|_SPL_B|2|B I1_|_SPL_B|D2 I1_|_SPL_B|2|MID_SHUNT  2.7439617672
LI1_|_SPL_B|2|RB I1_|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI1_|_SPL_B|A|1 I1_|_SPL_B|QA1 I1_|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_B|A|P I1_|_SPL_B|A|MID_SERIES 0  2e-13
RI1_|_SPL_B|A|B I1_|_SPL_B|QA1 I1_|_SPL_B|A|MID_SHUNT  2.7439617672
LI1_|_SPL_B|A|RB I1_|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI1_|_SPL_B|B|1 I1_|_SPL_B|QB1 I1_|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI1_|_SPL_B|B|P I1_|_SPL_B|B|MID_SERIES 0  2e-13
RI1_|_SPL_B|B|B I1_|_SPL_B|QB1 I1_|_SPL_B|B|MID_SHUNT  2.7439617672
LI1_|_SPL_B|B|RB I1_|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI1_|_DFF_A|I_1|B I1_|_DFF_A|A1 I1_|_DFF_A|I_1|MID  2e-12
II1_|_DFF_A|I_1|B 0 I1_|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_DFF_A|I_3|B I1_|_DFF_A|A3 I1_|_DFF_A|I_3|MID  2e-12
II1_|_DFF_A|I_3|B 0 I1_|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1_|_DFF_A|I_T|B I1_|_DFF_A|T1 I1_|_DFF_A|I_T|MID  2e-12
II1_|_DFF_A|I_T|B 0 I1_|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1_|_DFF_A|I_6|B I1_|_DFF_A|Q1 I1_|_DFF_A|I_6|MID  2e-12
II1_|_DFF_A|I_6|B 0 I1_|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1_|_DFF_A|1|1 I1_|_DFF_A|A1 I1_|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_A|1|P I1_|_DFF_A|1|MID_SERIES 0  2e-13
RI1_|_DFF_A|1|B I1_|_DFF_A|A1 I1_|_DFF_A|1|MID_SHUNT  2.7439617672
LI1_|_DFF_A|1|RB I1_|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_A|23|1 I1_|_DFF_A|A2 I1_|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI1_|_DFF_A|23|B I1_|_DFF_A|A2 I1_|_DFF_A|23|MID_SHUNT  3.84154647408
LI1_|_DFF_A|23|RB I1_|_DFF_A|23|MID_SHUNT I1_|_DFF_A|A3  2.1704737578552e-12
BI1_|_DFF_A|3|1 I1_|_DFF_A|A3 I1_|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_A|3|P I1_|_DFF_A|3|MID_SERIES 0  2e-13
RI1_|_DFF_A|3|B I1_|_DFF_A|A3 I1_|_DFF_A|3|MID_SHUNT  2.7439617672
LI1_|_DFF_A|3|RB I1_|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_A|4|1 I1_|_DFF_A|A4 I1_|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_A|4|P I1_|_DFF_A|4|MID_SERIES 0  2e-13
RI1_|_DFF_A|4|B I1_|_DFF_A|A4 I1_|_DFF_A|4|MID_SHUNT  2.7439617672
LI1_|_DFF_A|4|RB I1_|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_A|T|1 I1_|_DFF_A|T1 I1_|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_A|T|P I1_|_DFF_A|T|MID_SERIES 0  2e-13
RI1_|_DFF_A|T|B I1_|_DFF_A|T1 I1_|_DFF_A|T|MID_SHUNT  2.7439617672
LI1_|_DFF_A|T|RB I1_|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_A|45|1 I1_|_DFF_A|T2 I1_|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI1_|_DFF_A|45|B I1_|_DFF_A|T2 I1_|_DFF_A|45|MID_SHUNT  3.84154647408
LI1_|_DFF_A|45|RB I1_|_DFF_A|45|MID_SHUNT I1_|_DFF_A|A4  2.1704737578552e-12
BI1_|_DFF_A|6|1 I1_|_DFF_A|Q1 I1_|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_A|6|P I1_|_DFF_A|6|MID_SERIES 0  2e-13
RI1_|_DFF_A|6|B I1_|_DFF_A|Q1 I1_|_DFF_A|6|MID_SHUNT  2.7439617672
LI1_|_DFF_A|6|RB I1_|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI1_|_DFF_B|I_1|B I1_|_DFF_B|A1 I1_|_DFF_B|I_1|MID  2e-12
II1_|_DFF_B|I_1|B 0 I1_|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_DFF_B|I_3|B I1_|_DFF_B|A3 I1_|_DFF_B|I_3|MID  2e-12
II1_|_DFF_B|I_3|B 0 I1_|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1_|_DFF_B|I_T|B I1_|_DFF_B|T1 I1_|_DFF_B|I_T|MID  2e-12
II1_|_DFF_B|I_T|B 0 I1_|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1_|_DFF_B|I_6|B I1_|_DFF_B|Q1 I1_|_DFF_B|I_6|MID  2e-12
II1_|_DFF_B|I_6|B 0 I1_|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1_|_DFF_B|1|1 I1_|_DFF_B|A1 I1_|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_B|1|P I1_|_DFF_B|1|MID_SERIES 0  2e-13
RI1_|_DFF_B|1|B I1_|_DFF_B|A1 I1_|_DFF_B|1|MID_SHUNT  2.7439617672
LI1_|_DFF_B|1|RB I1_|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_B|23|1 I1_|_DFF_B|A2 I1_|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI1_|_DFF_B|23|B I1_|_DFF_B|A2 I1_|_DFF_B|23|MID_SHUNT  3.84154647408
LI1_|_DFF_B|23|RB I1_|_DFF_B|23|MID_SHUNT I1_|_DFF_B|A3  2.1704737578552e-12
BI1_|_DFF_B|3|1 I1_|_DFF_B|A3 I1_|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_B|3|P I1_|_DFF_B|3|MID_SERIES 0  2e-13
RI1_|_DFF_B|3|B I1_|_DFF_B|A3 I1_|_DFF_B|3|MID_SHUNT  2.7439617672
LI1_|_DFF_B|3|RB I1_|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_B|4|1 I1_|_DFF_B|A4 I1_|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_B|4|P I1_|_DFF_B|4|MID_SERIES 0  2e-13
RI1_|_DFF_B|4|B I1_|_DFF_B|A4 I1_|_DFF_B|4|MID_SHUNT  2.7439617672
LI1_|_DFF_B|4|RB I1_|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_B|T|1 I1_|_DFF_B|T1 I1_|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_B|T|P I1_|_DFF_B|T|MID_SERIES 0  2e-13
RI1_|_DFF_B|T|B I1_|_DFF_B|T1 I1_|_DFF_B|T|MID_SHUNT  2.7439617672
LI1_|_DFF_B|T|RB I1_|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI1_|_DFF_B|45|1 I1_|_DFF_B|T2 I1_|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI1_|_DFF_B|45|B I1_|_DFF_B|T2 I1_|_DFF_B|45|MID_SHUNT  3.84154647408
LI1_|_DFF_B|45|RB I1_|_DFF_B|45|MID_SHUNT I1_|_DFF_B|A4  2.1704737578552e-12
BI1_|_DFF_B|6|1 I1_|_DFF_B|Q1 I1_|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI1_|_DFF_B|6|P I1_|_DFF_B|6|MID_SERIES 0  2e-13
RI1_|_DFF_B|6|B I1_|_DFF_B|Q1 I1_|_DFF_B|6|MID_SHUNT  2.7439617672
LI1_|_DFF_B|6|RB I1_|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI1_|_XOR|I_A1|B I1_|_XOR|A1 I1_|_XOR|I_A1|MID  2e-12
II1_|_XOR|I_A1|B 0 I1_|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_XOR|I_A3|B I1_|_XOR|A3 I1_|_XOR|I_A3|MID  2e-12
II1_|_XOR|I_A3|B 0 I1_|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI1_|_XOR|I_B1|B I1_|_XOR|B1 I1_|_XOR|I_B1|MID  2e-12
II1_|_XOR|I_B1|B 0 I1_|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_XOR|I_B3|B I1_|_XOR|B3 I1_|_XOR|I_B3|MID  2e-12
II1_|_XOR|I_B3|B 0 I1_|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI1_|_XOR|I_Q1|B I1_|_XOR|Q1 I1_|_XOR|I_Q1|MID  2e-12
II1_|_XOR|I_Q1|B 0 I1_|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1_|_XOR|A1|1 I1_|_XOR|A1 I1_|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|A1|P I1_|_XOR|A1|MID_SERIES 0  5e-13
RI1_|_XOR|A1|B I1_|_XOR|A1 I1_|_XOR|A1|MID_SHUNT  2.7439617672
LI1_|_XOR|A1|RB I1_|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI1_|_XOR|A2|1 I1_|_XOR|A2 I1_|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|A2|P I1_|_XOR|A2|MID_SERIES 0  5e-13
RI1_|_XOR|A2|B I1_|_XOR|A2 I1_|_XOR|A2|MID_SHUNT  2.7439617672
LI1_|_XOR|A2|RB I1_|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI1_|_XOR|A3|1 I1_|_XOR|A2 I1_|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|A3|P I1_|_XOR|A3|MID_SERIES I1_|_XOR|A3  1.2e-12
RI1_|_XOR|A3|B I1_|_XOR|A2 I1_|_XOR|A3|MID_SHUNT  2.7439617672
LI1_|_XOR|A3|RB I1_|_XOR|A3|MID_SHUNT I1_|_XOR|A3  2.050338398468e-12
BI1_|_XOR|B1|1 I1_|_XOR|B1 I1_|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|B1|P I1_|_XOR|B1|MID_SERIES 0  5e-13
RI1_|_XOR|B1|B I1_|_XOR|B1 I1_|_XOR|B1|MID_SHUNT  2.7439617672
LI1_|_XOR|B1|RB I1_|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI1_|_XOR|B2|1 I1_|_XOR|B2 I1_|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|B2|P I1_|_XOR|B2|MID_SERIES 0  5e-13
RI1_|_XOR|B2|B I1_|_XOR|B2 I1_|_XOR|B2|MID_SHUNT  2.7439617672
LI1_|_XOR|B2|RB I1_|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI1_|_XOR|B3|1 I1_|_XOR|B2 I1_|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|B3|P I1_|_XOR|B3|MID_SERIES I1_|_XOR|B3  1.2e-12
RI1_|_XOR|B3|B I1_|_XOR|B2 I1_|_XOR|B3|MID_SHUNT  2.7439617672
LI1_|_XOR|B3|RB I1_|_XOR|B3|MID_SHUNT I1_|_XOR|B3  2.050338398468e-12
BI1_|_XOR|T1|1 I1_|_XOR|T1 I1_|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|T1|P I1_|_XOR|T1|MID_SERIES 0  5e-13
RI1_|_XOR|T1|B I1_|_XOR|T1 I1_|_XOR|T1|MID_SHUNT  2.7439617672
LI1_|_XOR|T1|RB I1_|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI1_|_XOR|T2|1 I1_|_XOR|T2 I1_|_XOR|ABTQ JJMIT AREA=2.0
RI1_|_XOR|T2|B I1_|_XOR|T2 I1_|_XOR|T2|MID_SHUNT  3.429952209
LI1_|_XOR|T2|RB I1_|_XOR|T2|MID_SHUNT I1_|_XOR|ABTQ  2.437922998085e-12
BI1_|_XOR|AB|1 I1_|_XOR|AB I1_|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI1_|_XOR|AB|P I1_|_XOR|AB|MID_SERIES I1_|_XOR|ABTQ  1.2e-12
RI1_|_XOR|AB|B I1_|_XOR|AB I1_|_XOR|AB|MID_SHUNT  3.429952209
LI1_|_XOR|AB|RB I1_|_XOR|AB|MID_SHUNT I1_|_XOR|ABTQ  2.437922998085e-12
BI1_|_XOR|ABTQ|1 I1_|_XOR|ABTQ I1_|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|ABTQ|P I1_|_XOR|ABTQ|MID_SERIES 0  5e-13
RI1_|_XOR|ABTQ|B I1_|_XOR|ABTQ I1_|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI1_|_XOR|ABTQ|RB I1_|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI1_|_XOR|Q1|1 I1_|_XOR|Q1 I1_|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI1_|_XOR|Q1|P I1_|_XOR|Q1|MID_SERIES 0  5e-13
RI1_|_XOR|Q1|B I1_|_XOR|Q1 I1_|_XOR|Q1|MID_SHUNT  2.7439617672
LI1_|_XOR|Q1|RB I1_|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI1_|_AND|I_A1|B I1_|_AND|A1 I1_|_AND|I_A1|MID  2e-12
II1_|_AND|I_A1|B 0 I1_|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_AND|I_B1|B I1_|_AND|B1 I1_|_AND|I_B1|MID  2e-12
II1_|_AND|I_B1|B 0 I1_|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1_|_AND|I_Q3|B I1_|_AND|Q3 I1_|_AND|I_Q3|MID  2e-12
II1_|_AND|I_Q3|B 0 I1_|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1_|_AND|I_Q2|B I1_|_AND|Q2 I1_|_AND|I_Q2|MID  2e-12
II1_|_AND|I_Q2|B 0 I1_|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1_|_AND|I_Q1|B I1_|_AND|Q1 I1_|_AND|I_Q1|MID  2e-12
II1_|_AND|I_Q1|B 0 I1_|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1_|_AND|A1|1 I1_|_AND|A1 I1_|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1_|_AND|A1|P I1_|_AND|A1|MID_SERIES 0  2e-13
RI1_|_AND|A1|B I1_|_AND|A1 I1_|_AND|A1|MID_SHUNT  2.7439617672
LI1_|_AND|A1|RB I1_|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1_|_AND|A2|1 I1_|_AND|A2 I1_|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1_|_AND|A2|P I1_|_AND|A2|MID_SERIES 0  2e-13
RI1_|_AND|A2|B I1_|_AND|A2 I1_|_AND|A2|MID_SHUNT  2.7439617672
LI1_|_AND|A2|RB I1_|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1_|_AND|A12|1 I1_|_AND|A2 I1_|_AND|A3 JJMIT AREA=1.7857142857142858
RI1_|_AND|A12|B I1_|_AND|A2 I1_|_AND|A12|MID_SHUNT  3.84154647408
LI1_|_AND|A12|RB I1_|_AND|A12|MID_SHUNT I1_|_AND|A3  2.1704737578552e-12
BI1_|_AND|B1|1 I1_|_AND|B1 I1_|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1_|_AND|B1|P I1_|_AND|B1|MID_SERIES 0  2e-13
RI1_|_AND|B1|B I1_|_AND|B1 I1_|_AND|B1|MID_SHUNT  2.7439617672
LI1_|_AND|B1|RB I1_|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1_|_AND|B2|1 I1_|_AND|B2 I1_|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1_|_AND|B2|P I1_|_AND|B2|MID_SERIES 0  2e-13
RI1_|_AND|B2|B I1_|_AND|B2 I1_|_AND|B2|MID_SHUNT  2.7439617672
LI1_|_AND|B2|RB I1_|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1_|_AND|B12|1 I1_|_AND|B2 I1_|_AND|B3 JJMIT AREA=1.7857142857142858
RI1_|_AND|B12|B I1_|_AND|B2 I1_|_AND|B12|MID_SHUNT  3.84154647408
LI1_|_AND|B12|RB I1_|_AND|B12|MID_SHUNT I1_|_AND|B3  2.1704737578552e-12
BI1_|_AND|Q2|1 I1_|_AND|Q2 I1_|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1_|_AND|Q2|P I1_|_AND|Q2|MID_SERIES 0  2e-13
RI1_|_AND|Q2|B I1_|_AND|Q2 I1_|_AND|Q2|MID_SHUNT  2.7439617672
LI1_|_AND|Q2|RB I1_|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1_|_AND|Q1|1 I1_|_AND|Q1 I1_|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1_|_AND|Q1|P I1_|_AND|Q1|MID_SERIES 0  2e-13
RI1_|_AND|Q1|B I1_|_AND|Q1 I1_|_AND|Q1|MID_SHUNT  2.7439617672
LI1_|_AND|Q1|RB I1_|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2_|_SPL_A|I_D1|B I2_|_SPL_A|D1 I2_|_SPL_A|I_D1|MID  2e-12
II2_|_SPL_A|I_D1|B 0 I2_|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_SPL_A|I_D2|B I2_|_SPL_A|D2 I2_|_SPL_A|I_D2|MID  2e-12
II2_|_SPL_A|I_D2|B 0 I2_|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI2_|_SPL_A|I_Q1|B I2_|_SPL_A|QA1 I2_|_SPL_A|I_Q1|MID  2e-12
II2_|_SPL_A|I_Q1|B 0 I2_|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_SPL_A|I_Q2|B I2_|_SPL_A|QB1 I2_|_SPL_A|I_Q2|MID  2e-12
II2_|_SPL_A|I_Q2|B 0 I2_|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI2_|_SPL_A|1|1 I2_|_SPL_A|D1 I2_|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_A|1|P I2_|_SPL_A|1|MID_SERIES 0  2e-13
RI2_|_SPL_A|1|B I2_|_SPL_A|D1 I2_|_SPL_A|1|MID_SHUNT  2.7439617672
LI2_|_SPL_A|1|RB I2_|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI2_|_SPL_A|2|1 I2_|_SPL_A|D2 I2_|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_A|2|P I2_|_SPL_A|2|MID_SERIES 0  2e-13
RI2_|_SPL_A|2|B I2_|_SPL_A|D2 I2_|_SPL_A|2|MID_SHUNT  2.7439617672
LI2_|_SPL_A|2|RB I2_|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI2_|_SPL_A|A|1 I2_|_SPL_A|QA1 I2_|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_A|A|P I2_|_SPL_A|A|MID_SERIES 0  2e-13
RI2_|_SPL_A|A|B I2_|_SPL_A|QA1 I2_|_SPL_A|A|MID_SHUNT  2.7439617672
LI2_|_SPL_A|A|RB I2_|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI2_|_SPL_A|B|1 I2_|_SPL_A|QB1 I2_|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_A|B|P I2_|_SPL_A|B|MID_SERIES 0  2e-13
RI2_|_SPL_A|B|B I2_|_SPL_A|QB1 I2_|_SPL_A|B|MID_SHUNT  2.7439617672
LI2_|_SPL_A|B|RB I2_|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI2_|_SPL_B|I_D1|B I2_|_SPL_B|D1 I2_|_SPL_B|I_D1|MID  2e-12
II2_|_SPL_B|I_D1|B 0 I2_|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_SPL_B|I_D2|B I2_|_SPL_B|D2 I2_|_SPL_B|I_D2|MID  2e-12
II2_|_SPL_B|I_D2|B 0 I2_|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI2_|_SPL_B|I_Q1|B I2_|_SPL_B|QA1 I2_|_SPL_B|I_Q1|MID  2e-12
II2_|_SPL_B|I_Q1|B 0 I2_|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_SPL_B|I_Q2|B I2_|_SPL_B|QB1 I2_|_SPL_B|I_Q2|MID  2e-12
II2_|_SPL_B|I_Q2|B 0 I2_|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI2_|_SPL_B|1|1 I2_|_SPL_B|D1 I2_|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_B|1|P I2_|_SPL_B|1|MID_SERIES 0  2e-13
RI2_|_SPL_B|1|B I2_|_SPL_B|D1 I2_|_SPL_B|1|MID_SHUNT  2.7439617672
LI2_|_SPL_B|1|RB I2_|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI2_|_SPL_B|2|1 I2_|_SPL_B|D2 I2_|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_B|2|P I2_|_SPL_B|2|MID_SERIES 0  2e-13
RI2_|_SPL_B|2|B I2_|_SPL_B|D2 I2_|_SPL_B|2|MID_SHUNT  2.7439617672
LI2_|_SPL_B|2|RB I2_|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI2_|_SPL_B|A|1 I2_|_SPL_B|QA1 I2_|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_B|A|P I2_|_SPL_B|A|MID_SERIES 0  2e-13
RI2_|_SPL_B|A|B I2_|_SPL_B|QA1 I2_|_SPL_B|A|MID_SHUNT  2.7439617672
LI2_|_SPL_B|A|RB I2_|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI2_|_SPL_B|B|1 I2_|_SPL_B|QB1 I2_|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI2_|_SPL_B|B|P I2_|_SPL_B|B|MID_SERIES 0  2e-13
RI2_|_SPL_B|B|B I2_|_SPL_B|QB1 I2_|_SPL_B|B|MID_SHUNT  2.7439617672
LI2_|_SPL_B|B|RB I2_|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI2_|_DFF_A|I_1|B I2_|_DFF_A|A1 I2_|_DFF_A|I_1|MID  2e-12
II2_|_DFF_A|I_1|B 0 I2_|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_DFF_A|I_3|B I2_|_DFF_A|A3 I2_|_DFF_A|I_3|MID  2e-12
II2_|_DFF_A|I_3|B 0 I2_|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2_|_DFF_A|I_T|B I2_|_DFF_A|T1 I2_|_DFF_A|I_T|MID  2e-12
II2_|_DFF_A|I_T|B 0 I2_|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2_|_DFF_A|I_6|B I2_|_DFF_A|Q1 I2_|_DFF_A|I_6|MID  2e-12
II2_|_DFF_A|I_6|B 0 I2_|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2_|_DFF_A|1|1 I2_|_DFF_A|A1 I2_|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_A|1|P I2_|_DFF_A|1|MID_SERIES 0  2e-13
RI2_|_DFF_A|1|B I2_|_DFF_A|A1 I2_|_DFF_A|1|MID_SHUNT  2.7439617672
LI2_|_DFF_A|1|RB I2_|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_A|23|1 I2_|_DFF_A|A2 I2_|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI2_|_DFF_A|23|B I2_|_DFF_A|A2 I2_|_DFF_A|23|MID_SHUNT  3.84154647408
LI2_|_DFF_A|23|RB I2_|_DFF_A|23|MID_SHUNT I2_|_DFF_A|A3  2.1704737578552e-12
BI2_|_DFF_A|3|1 I2_|_DFF_A|A3 I2_|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_A|3|P I2_|_DFF_A|3|MID_SERIES 0  2e-13
RI2_|_DFF_A|3|B I2_|_DFF_A|A3 I2_|_DFF_A|3|MID_SHUNT  2.7439617672
LI2_|_DFF_A|3|RB I2_|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_A|4|1 I2_|_DFF_A|A4 I2_|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_A|4|P I2_|_DFF_A|4|MID_SERIES 0  2e-13
RI2_|_DFF_A|4|B I2_|_DFF_A|A4 I2_|_DFF_A|4|MID_SHUNT  2.7439617672
LI2_|_DFF_A|4|RB I2_|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_A|T|1 I2_|_DFF_A|T1 I2_|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_A|T|P I2_|_DFF_A|T|MID_SERIES 0  2e-13
RI2_|_DFF_A|T|B I2_|_DFF_A|T1 I2_|_DFF_A|T|MID_SHUNT  2.7439617672
LI2_|_DFF_A|T|RB I2_|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_A|45|1 I2_|_DFF_A|T2 I2_|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI2_|_DFF_A|45|B I2_|_DFF_A|T2 I2_|_DFF_A|45|MID_SHUNT  3.84154647408
LI2_|_DFF_A|45|RB I2_|_DFF_A|45|MID_SHUNT I2_|_DFF_A|A4  2.1704737578552e-12
BI2_|_DFF_A|6|1 I2_|_DFF_A|Q1 I2_|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_A|6|P I2_|_DFF_A|6|MID_SERIES 0  2e-13
RI2_|_DFF_A|6|B I2_|_DFF_A|Q1 I2_|_DFF_A|6|MID_SHUNT  2.7439617672
LI2_|_DFF_A|6|RB I2_|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI2_|_DFF_B|I_1|B I2_|_DFF_B|A1 I2_|_DFF_B|I_1|MID  2e-12
II2_|_DFF_B|I_1|B 0 I2_|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_DFF_B|I_3|B I2_|_DFF_B|A3 I2_|_DFF_B|I_3|MID  2e-12
II2_|_DFF_B|I_3|B 0 I2_|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2_|_DFF_B|I_T|B I2_|_DFF_B|T1 I2_|_DFF_B|I_T|MID  2e-12
II2_|_DFF_B|I_T|B 0 I2_|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2_|_DFF_B|I_6|B I2_|_DFF_B|Q1 I2_|_DFF_B|I_6|MID  2e-12
II2_|_DFF_B|I_6|B 0 I2_|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2_|_DFF_B|1|1 I2_|_DFF_B|A1 I2_|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_B|1|P I2_|_DFF_B|1|MID_SERIES 0  2e-13
RI2_|_DFF_B|1|B I2_|_DFF_B|A1 I2_|_DFF_B|1|MID_SHUNT  2.7439617672
LI2_|_DFF_B|1|RB I2_|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_B|23|1 I2_|_DFF_B|A2 I2_|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI2_|_DFF_B|23|B I2_|_DFF_B|A2 I2_|_DFF_B|23|MID_SHUNT  3.84154647408
LI2_|_DFF_B|23|RB I2_|_DFF_B|23|MID_SHUNT I2_|_DFF_B|A3  2.1704737578552e-12
BI2_|_DFF_B|3|1 I2_|_DFF_B|A3 I2_|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_B|3|P I2_|_DFF_B|3|MID_SERIES 0  2e-13
RI2_|_DFF_B|3|B I2_|_DFF_B|A3 I2_|_DFF_B|3|MID_SHUNT  2.7439617672
LI2_|_DFF_B|3|RB I2_|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_B|4|1 I2_|_DFF_B|A4 I2_|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_B|4|P I2_|_DFF_B|4|MID_SERIES 0  2e-13
RI2_|_DFF_B|4|B I2_|_DFF_B|A4 I2_|_DFF_B|4|MID_SHUNT  2.7439617672
LI2_|_DFF_B|4|RB I2_|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_B|T|1 I2_|_DFF_B|T1 I2_|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_B|T|P I2_|_DFF_B|T|MID_SERIES 0  2e-13
RI2_|_DFF_B|T|B I2_|_DFF_B|T1 I2_|_DFF_B|T|MID_SHUNT  2.7439617672
LI2_|_DFF_B|T|RB I2_|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI2_|_DFF_B|45|1 I2_|_DFF_B|T2 I2_|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI2_|_DFF_B|45|B I2_|_DFF_B|T2 I2_|_DFF_B|45|MID_SHUNT  3.84154647408
LI2_|_DFF_B|45|RB I2_|_DFF_B|45|MID_SHUNT I2_|_DFF_B|A4  2.1704737578552e-12
BI2_|_DFF_B|6|1 I2_|_DFF_B|Q1 I2_|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI2_|_DFF_B|6|P I2_|_DFF_B|6|MID_SERIES 0  2e-13
RI2_|_DFF_B|6|B I2_|_DFF_B|Q1 I2_|_DFF_B|6|MID_SHUNT  2.7439617672
LI2_|_DFF_B|6|RB I2_|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI2_|_XOR|I_A1|B I2_|_XOR|A1 I2_|_XOR|I_A1|MID  2e-12
II2_|_XOR|I_A1|B 0 I2_|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_XOR|I_A3|B I2_|_XOR|A3 I2_|_XOR|I_A3|MID  2e-12
II2_|_XOR|I_A3|B 0 I2_|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI2_|_XOR|I_B1|B I2_|_XOR|B1 I2_|_XOR|I_B1|MID  2e-12
II2_|_XOR|I_B1|B 0 I2_|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_XOR|I_B3|B I2_|_XOR|B3 I2_|_XOR|I_B3|MID  2e-12
II2_|_XOR|I_B3|B 0 I2_|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI2_|_XOR|I_Q1|B I2_|_XOR|Q1 I2_|_XOR|I_Q1|MID  2e-12
II2_|_XOR|I_Q1|B 0 I2_|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2_|_XOR|A1|1 I2_|_XOR|A1 I2_|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|A1|P I2_|_XOR|A1|MID_SERIES 0  5e-13
RI2_|_XOR|A1|B I2_|_XOR|A1 I2_|_XOR|A1|MID_SHUNT  2.7439617672
LI2_|_XOR|A1|RB I2_|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI2_|_XOR|A2|1 I2_|_XOR|A2 I2_|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|A2|P I2_|_XOR|A2|MID_SERIES 0  5e-13
RI2_|_XOR|A2|B I2_|_XOR|A2 I2_|_XOR|A2|MID_SHUNT  2.7439617672
LI2_|_XOR|A2|RB I2_|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI2_|_XOR|A3|1 I2_|_XOR|A2 I2_|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|A3|P I2_|_XOR|A3|MID_SERIES I2_|_XOR|A3  1.2e-12
RI2_|_XOR|A3|B I2_|_XOR|A2 I2_|_XOR|A3|MID_SHUNT  2.7439617672
LI2_|_XOR|A3|RB I2_|_XOR|A3|MID_SHUNT I2_|_XOR|A3  2.050338398468e-12
BI2_|_XOR|B1|1 I2_|_XOR|B1 I2_|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|B1|P I2_|_XOR|B1|MID_SERIES 0  5e-13
RI2_|_XOR|B1|B I2_|_XOR|B1 I2_|_XOR|B1|MID_SHUNT  2.7439617672
LI2_|_XOR|B1|RB I2_|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI2_|_XOR|B2|1 I2_|_XOR|B2 I2_|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|B2|P I2_|_XOR|B2|MID_SERIES 0  5e-13
RI2_|_XOR|B2|B I2_|_XOR|B2 I2_|_XOR|B2|MID_SHUNT  2.7439617672
LI2_|_XOR|B2|RB I2_|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI2_|_XOR|B3|1 I2_|_XOR|B2 I2_|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|B3|P I2_|_XOR|B3|MID_SERIES I2_|_XOR|B3  1.2e-12
RI2_|_XOR|B3|B I2_|_XOR|B2 I2_|_XOR|B3|MID_SHUNT  2.7439617672
LI2_|_XOR|B3|RB I2_|_XOR|B3|MID_SHUNT I2_|_XOR|B3  2.050338398468e-12
BI2_|_XOR|T1|1 I2_|_XOR|T1 I2_|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|T1|P I2_|_XOR|T1|MID_SERIES 0  5e-13
RI2_|_XOR|T1|B I2_|_XOR|T1 I2_|_XOR|T1|MID_SHUNT  2.7439617672
LI2_|_XOR|T1|RB I2_|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI2_|_XOR|T2|1 I2_|_XOR|T2 I2_|_XOR|ABTQ JJMIT AREA=2.0
RI2_|_XOR|T2|B I2_|_XOR|T2 I2_|_XOR|T2|MID_SHUNT  3.429952209
LI2_|_XOR|T2|RB I2_|_XOR|T2|MID_SHUNT I2_|_XOR|ABTQ  2.437922998085e-12
BI2_|_XOR|AB|1 I2_|_XOR|AB I2_|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI2_|_XOR|AB|P I2_|_XOR|AB|MID_SERIES I2_|_XOR|ABTQ  1.2e-12
RI2_|_XOR|AB|B I2_|_XOR|AB I2_|_XOR|AB|MID_SHUNT  3.429952209
LI2_|_XOR|AB|RB I2_|_XOR|AB|MID_SHUNT I2_|_XOR|ABTQ  2.437922998085e-12
BI2_|_XOR|ABTQ|1 I2_|_XOR|ABTQ I2_|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|ABTQ|P I2_|_XOR|ABTQ|MID_SERIES 0  5e-13
RI2_|_XOR|ABTQ|B I2_|_XOR|ABTQ I2_|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI2_|_XOR|ABTQ|RB I2_|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI2_|_XOR|Q1|1 I2_|_XOR|Q1 I2_|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI2_|_XOR|Q1|P I2_|_XOR|Q1|MID_SERIES 0  5e-13
RI2_|_XOR|Q1|B I2_|_XOR|Q1 I2_|_XOR|Q1|MID_SHUNT  2.7439617672
LI2_|_XOR|Q1|RB I2_|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI2_|_AND|I_A1|B I2_|_AND|A1 I2_|_AND|I_A1|MID  2e-12
II2_|_AND|I_A1|B 0 I2_|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_AND|I_B1|B I2_|_AND|B1 I2_|_AND|I_B1|MID  2e-12
II2_|_AND|I_B1|B 0 I2_|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2_|_AND|I_Q3|B I2_|_AND|Q3 I2_|_AND|I_Q3|MID  2e-12
II2_|_AND|I_Q3|B 0 I2_|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2_|_AND|I_Q2|B I2_|_AND|Q2 I2_|_AND|I_Q2|MID  2e-12
II2_|_AND|I_Q2|B 0 I2_|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2_|_AND|I_Q1|B I2_|_AND|Q1 I2_|_AND|I_Q1|MID  2e-12
II2_|_AND|I_Q1|B 0 I2_|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2_|_AND|A1|1 I2_|_AND|A1 I2_|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2_|_AND|A1|P I2_|_AND|A1|MID_SERIES 0  2e-13
RI2_|_AND|A1|B I2_|_AND|A1 I2_|_AND|A1|MID_SHUNT  2.7439617672
LI2_|_AND|A1|RB I2_|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2_|_AND|A2|1 I2_|_AND|A2 I2_|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2_|_AND|A2|P I2_|_AND|A2|MID_SERIES 0  2e-13
RI2_|_AND|A2|B I2_|_AND|A2 I2_|_AND|A2|MID_SHUNT  2.7439617672
LI2_|_AND|A2|RB I2_|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2_|_AND|A12|1 I2_|_AND|A2 I2_|_AND|A3 JJMIT AREA=1.7857142857142858
RI2_|_AND|A12|B I2_|_AND|A2 I2_|_AND|A12|MID_SHUNT  3.84154647408
LI2_|_AND|A12|RB I2_|_AND|A12|MID_SHUNT I2_|_AND|A3  2.1704737578552e-12
BI2_|_AND|B1|1 I2_|_AND|B1 I2_|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2_|_AND|B1|P I2_|_AND|B1|MID_SERIES 0  2e-13
RI2_|_AND|B1|B I2_|_AND|B1 I2_|_AND|B1|MID_SHUNT  2.7439617672
LI2_|_AND|B1|RB I2_|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2_|_AND|B2|1 I2_|_AND|B2 I2_|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2_|_AND|B2|P I2_|_AND|B2|MID_SERIES 0  2e-13
RI2_|_AND|B2|B I2_|_AND|B2 I2_|_AND|B2|MID_SHUNT  2.7439617672
LI2_|_AND|B2|RB I2_|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2_|_AND|B12|1 I2_|_AND|B2 I2_|_AND|B3 JJMIT AREA=1.7857142857142858
RI2_|_AND|B12|B I2_|_AND|B2 I2_|_AND|B12|MID_SHUNT  3.84154647408
LI2_|_AND|B12|RB I2_|_AND|B12|MID_SHUNT I2_|_AND|B3  2.1704737578552e-12
BI2_|_AND|Q2|1 I2_|_AND|Q2 I2_|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2_|_AND|Q2|P I2_|_AND|Q2|MID_SERIES 0  2e-13
RI2_|_AND|Q2|B I2_|_AND|Q2 I2_|_AND|Q2|MID_SHUNT  2.7439617672
LI2_|_AND|Q2|RB I2_|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2_|_AND|Q1|1 I2_|_AND|Q1 I2_|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2_|_AND|Q1|P I2_|_AND|Q1|MID_SERIES 0  2e-13
RI2_|_AND|Q1|B I2_|_AND|Q1 I2_|_AND|Q1|MID_SHUNT  2.7439617672
LI2_|_AND|Q1|RB I2_|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3_|_SPL_A|I_D1|B I3_|_SPL_A|D1 I3_|_SPL_A|I_D1|MID  2e-12
II3_|_SPL_A|I_D1|B 0 I3_|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_SPL_A|I_D2|B I3_|_SPL_A|D2 I3_|_SPL_A|I_D2|MID  2e-12
II3_|_SPL_A|I_D2|B 0 I3_|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI3_|_SPL_A|I_Q1|B I3_|_SPL_A|QA1 I3_|_SPL_A|I_Q1|MID  2e-12
II3_|_SPL_A|I_Q1|B 0 I3_|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_SPL_A|I_Q2|B I3_|_SPL_A|QB1 I3_|_SPL_A|I_Q2|MID  2e-12
II3_|_SPL_A|I_Q2|B 0 I3_|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI3_|_SPL_A|1|1 I3_|_SPL_A|D1 I3_|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_A|1|P I3_|_SPL_A|1|MID_SERIES 0  2e-13
RI3_|_SPL_A|1|B I3_|_SPL_A|D1 I3_|_SPL_A|1|MID_SHUNT  2.7439617672
LI3_|_SPL_A|1|RB I3_|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI3_|_SPL_A|2|1 I3_|_SPL_A|D2 I3_|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_A|2|P I3_|_SPL_A|2|MID_SERIES 0  2e-13
RI3_|_SPL_A|2|B I3_|_SPL_A|D2 I3_|_SPL_A|2|MID_SHUNT  2.7439617672
LI3_|_SPL_A|2|RB I3_|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI3_|_SPL_A|A|1 I3_|_SPL_A|QA1 I3_|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_A|A|P I3_|_SPL_A|A|MID_SERIES 0  2e-13
RI3_|_SPL_A|A|B I3_|_SPL_A|QA1 I3_|_SPL_A|A|MID_SHUNT  2.7439617672
LI3_|_SPL_A|A|RB I3_|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI3_|_SPL_A|B|1 I3_|_SPL_A|QB1 I3_|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_A|B|P I3_|_SPL_A|B|MID_SERIES 0  2e-13
RI3_|_SPL_A|B|B I3_|_SPL_A|QB1 I3_|_SPL_A|B|MID_SHUNT  2.7439617672
LI3_|_SPL_A|B|RB I3_|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI3_|_SPL_B|I_D1|B I3_|_SPL_B|D1 I3_|_SPL_B|I_D1|MID  2e-12
II3_|_SPL_B|I_D1|B 0 I3_|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_SPL_B|I_D2|B I3_|_SPL_B|D2 I3_|_SPL_B|I_D2|MID  2e-12
II3_|_SPL_B|I_D2|B 0 I3_|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.000245)
LI3_|_SPL_B|I_Q1|B I3_|_SPL_B|QA1 I3_|_SPL_B|I_Q1|MID  2e-12
II3_|_SPL_B|I_Q1|B 0 I3_|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_SPL_B|I_Q2|B I3_|_SPL_B|QB1 I3_|_SPL_B|I_Q2|MID  2e-12
II3_|_SPL_B|I_Q2|B 0 I3_|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BI3_|_SPL_B|1|1 I3_|_SPL_B|D1 I3_|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_B|1|P I3_|_SPL_B|1|MID_SERIES 0  2e-13
RI3_|_SPL_B|1|B I3_|_SPL_B|D1 I3_|_SPL_B|1|MID_SHUNT  2.7439617672
LI3_|_SPL_B|1|RB I3_|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI3_|_SPL_B|2|1 I3_|_SPL_B|D2 I3_|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_B|2|P I3_|_SPL_B|2|MID_SERIES 0  2e-13
RI3_|_SPL_B|2|B I3_|_SPL_B|D2 I3_|_SPL_B|2|MID_SHUNT  2.7439617672
LI3_|_SPL_B|2|RB I3_|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI3_|_SPL_B|A|1 I3_|_SPL_B|QA1 I3_|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_B|A|P I3_|_SPL_B|A|MID_SERIES 0  2e-13
RI3_|_SPL_B|A|B I3_|_SPL_B|QA1 I3_|_SPL_B|A|MID_SHUNT  2.7439617672
LI3_|_SPL_B|A|RB I3_|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI3_|_SPL_B|B|1 I3_|_SPL_B|QB1 I3_|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI3_|_SPL_B|B|P I3_|_SPL_B|B|MID_SERIES 0  2e-13
RI3_|_SPL_B|B|B I3_|_SPL_B|QB1 I3_|_SPL_B|B|MID_SHUNT  2.7439617672
LI3_|_SPL_B|B|RB I3_|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI3_|_DFF_A|I_1|B I3_|_DFF_A|A1 I3_|_DFF_A|I_1|MID  2e-12
II3_|_DFF_A|I_1|B 0 I3_|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_DFF_A|I_3|B I3_|_DFF_A|A3 I3_|_DFF_A|I_3|MID  2e-12
II3_|_DFF_A|I_3|B 0 I3_|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3_|_DFF_A|I_T|B I3_|_DFF_A|T1 I3_|_DFF_A|I_T|MID  2e-12
II3_|_DFF_A|I_T|B 0 I3_|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3_|_DFF_A|I_6|B I3_|_DFF_A|Q1 I3_|_DFF_A|I_6|MID  2e-12
II3_|_DFF_A|I_6|B 0 I3_|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3_|_DFF_A|1|1 I3_|_DFF_A|A1 I3_|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_A|1|P I3_|_DFF_A|1|MID_SERIES 0  2e-13
RI3_|_DFF_A|1|B I3_|_DFF_A|A1 I3_|_DFF_A|1|MID_SHUNT  2.7439617672
LI3_|_DFF_A|1|RB I3_|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_A|23|1 I3_|_DFF_A|A2 I3_|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI3_|_DFF_A|23|B I3_|_DFF_A|A2 I3_|_DFF_A|23|MID_SHUNT  3.84154647408
LI3_|_DFF_A|23|RB I3_|_DFF_A|23|MID_SHUNT I3_|_DFF_A|A3  2.1704737578552e-12
BI3_|_DFF_A|3|1 I3_|_DFF_A|A3 I3_|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_A|3|P I3_|_DFF_A|3|MID_SERIES 0  2e-13
RI3_|_DFF_A|3|B I3_|_DFF_A|A3 I3_|_DFF_A|3|MID_SHUNT  2.7439617672
LI3_|_DFF_A|3|RB I3_|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_A|4|1 I3_|_DFF_A|A4 I3_|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_A|4|P I3_|_DFF_A|4|MID_SERIES 0  2e-13
RI3_|_DFF_A|4|B I3_|_DFF_A|A4 I3_|_DFF_A|4|MID_SHUNT  2.7439617672
LI3_|_DFF_A|4|RB I3_|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_A|T|1 I3_|_DFF_A|T1 I3_|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_A|T|P I3_|_DFF_A|T|MID_SERIES 0  2e-13
RI3_|_DFF_A|T|B I3_|_DFF_A|T1 I3_|_DFF_A|T|MID_SHUNT  2.7439617672
LI3_|_DFF_A|T|RB I3_|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_A|45|1 I3_|_DFF_A|T2 I3_|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI3_|_DFF_A|45|B I3_|_DFF_A|T2 I3_|_DFF_A|45|MID_SHUNT  3.84154647408
LI3_|_DFF_A|45|RB I3_|_DFF_A|45|MID_SHUNT I3_|_DFF_A|A4  2.1704737578552e-12
BI3_|_DFF_A|6|1 I3_|_DFF_A|Q1 I3_|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_A|6|P I3_|_DFF_A|6|MID_SERIES 0  2e-13
RI3_|_DFF_A|6|B I3_|_DFF_A|Q1 I3_|_DFF_A|6|MID_SHUNT  2.7439617672
LI3_|_DFF_A|6|RB I3_|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI3_|_DFF_B|I_1|B I3_|_DFF_B|A1 I3_|_DFF_B|I_1|MID  2e-12
II3_|_DFF_B|I_1|B 0 I3_|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_DFF_B|I_3|B I3_|_DFF_B|A3 I3_|_DFF_B|I_3|MID  2e-12
II3_|_DFF_B|I_3|B 0 I3_|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3_|_DFF_B|I_T|B I3_|_DFF_B|T1 I3_|_DFF_B|I_T|MID  2e-12
II3_|_DFF_B|I_T|B 0 I3_|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3_|_DFF_B|I_6|B I3_|_DFF_B|Q1 I3_|_DFF_B|I_6|MID  2e-12
II3_|_DFF_B|I_6|B 0 I3_|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3_|_DFF_B|1|1 I3_|_DFF_B|A1 I3_|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_B|1|P I3_|_DFF_B|1|MID_SERIES 0  2e-13
RI3_|_DFF_B|1|B I3_|_DFF_B|A1 I3_|_DFF_B|1|MID_SHUNT  2.7439617672
LI3_|_DFF_B|1|RB I3_|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_B|23|1 I3_|_DFF_B|A2 I3_|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI3_|_DFF_B|23|B I3_|_DFF_B|A2 I3_|_DFF_B|23|MID_SHUNT  3.84154647408
LI3_|_DFF_B|23|RB I3_|_DFF_B|23|MID_SHUNT I3_|_DFF_B|A3  2.1704737578552e-12
BI3_|_DFF_B|3|1 I3_|_DFF_B|A3 I3_|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_B|3|P I3_|_DFF_B|3|MID_SERIES 0  2e-13
RI3_|_DFF_B|3|B I3_|_DFF_B|A3 I3_|_DFF_B|3|MID_SHUNT  2.7439617672
LI3_|_DFF_B|3|RB I3_|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_B|4|1 I3_|_DFF_B|A4 I3_|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_B|4|P I3_|_DFF_B|4|MID_SERIES 0  2e-13
RI3_|_DFF_B|4|B I3_|_DFF_B|A4 I3_|_DFF_B|4|MID_SHUNT  2.7439617672
LI3_|_DFF_B|4|RB I3_|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_B|T|1 I3_|_DFF_B|T1 I3_|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_B|T|P I3_|_DFF_B|T|MID_SERIES 0  2e-13
RI3_|_DFF_B|T|B I3_|_DFF_B|T1 I3_|_DFF_B|T|MID_SHUNT  2.7439617672
LI3_|_DFF_B|T|RB I3_|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI3_|_DFF_B|45|1 I3_|_DFF_B|T2 I3_|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI3_|_DFF_B|45|B I3_|_DFF_B|T2 I3_|_DFF_B|45|MID_SHUNT  3.84154647408
LI3_|_DFF_B|45|RB I3_|_DFF_B|45|MID_SHUNT I3_|_DFF_B|A4  2.1704737578552e-12
BI3_|_DFF_B|6|1 I3_|_DFF_B|Q1 I3_|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI3_|_DFF_B|6|P I3_|_DFF_B|6|MID_SERIES 0  2e-13
RI3_|_DFF_B|6|B I3_|_DFF_B|Q1 I3_|_DFF_B|6|MID_SHUNT  2.7439617672
LI3_|_DFF_B|6|RB I3_|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI3_|_XOR|I_A1|B I3_|_XOR|A1 I3_|_XOR|I_A1|MID  2e-12
II3_|_XOR|I_A1|B 0 I3_|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_XOR|I_A3|B I3_|_XOR|A3 I3_|_XOR|I_A3|MID  2e-12
II3_|_XOR|I_A3|B 0 I3_|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI3_|_XOR|I_B1|B I3_|_XOR|B1 I3_|_XOR|I_B1|MID  2e-12
II3_|_XOR|I_B1|B 0 I3_|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_XOR|I_B3|B I3_|_XOR|B3 I3_|_XOR|I_B3|MID  2e-12
II3_|_XOR|I_B3|B 0 I3_|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI3_|_XOR|I_Q1|B I3_|_XOR|Q1 I3_|_XOR|I_Q1|MID  2e-12
II3_|_XOR|I_Q1|B 0 I3_|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3_|_XOR|A1|1 I3_|_XOR|A1 I3_|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|A1|P I3_|_XOR|A1|MID_SERIES 0  5e-13
RI3_|_XOR|A1|B I3_|_XOR|A1 I3_|_XOR|A1|MID_SHUNT  2.7439617672
LI3_|_XOR|A1|RB I3_|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI3_|_XOR|A2|1 I3_|_XOR|A2 I3_|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|A2|P I3_|_XOR|A2|MID_SERIES 0  5e-13
RI3_|_XOR|A2|B I3_|_XOR|A2 I3_|_XOR|A2|MID_SHUNT  2.7439617672
LI3_|_XOR|A2|RB I3_|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI3_|_XOR|A3|1 I3_|_XOR|A2 I3_|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|A3|P I3_|_XOR|A3|MID_SERIES I3_|_XOR|A3  1.2e-12
RI3_|_XOR|A3|B I3_|_XOR|A2 I3_|_XOR|A3|MID_SHUNT  2.7439617672
LI3_|_XOR|A3|RB I3_|_XOR|A3|MID_SHUNT I3_|_XOR|A3  2.050338398468e-12
BI3_|_XOR|B1|1 I3_|_XOR|B1 I3_|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|B1|P I3_|_XOR|B1|MID_SERIES 0  5e-13
RI3_|_XOR|B1|B I3_|_XOR|B1 I3_|_XOR|B1|MID_SHUNT  2.7439617672
LI3_|_XOR|B1|RB I3_|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI3_|_XOR|B2|1 I3_|_XOR|B2 I3_|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|B2|P I3_|_XOR|B2|MID_SERIES 0  5e-13
RI3_|_XOR|B2|B I3_|_XOR|B2 I3_|_XOR|B2|MID_SHUNT  2.7439617672
LI3_|_XOR|B2|RB I3_|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI3_|_XOR|B3|1 I3_|_XOR|B2 I3_|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|B3|P I3_|_XOR|B3|MID_SERIES I3_|_XOR|B3  1.2e-12
RI3_|_XOR|B3|B I3_|_XOR|B2 I3_|_XOR|B3|MID_SHUNT  2.7439617672
LI3_|_XOR|B3|RB I3_|_XOR|B3|MID_SHUNT I3_|_XOR|B3  2.050338398468e-12
BI3_|_XOR|T1|1 I3_|_XOR|T1 I3_|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|T1|P I3_|_XOR|T1|MID_SERIES 0  5e-13
RI3_|_XOR|T1|B I3_|_XOR|T1 I3_|_XOR|T1|MID_SHUNT  2.7439617672
LI3_|_XOR|T1|RB I3_|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI3_|_XOR|T2|1 I3_|_XOR|T2 I3_|_XOR|ABTQ JJMIT AREA=2.0
RI3_|_XOR|T2|B I3_|_XOR|T2 I3_|_XOR|T2|MID_SHUNT  3.429952209
LI3_|_XOR|T2|RB I3_|_XOR|T2|MID_SHUNT I3_|_XOR|ABTQ  2.437922998085e-12
BI3_|_XOR|AB|1 I3_|_XOR|AB I3_|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI3_|_XOR|AB|P I3_|_XOR|AB|MID_SERIES I3_|_XOR|ABTQ  1.2e-12
RI3_|_XOR|AB|B I3_|_XOR|AB I3_|_XOR|AB|MID_SHUNT  3.429952209
LI3_|_XOR|AB|RB I3_|_XOR|AB|MID_SHUNT I3_|_XOR|ABTQ  2.437922998085e-12
BI3_|_XOR|ABTQ|1 I3_|_XOR|ABTQ I3_|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|ABTQ|P I3_|_XOR|ABTQ|MID_SERIES 0  5e-13
RI3_|_XOR|ABTQ|B I3_|_XOR|ABTQ I3_|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI3_|_XOR|ABTQ|RB I3_|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI3_|_XOR|Q1|1 I3_|_XOR|Q1 I3_|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI3_|_XOR|Q1|P I3_|_XOR|Q1|MID_SERIES 0  5e-13
RI3_|_XOR|Q1|B I3_|_XOR|Q1 I3_|_XOR|Q1|MID_SHUNT  2.7439617672
LI3_|_XOR|Q1|RB I3_|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI3_|_AND|I_A1|B I3_|_AND|A1 I3_|_AND|I_A1|MID  2e-12
II3_|_AND|I_A1|B 0 I3_|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_AND|I_B1|B I3_|_AND|B1 I3_|_AND|I_B1|MID  2e-12
II3_|_AND|I_B1|B 0 I3_|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3_|_AND|I_Q3|B I3_|_AND|Q3 I3_|_AND|I_Q3|MID  2e-12
II3_|_AND|I_Q3|B 0 I3_|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3_|_AND|I_Q2|B I3_|_AND|Q2 I3_|_AND|I_Q2|MID  2e-12
II3_|_AND|I_Q2|B 0 I3_|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3_|_AND|I_Q1|B I3_|_AND|Q1 I3_|_AND|I_Q1|MID  2e-12
II3_|_AND|I_Q1|B 0 I3_|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3_|_AND|A1|1 I3_|_AND|A1 I3_|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3_|_AND|A1|P I3_|_AND|A1|MID_SERIES 0  2e-13
RI3_|_AND|A1|B I3_|_AND|A1 I3_|_AND|A1|MID_SHUNT  2.7439617672
LI3_|_AND|A1|RB I3_|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3_|_AND|A2|1 I3_|_AND|A2 I3_|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3_|_AND|A2|P I3_|_AND|A2|MID_SERIES 0  2e-13
RI3_|_AND|A2|B I3_|_AND|A2 I3_|_AND|A2|MID_SHUNT  2.7439617672
LI3_|_AND|A2|RB I3_|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3_|_AND|A12|1 I3_|_AND|A2 I3_|_AND|A3 JJMIT AREA=1.7857142857142858
RI3_|_AND|A12|B I3_|_AND|A2 I3_|_AND|A12|MID_SHUNT  3.84154647408
LI3_|_AND|A12|RB I3_|_AND|A12|MID_SHUNT I3_|_AND|A3  2.1704737578552e-12
BI3_|_AND|B1|1 I3_|_AND|B1 I3_|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3_|_AND|B1|P I3_|_AND|B1|MID_SERIES 0  2e-13
RI3_|_AND|B1|B I3_|_AND|B1 I3_|_AND|B1|MID_SHUNT  2.7439617672
LI3_|_AND|B1|RB I3_|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3_|_AND|B2|1 I3_|_AND|B2 I3_|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3_|_AND|B2|P I3_|_AND|B2|MID_SERIES 0  2e-13
RI3_|_AND|B2|B I3_|_AND|B2 I3_|_AND|B2|MID_SHUNT  2.7439617672
LI3_|_AND|B2|RB I3_|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3_|_AND|B12|1 I3_|_AND|B2 I3_|_AND|B3 JJMIT AREA=1.7857142857142858
RI3_|_AND|B12|B I3_|_AND|B2 I3_|_AND|B12|MID_SHUNT  3.84154647408
LI3_|_AND|B12|RB I3_|_AND|B12|MID_SHUNT I3_|_AND|B3  2.1704737578552e-12
BI3_|_AND|Q2|1 I3_|_AND|Q2 I3_|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3_|_AND|Q2|P I3_|_AND|Q2|MID_SERIES 0  2e-13
RI3_|_AND|Q2|B I3_|_AND|Q2 I3_|_AND|Q2|MID_SHUNT  2.7439617672
LI3_|_AND|Q2|RB I3_|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3_|_AND|Q1|1 I3_|_AND|Q1 I3_|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3_|_AND|Q1|P I3_|_AND|Q1|MID_SERIES 0  2e-13
RI3_|_AND|Q1|B I3_|_AND|Q1 I3_|_AND|Q1|MID_SHUNT  2.7439617672
LI3_|_AND|Q1|RB I3_|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0_|SPL1|I_D1|B SPL_IP2_0_|SPL1|D1 SPL_IP2_0_|SPL1|I_D1|MID  2e-12
ISPL_IP2_0_|SPL1|I_D1|B 0 SPL_IP2_0_|SPL1|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0_|SPL1|I_D2|B SPL_IP2_0_|SPL1|D2 SPL_IP2_0_|SPL1|I_D2|MID  2e-12
ISPL_IP2_0_|SPL1|I_D2|B 0 SPL_IP2_0_|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IP2_0_|SPL1|I_Q1|B SPL_IP2_0_|SPL1|QA1 SPL_IP2_0_|SPL1|I_Q1|MID  2e-12
ISPL_IP2_0_|SPL1|I_Q1|B 0 SPL_IP2_0_|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0_|SPL1|I_Q2|B SPL_IP2_0_|SPL1|QB1 SPL_IP2_0_|SPL1|I_Q2|MID  2e-12
ISPL_IP2_0_|SPL1|I_Q2|B 0 SPL_IP2_0_|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IP2_0_|SPL1|1|1 SPL_IP2_0_|SPL1|D1 SPL_IP2_0_|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL1|1|P SPL_IP2_0_|SPL1|1|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL1|1|B SPL_IP2_0_|SPL1|D1 SPL_IP2_0_|SPL1|1|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL1|1|RB SPL_IP2_0_|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0_|SPL1|2|1 SPL_IP2_0_|SPL1|D2 SPL_IP2_0_|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL1|2|P SPL_IP2_0_|SPL1|2|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL1|2|B SPL_IP2_0_|SPL1|D2 SPL_IP2_0_|SPL1|2|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL1|2|RB SPL_IP2_0_|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0_|SPL1|A|1 SPL_IP2_0_|SPL1|QA1 SPL_IP2_0_|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL1|A|P SPL_IP2_0_|SPL1|A|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL1|A|B SPL_IP2_0_|SPL1|QA1 SPL_IP2_0_|SPL1|A|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL1|A|RB SPL_IP2_0_|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0_|SPL1|B|1 SPL_IP2_0_|SPL1|QB1 SPL_IP2_0_|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL1|B|P SPL_IP2_0_|SPL1|B|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL1|B|B SPL_IP2_0_|SPL1|QB1 SPL_IP2_0_|SPL1|B|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL1|B|RB SPL_IP2_0_|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0_|SPL2|I_D1|B SPL_IP2_0_|SPL2|D1 SPL_IP2_0_|SPL2|I_D1|MID  2e-12
ISPL_IP2_0_|SPL2|I_D1|B 0 SPL_IP2_0_|SPL2|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0_|SPL2|I_D2|B SPL_IP2_0_|SPL2|D2 SPL_IP2_0_|SPL2|I_D2|MID  2e-12
ISPL_IP2_0_|SPL2|I_D2|B 0 SPL_IP2_0_|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_IP2_0_|SPL2|I_Q1|B SPL_IP2_0_|SPL2|QA1 SPL_IP2_0_|SPL2|I_Q1|MID  2e-12
ISPL_IP2_0_|SPL2|I_Q1|B 0 SPL_IP2_0_|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_IP2_0_|SPL2|I_Q2|B SPL_IP2_0_|SPL2|QB1 SPL_IP2_0_|SPL2|I_Q2|MID  2e-12
ISPL_IP2_0_|SPL2|I_Q2|B 0 SPL_IP2_0_|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_IP2_0_|SPL2|1|1 SPL_IP2_0_|SPL2|D1 SPL_IP2_0_|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL2|1|P SPL_IP2_0_|SPL2|1|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL2|1|B SPL_IP2_0_|SPL2|D1 SPL_IP2_0_|SPL2|1|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL2|1|RB SPL_IP2_0_|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0_|SPL2|2|1 SPL_IP2_0_|SPL2|D2 SPL_IP2_0_|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL2|2|P SPL_IP2_0_|SPL2|2|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL2|2|B SPL_IP2_0_|SPL2|D2 SPL_IP2_0_|SPL2|2|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL2|2|RB SPL_IP2_0_|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0_|SPL2|A|1 SPL_IP2_0_|SPL2|QA1 SPL_IP2_0_|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL2|A|P SPL_IP2_0_|SPL2|A|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL2|A|B SPL_IP2_0_|SPL2|QA1 SPL_IP2_0_|SPL2|A|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL2|A|RB SPL_IP2_0_|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0_|SPL2|B|1 SPL_IP2_0_|SPL2|QB1 SPL_IP2_0_|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0_|SPL2|B|P SPL_IP2_0_|SPL2|B|MID_SERIES 0  2e-13
RSPL_IP2_0_|SPL2|B|B SPL_IP2_0_|SPL2|QB1 SPL_IP2_0_|SPL2|B|MID_SHUNT  2.7439617672
LSPL_IP2_0_|SPL2|B|RB SPL_IP2_0_|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01_|P|I_1|B _PG0_01_|P|A1 _PG0_01_|P|I_1|MID  2e-12
I_PG0_01_|P|I_1|B 0 _PG0_01_|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01_|P|I_3|B _PG0_01_|P|A3 _PG0_01_|P|I_3|MID  2e-12
I_PG0_01_|P|I_3|B 0 _PG0_01_|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01_|P|I_T|B _PG0_01_|P|T1 _PG0_01_|P|I_T|MID  2e-12
I_PG0_01_|P|I_T|B 0 _PG0_01_|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01_|P|I_6|B _PG0_01_|P|Q1 _PG0_01_|P|I_6|MID  2e-12
I_PG0_01_|P|I_6|B 0 _PG0_01_|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01_|P|1|1 _PG0_01_|P|A1 _PG0_01_|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|P|1|P _PG0_01_|P|1|MID_SERIES 0  2e-13
R_PG0_01_|P|1|B _PG0_01_|P|A1 _PG0_01_|P|1|MID_SHUNT  2.7439617672
L_PG0_01_|P|1|RB _PG0_01_|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|P|23|1 _PG0_01_|P|A2 _PG0_01_|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_01_|P|23|B _PG0_01_|P|A2 _PG0_01_|P|23|MID_SHUNT  3.84154647408
L_PG0_01_|P|23|RB _PG0_01_|P|23|MID_SHUNT _PG0_01_|P|A3  2.1704737578552e-12
B_PG0_01_|P|3|1 _PG0_01_|P|A3 _PG0_01_|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|P|3|P _PG0_01_|P|3|MID_SERIES 0  2e-13
R_PG0_01_|P|3|B _PG0_01_|P|A3 _PG0_01_|P|3|MID_SHUNT  2.7439617672
L_PG0_01_|P|3|RB _PG0_01_|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|P|4|1 _PG0_01_|P|A4 _PG0_01_|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|P|4|P _PG0_01_|P|4|MID_SERIES 0  2e-13
R_PG0_01_|P|4|B _PG0_01_|P|A4 _PG0_01_|P|4|MID_SHUNT  2.7439617672
L_PG0_01_|P|4|RB _PG0_01_|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|P|T|1 _PG0_01_|P|T1 _PG0_01_|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|P|T|P _PG0_01_|P|T|MID_SERIES 0  2e-13
R_PG0_01_|P|T|B _PG0_01_|P|T1 _PG0_01_|P|T|MID_SHUNT  2.7439617672
L_PG0_01_|P|T|RB _PG0_01_|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|P|45|1 _PG0_01_|P|T2 _PG0_01_|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_01_|P|45|B _PG0_01_|P|T2 _PG0_01_|P|45|MID_SHUNT  3.84154647408
L_PG0_01_|P|45|RB _PG0_01_|P|45|MID_SHUNT _PG0_01_|P|A4  2.1704737578552e-12
B_PG0_01_|P|6|1 _PG0_01_|P|Q1 _PG0_01_|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|P|6|P _PG0_01_|P|6|MID_SERIES 0  2e-13
R_PG0_01_|P|6|B _PG0_01_|P|Q1 _PG0_01_|P|6|MID_SHUNT  2.7439617672
L_PG0_01_|P|6|RB _PG0_01_|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_01_|G|I_1|B _PG0_01_|G|A1 _PG0_01_|G|I_1|MID  2e-12
I_PG0_01_|G|I_1|B 0 _PG0_01_|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01_|G|I_3|B _PG0_01_|G|A3 _PG0_01_|G|I_3|MID  2e-12
I_PG0_01_|G|I_3|B 0 _PG0_01_|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01_|G|I_T|B _PG0_01_|G|T1 _PG0_01_|G|I_T|MID  2e-12
I_PG0_01_|G|I_T|B 0 _PG0_01_|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01_|G|I_6|B _PG0_01_|G|Q1 _PG0_01_|G|I_6|MID  2e-12
I_PG0_01_|G|I_6|B 0 _PG0_01_|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01_|G|1|1 _PG0_01_|G|A1 _PG0_01_|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|G|1|P _PG0_01_|G|1|MID_SERIES 0  2e-13
R_PG0_01_|G|1|B _PG0_01_|G|A1 _PG0_01_|G|1|MID_SHUNT  2.7439617672
L_PG0_01_|G|1|RB _PG0_01_|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|G|23|1 _PG0_01_|G|A2 _PG0_01_|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_01_|G|23|B _PG0_01_|G|A2 _PG0_01_|G|23|MID_SHUNT  3.84154647408
L_PG0_01_|G|23|RB _PG0_01_|G|23|MID_SHUNT _PG0_01_|G|A3  2.1704737578552e-12
B_PG0_01_|G|3|1 _PG0_01_|G|A3 _PG0_01_|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|G|3|P _PG0_01_|G|3|MID_SERIES 0  2e-13
R_PG0_01_|G|3|B _PG0_01_|G|A3 _PG0_01_|G|3|MID_SHUNT  2.7439617672
L_PG0_01_|G|3|RB _PG0_01_|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|G|4|1 _PG0_01_|G|A4 _PG0_01_|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|G|4|P _PG0_01_|G|4|MID_SERIES 0  2e-13
R_PG0_01_|G|4|B _PG0_01_|G|A4 _PG0_01_|G|4|MID_SHUNT  2.7439617672
L_PG0_01_|G|4|RB _PG0_01_|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|G|T|1 _PG0_01_|G|T1 _PG0_01_|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|G|T|P _PG0_01_|G|T|MID_SERIES 0  2e-13
R_PG0_01_|G|T|B _PG0_01_|G|T1 _PG0_01_|G|T|MID_SHUNT  2.7439617672
L_PG0_01_|G|T|RB _PG0_01_|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01_|G|45|1 _PG0_01_|G|T2 _PG0_01_|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_01_|G|45|B _PG0_01_|G|T2 _PG0_01_|G|45|MID_SHUNT  3.84154647408
L_PG0_01_|G|45|RB _PG0_01_|G|45|MID_SHUNT _PG0_01_|G|A4  2.1704737578552e-12
B_PG0_01_|G|6|1 _PG0_01_|G|Q1 _PG0_01_|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01_|G|6|P _PG0_01_|G|6|MID_SERIES 0  2e-13
R_PG0_01_|G|6|B _PG0_01_|G|Q1 _PG0_01_|G|6|MID_SHUNT  2.7439617672
L_PG0_01_|G|6|RB _PG0_01_|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01_|_SPL_G1|I_D1|B _PG1_01_|_SPL_G1|D1 _PG1_01_|_SPL_G1|I_D1|MID  2e-12
I_PG1_01_|_SPL_G1|I_D1|B 0 _PG1_01_|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_SPL_G1|I_D2|B _PG1_01_|_SPL_G1|D2 _PG1_01_|_SPL_G1|I_D2|MID  2e-12
I_PG1_01_|_SPL_G1|I_D2|B 0 _PG1_01_|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PG1_01_|_SPL_G1|I_Q1|B _PG1_01_|_SPL_G1|QA1 _PG1_01_|_SPL_G1|I_Q1|MID  2e-12
I_PG1_01_|_SPL_G1|I_Q1|B 0 _PG1_01_|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_SPL_G1|I_Q2|B _PG1_01_|_SPL_G1|QB1 _PG1_01_|_SPL_G1|I_Q2|MID  2e-12
I_PG1_01_|_SPL_G1|I_Q2|B 0 _PG1_01_|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01_|_SPL_G1|1|1 _PG1_01_|_SPL_G1|D1 _PG1_01_|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_SPL_G1|1|P _PG1_01_|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG1_01_|_SPL_G1|1|B _PG1_01_|_SPL_G1|D1 _PG1_01_|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG1_01_|_SPL_G1|1|RB _PG1_01_|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_SPL_G1|2|1 _PG1_01_|_SPL_G1|D2 _PG1_01_|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_SPL_G1|2|P _PG1_01_|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG1_01_|_SPL_G1|2|B _PG1_01_|_SPL_G1|D2 _PG1_01_|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG1_01_|_SPL_G1|2|RB _PG1_01_|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_SPL_G1|A|1 _PG1_01_|_SPL_G1|QA1 _PG1_01_|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_SPL_G1|A|P _PG1_01_|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG1_01_|_SPL_G1|A|B _PG1_01_|_SPL_G1|QA1 _PG1_01_|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG1_01_|_SPL_G1|A|RB _PG1_01_|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_SPL_G1|B|1 _PG1_01_|_SPL_G1|QB1 _PG1_01_|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_SPL_G1|B|P _PG1_01_|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG1_01_|_SPL_G1|B|B _PG1_01_|_SPL_G1|QB1 _PG1_01_|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG1_01_|_SPL_G1|B|RB _PG1_01_|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01_|_PG|I_A1|B _PG1_01_|_PG|A1 _PG1_01_|_PG|I_A1|MID  2e-12
I_PG1_01_|_PG|I_A1|B 0 _PG1_01_|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_PG|I_B1|B _PG1_01_|_PG|B1 _PG1_01_|_PG|I_B1|MID  2e-12
I_PG1_01_|_PG|I_B1|B 0 _PG1_01_|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_PG|I_Q3|B _PG1_01_|_PG|Q3 _PG1_01_|_PG|I_Q3|MID  2e-12
I_PG1_01_|_PG|I_Q3|B 0 _PG1_01_|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01_|_PG|I_Q2|B _PG1_01_|_PG|Q2 _PG1_01_|_PG|I_Q2|MID  2e-12
I_PG1_01_|_PG|I_Q2|B 0 _PG1_01_|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_PG|I_Q1|B _PG1_01_|_PG|Q1 _PG1_01_|_PG|I_Q1|MID  2e-12
I_PG1_01_|_PG|I_Q1|B 0 _PG1_01_|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01_|_PG|A1|1 _PG1_01_|_PG|A1 _PG1_01_|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_PG|A1|P _PG1_01_|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01_|_PG|A1|B _PG1_01_|_PG|A1 _PG1_01_|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01_|_PG|A1|RB _PG1_01_|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_PG|A2|1 _PG1_01_|_PG|A2 _PG1_01_|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_PG|A2|P _PG1_01_|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01_|_PG|A2|B _PG1_01_|_PG|A2 _PG1_01_|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01_|_PG|A2|RB _PG1_01_|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_PG|A12|1 _PG1_01_|_PG|A2 _PG1_01_|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_PG|A12|B _PG1_01_|_PG|A2 _PG1_01_|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01_|_PG|A12|RB _PG1_01_|_PG|A12|MID_SHUNT _PG1_01_|_PG|A3  2.1704737578552e-12
B_PG1_01_|_PG|B1|1 _PG1_01_|_PG|B1 _PG1_01_|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_PG|B1|P _PG1_01_|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01_|_PG|B1|B _PG1_01_|_PG|B1 _PG1_01_|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01_|_PG|B1|RB _PG1_01_|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_PG|B2|1 _PG1_01_|_PG|B2 _PG1_01_|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_PG|B2|P _PG1_01_|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01_|_PG|B2|B _PG1_01_|_PG|B2 _PG1_01_|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01_|_PG|B2|RB _PG1_01_|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_PG|B12|1 _PG1_01_|_PG|B2 _PG1_01_|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_PG|B12|B _PG1_01_|_PG|B2 _PG1_01_|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01_|_PG|B12|RB _PG1_01_|_PG|B12|MID_SHUNT _PG1_01_|_PG|B3  2.1704737578552e-12
B_PG1_01_|_PG|Q2|1 _PG1_01_|_PG|Q2 _PG1_01_|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_PG|Q2|P _PG1_01_|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01_|_PG|Q2|B _PG1_01_|_PG|Q2 _PG1_01_|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01_|_PG|Q2|RB _PG1_01_|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_PG|Q1|1 _PG1_01_|_PG|Q1 _PG1_01_|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_PG|Q1|P _PG1_01_|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01_|_PG|Q1|B _PG1_01_|_PG|Q1 _PG1_01_|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01_|_PG|Q1|RB _PG1_01_|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01_|_GG|I_A1|B _PG1_01_|_GG|A1 _PG1_01_|_GG|I_A1|MID  2e-12
I_PG1_01_|_GG|I_A1|B 0 _PG1_01_|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_GG|I_B1|B _PG1_01_|_GG|B1 _PG1_01_|_GG|I_B1|MID  2e-12
I_PG1_01_|_GG|I_B1|B 0 _PG1_01_|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_GG|I_Q3|B _PG1_01_|_GG|Q3 _PG1_01_|_GG|I_Q3|MID  2e-12
I_PG1_01_|_GG|I_Q3|B 0 _PG1_01_|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01_|_GG|I_Q2|B _PG1_01_|_GG|Q2 _PG1_01_|_GG|I_Q2|MID  2e-12
I_PG1_01_|_GG|I_Q2|B 0 _PG1_01_|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_GG|I_Q1|B _PG1_01_|_GG|Q1 _PG1_01_|_GG|I_Q1|MID  2e-12
I_PG1_01_|_GG|I_Q1|B 0 _PG1_01_|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01_|_GG|A1|1 _PG1_01_|_GG|A1 _PG1_01_|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_GG|A1|P _PG1_01_|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01_|_GG|A1|B _PG1_01_|_GG|A1 _PG1_01_|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01_|_GG|A1|RB _PG1_01_|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_GG|A2|1 _PG1_01_|_GG|A2 _PG1_01_|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_GG|A2|P _PG1_01_|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01_|_GG|A2|B _PG1_01_|_GG|A2 _PG1_01_|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01_|_GG|A2|RB _PG1_01_|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_GG|A12|1 _PG1_01_|_GG|A2 _PG1_01_|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_GG|A12|B _PG1_01_|_GG|A2 _PG1_01_|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01_|_GG|A12|RB _PG1_01_|_GG|A12|MID_SHUNT _PG1_01_|_GG|A3  2.1704737578552e-12
B_PG1_01_|_GG|B1|1 _PG1_01_|_GG|B1 _PG1_01_|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_GG|B1|P _PG1_01_|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01_|_GG|B1|B _PG1_01_|_GG|B1 _PG1_01_|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01_|_GG|B1|RB _PG1_01_|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_GG|B2|1 _PG1_01_|_GG|B2 _PG1_01_|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_GG|B2|P _PG1_01_|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01_|_GG|B2|B _PG1_01_|_GG|B2 _PG1_01_|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01_|_GG|B2|RB _PG1_01_|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_GG|B12|1 _PG1_01_|_GG|B2 _PG1_01_|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_GG|B12|B _PG1_01_|_GG|B2 _PG1_01_|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01_|_GG|B12|RB _PG1_01_|_GG|B12|MID_SHUNT _PG1_01_|_GG|B3  2.1704737578552e-12
B_PG1_01_|_GG|Q2|1 _PG1_01_|_GG|Q2 _PG1_01_|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_GG|Q2|P _PG1_01_|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01_|_GG|Q2|B _PG1_01_|_GG|Q2 _PG1_01_|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01_|_GG|Q2|RB _PG1_01_|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_GG|Q1|1 _PG1_01_|_GG|Q1 _PG1_01_|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_GG|Q1|P _PG1_01_|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01_|_GG|Q1|B _PG1_01_|_GG|Q1 _PG1_01_|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01_|_GG|Q1|RB _PG1_01_|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01_|_DFF_PG|I_1|B _PG1_01_|_DFF_PG|A1 _PG1_01_|_DFF_PG|I_1|MID  2e-12
I_PG1_01_|_DFF_PG|I_1|B 0 _PG1_01_|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_DFF_PG|I_3|B _PG1_01_|_DFF_PG|A3 _PG1_01_|_DFF_PG|I_3|MID  2e-12
I_PG1_01_|_DFF_PG|I_3|B 0 _PG1_01_|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01_|_DFF_PG|I_T|B _PG1_01_|_DFF_PG|T1 _PG1_01_|_DFF_PG|I_T|MID  2e-12
I_PG1_01_|_DFF_PG|I_T|B 0 _PG1_01_|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_DFF_PG|I_6|B _PG1_01_|_DFF_PG|Q1 _PG1_01_|_DFF_PG|I_6|MID  2e-12
I_PG1_01_|_DFF_PG|I_6|B 0 _PG1_01_|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01_|_DFF_PG|1|1 _PG1_01_|_DFF_PG|A1 _PG1_01_|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_PG|1|P _PG1_01_|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_PG|1|B _PG1_01_|_DFF_PG|A1 _PG1_01_|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_PG|1|RB _PG1_01_|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_PG|23|1 _PG1_01_|_DFF_PG|A2 _PG1_01_|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_DFF_PG|23|B _PG1_01_|_DFF_PG|A2 _PG1_01_|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG1_01_|_DFF_PG|23|RB _PG1_01_|_DFF_PG|23|MID_SHUNT _PG1_01_|_DFF_PG|A3  2.1704737578552e-12
B_PG1_01_|_DFF_PG|3|1 _PG1_01_|_DFF_PG|A3 _PG1_01_|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_PG|3|P _PG1_01_|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_PG|3|B _PG1_01_|_DFF_PG|A3 _PG1_01_|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_PG|3|RB _PG1_01_|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_PG|4|1 _PG1_01_|_DFF_PG|A4 _PG1_01_|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_PG|4|P _PG1_01_|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_PG|4|B _PG1_01_|_DFF_PG|A4 _PG1_01_|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_PG|4|RB _PG1_01_|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_PG|T|1 _PG1_01_|_DFF_PG|T1 _PG1_01_|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_PG|T|P _PG1_01_|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_PG|T|B _PG1_01_|_DFF_PG|T1 _PG1_01_|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_PG|T|RB _PG1_01_|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_PG|45|1 _PG1_01_|_DFF_PG|T2 _PG1_01_|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01_|_DFF_PG|45|B _PG1_01_|_DFF_PG|T2 _PG1_01_|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG1_01_|_DFF_PG|45|RB _PG1_01_|_DFF_PG|45|MID_SHUNT _PG1_01_|_DFF_PG|A4  2.1704737578552e-12
B_PG1_01_|_DFF_PG|6|1 _PG1_01_|_DFF_PG|Q1 _PG1_01_|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_PG|6|P _PG1_01_|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_PG|6|B _PG1_01_|_DFF_PG|Q1 _PG1_01_|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_PG|6|RB _PG1_01_|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01_|_DFF_GG|I_1|B _PG1_01_|_DFF_GG|A1 _PG1_01_|_DFF_GG|I_1|MID  2e-12
I_PG1_01_|_DFF_GG|I_1|B 0 _PG1_01_|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_DFF_GG|I_3|B _PG1_01_|_DFF_GG|A3 _PG1_01_|_DFF_GG|I_3|MID  2e-12
I_PG1_01_|_DFF_GG|I_3|B 0 _PG1_01_|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01_|_DFF_GG|I_T|B _PG1_01_|_DFF_GG|T1 _PG1_01_|_DFF_GG|I_T|MID  2e-12
I_PG1_01_|_DFF_GG|I_T|B 0 _PG1_01_|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_DFF_GG|I_6|B _PG1_01_|_DFF_GG|Q1 _PG1_01_|_DFF_GG|I_6|MID  2e-12
I_PG1_01_|_DFF_GG|I_6|B 0 _PG1_01_|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01_|_DFF_GG|1|1 _PG1_01_|_DFF_GG|A1 _PG1_01_|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_GG|1|P _PG1_01_|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_GG|1|B _PG1_01_|_DFF_GG|A1 _PG1_01_|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_GG|1|RB _PG1_01_|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_GG|23|1 _PG1_01_|_DFF_GG|A2 _PG1_01_|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_DFF_GG|23|B _PG1_01_|_DFF_GG|A2 _PG1_01_|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG1_01_|_DFF_GG|23|RB _PG1_01_|_DFF_GG|23|MID_SHUNT _PG1_01_|_DFF_GG|A3  2.1704737578552e-12
B_PG1_01_|_DFF_GG|3|1 _PG1_01_|_DFF_GG|A3 _PG1_01_|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_GG|3|P _PG1_01_|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_GG|3|B _PG1_01_|_DFF_GG|A3 _PG1_01_|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_GG|3|RB _PG1_01_|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_GG|4|1 _PG1_01_|_DFF_GG|A4 _PG1_01_|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_GG|4|P _PG1_01_|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_GG|4|B _PG1_01_|_DFF_GG|A4 _PG1_01_|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_GG|4|RB _PG1_01_|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_GG|T|1 _PG1_01_|_DFF_GG|T1 _PG1_01_|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_GG|T|P _PG1_01_|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_GG|T|B _PG1_01_|_DFF_GG|T1 _PG1_01_|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_GG|T|RB _PG1_01_|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_DFF_GG|45|1 _PG1_01_|_DFF_GG|T2 _PG1_01_|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01_|_DFF_GG|45|B _PG1_01_|_DFF_GG|T2 _PG1_01_|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG1_01_|_DFF_GG|45|RB _PG1_01_|_DFF_GG|45|MID_SHUNT _PG1_01_|_DFF_GG|A4  2.1704737578552e-12
B_PG1_01_|_DFF_GG|6|1 _PG1_01_|_DFF_GG|Q1 _PG1_01_|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_DFF_GG|6|P _PG1_01_|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG1_01_|_DFF_GG|6|B _PG1_01_|_DFF_GG|Q1 _PG1_01_|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG1_01_|_DFF_GG|6|RB _PG1_01_|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01_|_AND_G|I_A1|B _PG1_01_|_AND_G|A1 _PG1_01_|_AND_G|I_A1|MID  2e-12
I_PG1_01_|_AND_G|I_A1|B 0 _PG1_01_|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_AND_G|I_B1|B _PG1_01_|_AND_G|B1 _PG1_01_|_AND_G|I_B1|MID  2e-12
I_PG1_01_|_AND_G|I_B1|B 0 _PG1_01_|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_AND_G|I_Q3|B _PG1_01_|_AND_G|Q3 _PG1_01_|_AND_G|I_Q3|MID  2e-12
I_PG1_01_|_AND_G|I_Q3|B 0 _PG1_01_|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01_|_AND_G|I_Q2|B _PG1_01_|_AND_G|Q2 _PG1_01_|_AND_G|I_Q2|MID  2e-12
I_PG1_01_|_AND_G|I_Q2|B 0 _PG1_01_|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01_|_AND_G|I_Q1|B _PG1_01_|_AND_G|Q1 _PG1_01_|_AND_G|I_Q1|MID  2e-12
I_PG1_01_|_AND_G|I_Q1|B 0 _PG1_01_|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01_|_AND_G|A1|1 _PG1_01_|_AND_G|A1 _PG1_01_|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_AND_G|A1|P _PG1_01_|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01_|_AND_G|A1|B _PG1_01_|_AND_G|A1 _PG1_01_|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01_|_AND_G|A1|RB _PG1_01_|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_AND_G|A2|1 _PG1_01_|_AND_G|A2 _PG1_01_|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_AND_G|A2|P _PG1_01_|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01_|_AND_G|A2|B _PG1_01_|_AND_G|A2 _PG1_01_|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01_|_AND_G|A2|RB _PG1_01_|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_AND_G|A12|1 _PG1_01_|_AND_G|A2 _PG1_01_|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_AND_G|A12|B _PG1_01_|_AND_G|A2 _PG1_01_|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01_|_AND_G|A12|RB _PG1_01_|_AND_G|A12|MID_SHUNT _PG1_01_|_AND_G|A3  2.1704737578552e-12
B_PG1_01_|_AND_G|B1|1 _PG1_01_|_AND_G|B1 _PG1_01_|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_AND_G|B1|P _PG1_01_|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01_|_AND_G|B1|B _PG1_01_|_AND_G|B1 _PG1_01_|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01_|_AND_G|B1|RB _PG1_01_|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_AND_G|B2|1 _PG1_01_|_AND_G|B2 _PG1_01_|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_AND_G|B2|P _PG1_01_|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01_|_AND_G|B2|B _PG1_01_|_AND_G|B2 _PG1_01_|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01_|_AND_G|B2|RB _PG1_01_|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_AND_G|B12|1 _PG1_01_|_AND_G|B2 _PG1_01_|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01_|_AND_G|B12|B _PG1_01_|_AND_G|B2 _PG1_01_|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01_|_AND_G|B12|RB _PG1_01_|_AND_G|B12|MID_SHUNT _PG1_01_|_AND_G|B3  2.1704737578552e-12
B_PG1_01_|_AND_G|Q2|1 _PG1_01_|_AND_G|Q2 _PG1_01_|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_AND_G|Q2|P _PG1_01_|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01_|_AND_G|Q2|B _PG1_01_|_AND_G|Q2 _PG1_01_|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01_|_AND_G|Q2|RB _PG1_01_|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01_|_AND_G|Q1|1 _PG1_01_|_AND_G|Q1 _PG1_01_|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01_|_AND_G|Q1|P _PG1_01_|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01_|_AND_G|Q1|B _PG1_01_|_AND_G|Q1 _PG1_01_|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01_|_AND_G|Q1|RB _PG1_01_|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_01_|P|I_1|B _PG2_01_|P|A1 _PG2_01_|P|I_1|MID  2e-12
I_PG2_01_|P|I_1|B 0 _PG2_01_|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01_|P|I_3|B _PG2_01_|P|A3 _PG2_01_|P|I_3|MID  2e-12
I_PG2_01_|P|I_3|B 0 _PG2_01_|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01_|P|I_T|B _PG2_01_|P|T1 _PG2_01_|P|I_T|MID  2e-12
I_PG2_01_|P|I_T|B 0 _PG2_01_|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01_|P|I_6|B _PG2_01_|P|Q1 _PG2_01_|P|I_6|MID  2e-12
I_PG2_01_|P|I_6|B 0 _PG2_01_|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01_|P|1|1 _PG2_01_|P|A1 _PG2_01_|P|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|P|1|P _PG2_01_|P|1|MID_SERIES 0  2e-13
R_PG2_01_|P|1|B _PG2_01_|P|A1 _PG2_01_|P|1|MID_SHUNT  2.7439617672
L_PG2_01_|P|1|RB _PG2_01_|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|P|23|1 _PG2_01_|P|A2 _PG2_01_|P|A3 JJMIT AREA=1.7857142857142858
R_PG2_01_|P|23|B _PG2_01_|P|A2 _PG2_01_|P|23|MID_SHUNT  3.84154647408
L_PG2_01_|P|23|RB _PG2_01_|P|23|MID_SHUNT _PG2_01_|P|A3  2.1704737578552e-12
B_PG2_01_|P|3|1 _PG2_01_|P|A3 _PG2_01_|P|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|P|3|P _PG2_01_|P|3|MID_SERIES 0  2e-13
R_PG2_01_|P|3|B _PG2_01_|P|A3 _PG2_01_|P|3|MID_SHUNT  2.7439617672
L_PG2_01_|P|3|RB _PG2_01_|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|P|4|1 _PG2_01_|P|A4 _PG2_01_|P|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|P|4|P _PG2_01_|P|4|MID_SERIES 0  2e-13
R_PG2_01_|P|4|B _PG2_01_|P|A4 _PG2_01_|P|4|MID_SHUNT  2.7439617672
L_PG2_01_|P|4|RB _PG2_01_|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|P|T|1 _PG2_01_|P|T1 _PG2_01_|P|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|P|T|P _PG2_01_|P|T|MID_SERIES 0  2e-13
R_PG2_01_|P|T|B _PG2_01_|P|T1 _PG2_01_|P|T|MID_SHUNT  2.7439617672
L_PG2_01_|P|T|RB _PG2_01_|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|P|45|1 _PG2_01_|P|T2 _PG2_01_|P|A4 JJMIT AREA=1.7857142857142858
R_PG2_01_|P|45|B _PG2_01_|P|T2 _PG2_01_|P|45|MID_SHUNT  3.84154647408
L_PG2_01_|P|45|RB _PG2_01_|P|45|MID_SHUNT _PG2_01_|P|A4  2.1704737578552e-12
B_PG2_01_|P|6|1 _PG2_01_|P|Q1 _PG2_01_|P|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|P|6|P _PG2_01_|P|6|MID_SERIES 0  2e-13
R_PG2_01_|P|6|B _PG2_01_|P|Q1 _PG2_01_|P|6|MID_SHUNT  2.7439617672
L_PG2_01_|P|6|RB _PG2_01_|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_01_|G|I_1|B _PG2_01_|G|A1 _PG2_01_|G|I_1|MID  2e-12
I_PG2_01_|G|I_1|B 0 _PG2_01_|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01_|G|I_3|B _PG2_01_|G|A3 _PG2_01_|G|I_3|MID  2e-12
I_PG2_01_|G|I_3|B 0 _PG2_01_|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01_|G|I_T|B _PG2_01_|G|T1 _PG2_01_|G|I_T|MID  2e-12
I_PG2_01_|G|I_T|B 0 _PG2_01_|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01_|G|I_6|B _PG2_01_|G|Q1 _PG2_01_|G|I_6|MID  2e-12
I_PG2_01_|G|I_6|B 0 _PG2_01_|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01_|G|1|1 _PG2_01_|G|A1 _PG2_01_|G|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|G|1|P _PG2_01_|G|1|MID_SERIES 0  2e-13
R_PG2_01_|G|1|B _PG2_01_|G|A1 _PG2_01_|G|1|MID_SHUNT  2.7439617672
L_PG2_01_|G|1|RB _PG2_01_|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|G|23|1 _PG2_01_|G|A2 _PG2_01_|G|A3 JJMIT AREA=1.7857142857142858
R_PG2_01_|G|23|B _PG2_01_|G|A2 _PG2_01_|G|23|MID_SHUNT  3.84154647408
L_PG2_01_|G|23|RB _PG2_01_|G|23|MID_SHUNT _PG2_01_|G|A3  2.1704737578552e-12
B_PG2_01_|G|3|1 _PG2_01_|G|A3 _PG2_01_|G|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|G|3|P _PG2_01_|G|3|MID_SERIES 0  2e-13
R_PG2_01_|G|3|B _PG2_01_|G|A3 _PG2_01_|G|3|MID_SHUNT  2.7439617672
L_PG2_01_|G|3|RB _PG2_01_|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|G|4|1 _PG2_01_|G|A4 _PG2_01_|G|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|G|4|P _PG2_01_|G|4|MID_SERIES 0  2e-13
R_PG2_01_|G|4|B _PG2_01_|G|A4 _PG2_01_|G|4|MID_SHUNT  2.7439617672
L_PG2_01_|G|4|RB _PG2_01_|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|G|T|1 _PG2_01_|G|T1 _PG2_01_|G|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|G|T|P _PG2_01_|G|T|MID_SERIES 0  2e-13
R_PG2_01_|G|T|B _PG2_01_|G|T1 _PG2_01_|G|T|MID_SHUNT  2.7439617672
L_PG2_01_|G|T|RB _PG2_01_|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01_|G|45|1 _PG2_01_|G|T2 _PG2_01_|G|A4 JJMIT AREA=1.7857142857142858
R_PG2_01_|G|45|B _PG2_01_|G|T2 _PG2_01_|G|45|MID_SHUNT  3.84154647408
L_PG2_01_|G|45|RB _PG2_01_|G|45|MID_SHUNT _PG2_01_|G|A4  2.1704737578552e-12
B_PG2_01_|G|6|1 _PG2_01_|G|Q1 _PG2_01_|G|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01_|G|6|P _PG2_01_|G|6|MID_SERIES 0  2e-13
R_PG2_01_|G|6|B _PG2_01_|G|Q1 _PG2_01_|G|6|MID_SHUNT  2.7439617672
L_PG2_01_|G|6|RB _PG2_01_|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_SPL_G1|I_D1|B _PG3_01_|_SPL_G1|D1 _PG3_01_|_SPL_G1|I_D1|MID  2e-12
I_PG3_01_|_SPL_G1|I_D1|B 0 _PG3_01_|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_SPL_G1|I_D2|B _PG3_01_|_SPL_G1|D2 _PG3_01_|_SPL_G1|I_D2|MID  2e-12
I_PG3_01_|_SPL_G1|I_D2|B 0 _PG3_01_|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PG3_01_|_SPL_G1|I_Q1|B _PG3_01_|_SPL_G1|QA1 _PG3_01_|_SPL_G1|I_Q1|MID  2e-12
I_PG3_01_|_SPL_G1|I_Q1|B 0 _PG3_01_|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_SPL_G1|I_Q2|B _PG3_01_|_SPL_G1|QB1 _PG3_01_|_SPL_G1|I_Q2|MID  2e-12
I_PG3_01_|_SPL_G1|I_Q2|B 0 _PG3_01_|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_SPL_G1|1|1 _PG3_01_|_SPL_G1|D1 _PG3_01_|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_G1|1|P _PG3_01_|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_G1|1|B _PG3_01_|_SPL_G1|D1 _PG3_01_|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_G1|1|RB _PG3_01_|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_SPL_G1|2|1 _PG3_01_|_SPL_G1|D2 _PG3_01_|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_G1|2|P _PG3_01_|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_G1|2|B _PG3_01_|_SPL_G1|D2 _PG3_01_|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_G1|2|RB _PG3_01_|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_SPL_G1|A|1 _PG3_01_|_SPL_G1|QA1 _PG3_01_|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_G1|A|P _PG3_01_|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_G1|A|B _PG3_01_|_SPL_G1|QA1 _PG3_01_|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_G1|A|RB _PG3_01_|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_SPL_G1|B|1 _PG3_01_|_SPL_G1|QB1 _PG3_01_|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_G1|B|P _PG3_01_|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_G1|B|B _PG3_01_|_SPL_G1|QB1 _PG3_01_|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_G1|B|RB _PG3_01_|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_SPL_P1|I_D1|B _PG3_01_|_SPL_P1|D1 _PG3_01_|_SPL_P1|I_D1|MID  2e-12
I_PG3_01_|_SPL_P1|I_D1|B 0 _PG3_01_|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_SPL_P1|I_D2|B _PG3_01_|_SPL_P1|D2 _PG3_01_|_SPL_P1|I_D2|MID  2e-12
I_PG3_01_|_SPL_P1|I_D2|B 0 _PG3_01_|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PG3_01_|_SPL_P1|I_Q1|B _PG3_01_|_SPL_P1|QA1 _PG3_01_|_SPL_P1|I_Q1|MID  2e-12
I_PG3_01_|_SPL_P1|I_Q1|B 0 _PG3_01_|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_SPL_P1|I_Q2|B _PG3_01_|_SPL_P1|QB1 _PG3_01_|_SPL_P1|I_Q2|MID  2e-12
I_PG3_01_|_SPL_P1|I_Q2|B 0 _PG3_01_|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_SPL_P1|1|1 _PG3_01_|_SPL_P1|D1 _PG3_01_|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_P1|1|P _PG3_01_|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_P1|1|B _PG3_01_|_SPL_P1|D1 _PG3_01_|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_P1|1|RB _PG3_01_|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_SPL_P1|2|1 _PG3_01_|_SPL_P1|D2 _PG3_01_|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_P1|2|P _PG3_01_|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_P1|2|B _PG3_01_|_SPL_P1|D2 _PG3_01_|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_P1|2|RB _PG3_01_|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_SPL_P1|A|1 _PG3_01_|_SPL_P1|QA1 _PG3_01_|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_P1|A|P _PG3_01_|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_P1|A|B _PG3_01_|_SPL_P1|QA1 _PG3_01_|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_P1|A|RB _PG3_01_|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_SPL_P1|B|1 _PG3_01_|_SPL_P1|QB1 _PG3_01_|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_SPL_P1|B|P _PG3_01_|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_01_|_SPL_P1|B|B _PG3_01_|_SPL_P1|QB1 _PG3_01_|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_01_|_SPL_P1|B|RB _PG3_01_|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_PG|I_A1|B _PG3_01_|_PG|A1 _PG3_01_|_PG|I_A1|MID  2e-12
I_PG3_01_|_PG|I_A1|B 0 _PG3_01_|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_PG|I_B1|B _PG3_01_|_PG|B1 _PG3_01_|_PG|I_B1|MID  2e-12
I_PG3_01_|_PG|I_B1|B 0 _PG3_01_|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_PG|I_Q3|B _PG3_01_|_PG|Q3 _PG3_01_|_PG|I_Q3|MID  2e-12
I_PG3_01_|_PG|I_Q3|B 0 _PG3_01_|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01_|_PG|I_Q2|B _PG3_01_|_PG|Q2 _PG3_01_|_PG|I_Q2|MID  2e-12
I_PG3_01_|_PG|I_Q2|B 0 _PG3_01_|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_PG|I_Q1|B _PG3_01_|_PG|Q1 _PG3_01_|_PG|I_Q1|MID  2e-12
I_PG3_01_|_PG|I_Q1|B 0 _PG3_01_|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_PG|A1|1 _PG3_01_|_PG|A1 _PG3_01_|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_PG|A1|P _PG3_01_|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01_|_PG|A1|B _PG3_01_|_PG|A1 _PG3_01_|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01_|_PG|A1|RB _PG3_01_|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_PG|A2|1 _PG3_01_|_PG|A2 _PG3_01_|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_PG|A2|P _PG3_01_|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01_|_PG|A2|B _PG3_01_|_PG|A2 _PG3_01_|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01_|_PG|A2|RB _PG3_01_|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_PG|A12|1 _PG3_01_|_PG|A2 _PG3_01_|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_PG|A12|B _PG3_01_|_PG|A2 _PG3_01_|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01_|_PG|A12|RB _PG3_01_|_PG|A12|MID_SHUNT _PG3_01_|_PG|A3  2.1704737578552e-12
B_PG3_01_|_PG|B1|1 _PG3_01_|_PG|B1 _PG3_01_|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_PG|B1|P _PG3_01_|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01_|_PG|B1|B _PG3_01_|_PG|B1 _PG3_01_|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01_|_PG|B1|RB _PG3_01_|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_PG|B2|1 _PG3_01_|_PG|B2 _PG3_01_|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_PG|B2|P _PG3_01_|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01_|_PG|B2|B _PG3_01_|_PG|B2 _PG3_01_|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01_|_PG|B2|RB _PG3_01_|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_PG|B12|1 _PG3_01_|_PG|B2 _PG3_01_|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_PG|B12|B _PG3_01_|_PG|B2 _PG3_01_|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01_|_PG|B12|RB _PG3_01_|_PG|B12|MID_SHUNT _PG3_01_|_PG|B3  2.1704737578552e-12
B_PG3_01_|_PG|Q2|1 _PG3_01_|_PG|Q2 _PG3_01_|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_PG|Q2|P _PG3_01_|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01_|_PG|Q2|B _PG3_01_|_PG|Q2 _PG3_01_|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01_|_PG|Q2|RB _PG3_01_|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_PG|Q1|1 _PG3_01_|_PG|Q1 _PG3_01_|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_PG|Q1|P _PG3_01_|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01_|_PG|Q1|B _PG3_01_|_PG|Q1 _PG3_01_|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01_|_PG|Q1|RB _PG3_01_|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_GG|I_A1|B _PG3_01_|_GG|A1 _PG3_01_|_GG|I_A1|MID  2e-12
I_PG3_01_|_GG|I_A1|B 0 _PG3_01_|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_GG|I_B1|B _PG3_01_|_GG|B1 _PG3_01_|_GG|I_B1|MID  2e-12
I_PG3_01_|_GG|I_B1|B 0 _PG3_01_|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_GG|I_Q3|B _PG3_01_|_GG|Q3 _PG3_01_|_GG|I_Q3|MID  2e-12
I_PG3_01_|_GG|I_Q3|B 0 _PG3_01_|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01_|_GG|I_Q2|B _PG3_01_|_GG|Q2 _PG3_01_|_GG|I_Q2|MID  2e-12
I_PG3_01_|_GG|I_Q2|B 0 _PG3_01_|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_GG|I_Q1|B _PG3_01_|_GG|Q1 _PG3_01_|_GG|I_Q1|MID  2e-12
I_PG3_01_|_GG|I_Q1|B 0 _PG3_01_|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_GG|A1|1 _PG3_01_|_GG|A1 _PG3_01_|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_GG|A1|P _PG3_01_|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01_|_GG|A1|B _PG3_01_|_GG|A1 _PG3_01_|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01_|_GG|A1|RB _PG3_01_|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_GG|A2|1 _PG3_01_|_GG|A2 _PG3_01_|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_GG|A2|P _PG3_01_|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01_|_GG|A2|B _PG3_01_|_GG|A2 _PG3_01_|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01_|_GG|A2|RB _PG3_01_|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_GG|A12|1 _PG3_01_|_GG|A2 _PG3_01_|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_GG|A12|B _PG3_01_|_GG|A2 _PG3_01_|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01_|_GG|A12|RB _PG3_01_|_GG|A12|MID_SHUNT _PG3_01_|_GG|A3  2.1704737578552e-12
B_PG3_01_|_GG|B1|1 _PG3_01_|_GG|B1 _PG3_01_|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_GG|B1|P _PG3_01_|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01_|_GG|B1|B _PG3_01_|_GG|B1 _PG3_01_|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01_|_GG|B1|RB _PG3_01_|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_GG|B2|1 _PG3_01_|_GG|B2 _PG3_01_|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_GG|B2|P _PG3_01_|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01_|_GG|B2|B _PG3_01_|_GG|B2 _PG3_01_|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01_|_GG|B2|RB _PG3_01_|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_GG|B12|1 _PG3_01_|_GG|B2 _PG3_01_|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_GG|B12|B _PG3_01_|_GG|B2 _PG3_01_|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01_|_GG|B12|RB _PG3_01_|_GG|B12|MID_SHUNT _PG3_01_|_GG|B3  2.1704737578552e-12
B_PG3_01_|_GG|Q2|1 _PG3_01_|_GG|Q2 _PG3_01_|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_GG|Q2|P _PG3_01_|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01_|_GG|Q2|B _PG3_01_|_GG|Q2 _PG3_01_|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01_|_GG|Q2|RB _PG3_01_|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_GG|Q1|1 _PG3_01_|_GG|Q1 _PG3_01_|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_GG|Q1|P _PG3_01_|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01_|_GG|Q1|B _PG3_01_|_GG|Q1 _PG3_01_|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01_|_GG|Q1|RB _PG3_01_|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_DFF_P0|I_1|B _PG3_01_|_DFF_P0|A1 _PG3_01_|_DFF_P0|I_1|MID  2e-12
I_PG3_01_|_DFF_P0|I_1|B 0 _PG3_01_|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_P0|I_3|B _PG3_01_|_DFF_P0|A3 _PG3_01_|_DFF_P0|I_3|MID  2e-12
I_PG3_01_|_DFF_P0|I_3|B 0 _PG3_01_|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01_|_DFF_P0|I_T|B _PG3_01_|_DFF_P0|T1 _PG3_01_|_DFF_P0|I_T|MID  2e-12
I_PG3_01_|_DFF_P0|I_T|B 0 _PG3_01_|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_P0|I_6|B _PG3_01_|_DFF_P0|Q1 _PG3_01_|_DFF_P0|I_6|MID  2e-12
I_PG3_01_|_DFF_P0|I_6|B 0 _PG3_01_|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_DFF_P0|1|1 _PG3_01_|_DFF_P0|A1 _PG3_01_|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P0|1|P _PG3_01_|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P0|1|B _PG3_01_|_DFF_P0|A1 _PG3_01_|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P0|1|RB _PG3_01_|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P0|23|1 _PG3_01_|_DFF_P0|A2 _PG3_01_|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_P0|23|B _PG3_01_|_DFF_P0|A2 _PG3_01_|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_P0|23|RB _PG3_01_|_DFF_P0|23|MID_SHUNT _PG3_01_|_DFF_P0|A3  2.1704737578552e-12
B_PG3_01_|_DFF_P0|3|1 _PG3_01_|_DFF_P0|A3 _PG3_01_|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P0|3|P _PG3_01_|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P0|3|B _PG3_01_|_DFF_P0|A3 _PG3_01_|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P0|3|RB _PG3_01_|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P0|4|1 _PG3_01_|_DFF_P0|A4 _PG3_01_|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P0|4|P _PG3_01_|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P0|4|B _PG3_01_|_DFF_P0|A4 _PG3_01_|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P0|4|RB _PG3_01_|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P0|T|1 _PG3_01_|_DFF_P0|T1 _PG3_01_|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P0|T|P _PG3_01_|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P0|T|B _PG3_01_|_DFF_P0|T1 _PG3_01_|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P0|T|RB _PG3_01_|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P0|45|1 _PG3_01_|_DFF_P0|T2 _PG3_01_|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_P0|45|B _PG3_01_|_DFF_P0|T2 _PG3_01_|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_P0|45|RB _PG3_01_|_DFF_P0|45|MID_SHUNT _PG3_01_|_DFF_P0|A4  2.1704737578552e-12
B_PG3_01_|_DFF_P0|6|1 _PG3_01_|_DFF_P0|Q1 _PG3_01_|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P0|6|P _PG3_01_|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P0|6|B _PG3_01_|_DFF_P0|Q1 _PG3_01_|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P0|6|RB _PG3_01_|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_DFF_P1|I_1|B _PG3_01_|_DFF_P1|A1 _PG3_01_|_DFF_P1|I_1|MID  2e-12
I_PG3_01_|_DFF_P1|I_1|B 0 _PG3_01_|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_P1|I_3|B _PG3_01_|_DFF_P1|A3 _PG3_01_|_DFF_P1|I_3|MID  2e-12
I_PG3_01_|_DFF_P1|I_3|B 0 _PG3_01_|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01_|_DFF_P1|I_T|B _PG3_01_|_DFF_P1|T1 _PG3_01_|_DFF_P1|I_T|MID  2e-12
I_PG3_01_|_DFF_P1|I_T|B 0 _PG3_01_|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_P1|I_6|B _PG3_01_|_DFF_P1|Q1 _PG3_01_|_DFF_P1|I_6|MID  2e-12
I_PG3_01_|_DFF_P1|I_6|B 0 _PG3_01_|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_DFF_P1|1|1 _PG3_01_|_DFF_P1|A1 _PG3_01_|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P1|1|P _PG3_01_|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P1|1|B _PG3_01_|_DFF_P1|A1 _PG3_01_|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P1|1|RB _PG3_01_|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P1|23|1 _PG3_01_|_DFF_P1|A2 _PG3_01_|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_P1|23|B _PG3_01_|_DFF_P1|A2 _PG3_01_|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_P1|23|RB _PG3_01_|_DFF_P1|23|MID_SHUNT _PG3_01_|_DFF_P1|A3  2.1704737578552e-12
B_PG3_01_|_DFF_P1|3|1 _PG3_01_|_DFF_P1|A3 _PG3_01_|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P1|3|P _PG3_01_|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P1|3|B _PG3_01_|_DFF_P1|A3 _PG3_01_|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P1|3|RB _PG3_01_|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P1|4|1 _PG3_01_|_DFF_P1|A4 _PG3_01_|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P1|4|P _PG3_01_|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P1|4|B _PG3_01_|_DFF_P1|A4 _PG3_01_|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P1|4|RB _PG3_01_|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P1|T|1 _PG3_01_|_DFF_P1|T1 _PG3_01_|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P1|T|P _PG3_01_|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P1|T|B _PG3_01_|_DFF_P1|T1 _PG3_01_|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P1|T|RB _PG3_01_|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_P1|45|1 _PG3_01_|_DFF_P1|T2 _PG3_01_|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_P1|45|B _PG3_01_|_DFF_P1|T2 _PG3_01_|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_P1|45|RB _PG3_01_|_DFF_P1|45|MID_SHUNT _PG3_01_|_DFF_P1|A4  2.1704737578552e-12
B_PG3_01_|_DFF_P1|6|1 _PG3_01_|_DFF_P1|Q1 _PG3_01_|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_P1|6|P _PG3_01_|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_P1|6|B _PG3_01_|_DFF_P1|Q1 _PG3_01_|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_P1|6|RB _PG3_01_|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_DFF_PG|I_1|B _PG3_01_|_DFF_PG|A1 _PG3_01_|_DFF_PG|I_1|MID  2e-12
I_PG3_01_|_DFF_PG|I_1|B 0 _PG3_01_|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_PG|I_3|B _PG3_01_|_DFF_PG|A3 _PG3_01_|_DFF_PG|I_3|MID  2e-12
I_PG3_01_|_DFF_PG|I_3|B 0 _PG3_01_|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01_|_DFF_PG|I_T|B _PG3_01_|_DFF_PG|T1 _PG3_01_|_DFF_PG|I_T|MID  2e-12
I_PG3_01_|_DFF_PG|I_T|B 0 _PG3_01_|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_PG|I_6|B _PG3_01_|_DFF_PG|Q1 _PG3_01_|_DFF_PG|I_6|MID  2e-12
I_PG3_01_|_DFF_PG|I_6|B 0 _PG3_01_|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_DFF_PG|1|1 _PG3_01_|_DFF_PG|A1 _PG3_01_|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_PG|1|P _PG3_01_|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_PG|1|B _PG3_01_|_DFF_PG|A1 _PG3_01_|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_PG|1|RB _PG3_01_|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_PG|23|1 _PG3_01_|_DFF_PG|A2 _PG3_01_|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_PG|23|B _PG3_01_|_DFF_PG|A2 _PG3_01_|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_PG|23|RB _PG3_01_|_DFF_PG|23|MID_SHUNT _PG3_01_|_DFF_PG|A3  2.1704737578552e-12
B_PG3_01_|_DFF_PG|3|1 _PG3_01_|_DFF_PG|A3 _PG3_01_|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_PG|3|P _PG3_01_|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_PG|3|B _PG3_01_|_DFF_PG|A3 _PG3_01_|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_PG|3|RB _PG3_01_|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_PG|4|1 _PG3_01_|_DFF_PG|A4 _PG3_01_|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_PG|4|P _PG3_01_|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_PG|4|B _PG3_01_|_DFF_PG|A4 _PG3_01_|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_PG|4|RB _PG3_01_|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_PG|T|1 _PG3_01_|_DFF_PG|T1 _PG3_01_|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_PG|T|P _PG3_01_|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_PG|T|B _PG3_01_|_DFF_PG|T1 _PG3_01_|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_PG|T|RB _PG3_01_|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_PG|45|1 _PG3_01_|_DFF_PG|T2 _PG3_01_|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_PG|45|B _PG3_01_|_DFF_PG|T2 _PG3_01_|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_PG|45|RB _PG3_01_|_DFF_PG|45|MID_SHUNT _PG3_01_|_DFF_PG|A4  2.1704737578552e-12
B_PG3_01_|_DFF_PG|6|1 _PG3_01_|_DFF_PG|Q1 _PG3_01_|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_PG|6|P _PG3_01_|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_PG|6|B _PG3_01_|_DFF_PG|Q1 _PG3_01_|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_PG|6|RB _PG3_01_|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_DFF_GG|I_1|B _PG3_01_|_DFF_GG|A1 _PG3_01_|_DFF_GG|I_1|MID  2e-12
I_PG3_01_|_DFF_GG|I_1|B 0 _PG3_01_|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_GG|I_3|B _PG3_01_|_DFF_GG|A3 _PG3_01_|_DFF_GG|I_3|MID  2e-12
I_PG3_01_|_DFF_GG|I_3|B 0 _PG3_01_|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01_|_DFF_GG|I_T|B _PG3_01_|_DFF_GG|T1 _PG3_01_|_DFF_GG|I_T|MID  2e-12
I_PG3_01_|_DFF_GG|I_T|B 0 _PG3_01_|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_DFF_GG|I_6|B _PG3_01_|_DFF_GG|Q1 _PG3_01_|_DFF_GG|I_6|MID  2e-12
I_PG3_01_|_DFF_GG|I_6|B 0 _PG3_01_|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_DFF_GG|1|1 _PG3_01_|_DFF_GG|A1 _PG3_01_|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_GG|1|P _PG3_01_|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_GG|1|B _PG3_01_|_DFF_GG|A1 _PG3_01_|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_GG|1|RB _PG3_01_|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_GG|23|1 _PG3_01_|_DFF_GG|A2 _PG3_01_|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_GG|23|B _PG3_01_|_DFF_GG|A2 _PG3_01_|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_GG|23|RB _PG3_01_|_DFF_GG|23|MID_SHUNT _PG3_01_|_DFF_GG|A3  2.1704737578552e-12
B_PG3_01_|_DFF_GG|3|1 _PG3_01_|_DFF_GG|A3 _PG3_01_|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_GG|3|P _PG3_01_|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_GG|3|B _PG3_01_|_DFF_GG|A3 _PG3_01_|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_GG|3|RB _PG3_01_|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_GG|4|1 _PG3_01_|_DFF_GG|A4 _PG3_01_|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_GG|4|P _PG3_01_|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_GG|4|B _PG3_01_|_DFF_GG|A4 _PG3_01_|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_GG|4|RB _PG3_01_|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_GG|T|1 _PG3_01_|_DFF_GG|T1 _PG3_01_|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_GG|T|P _PG3_01_|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_GG|T|B _PG3_01_|_DFF_GG|T1 _PG3_01_|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_GG|T|RB _PG3_01_|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_DFF_GG|45|1 _PG3_01_|_DFF_GG|T2 _PG3_01_|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01_|_DFF_GG|45|B _PG3_01_|_DFF_GG|T2 _PG3_01_|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_01_|_DFF_GG|45|RB _PG3_01_|_DFF_GG|45|MID_SHUNT _PG3_01_|_DFF_GG|A4  2.1704737578552e-12
B_PG3_01_|_DFF_GG|6|1 _PG3_01_|_DFF_GG|Q1 _PG3_01_|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_DFF_GG|6|P _PG3_01_|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_01_|_DFF_GG|6|B _PG3_01_|_DFF_GG|Q1 _PG3_01_|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_01_|_DFF_GG|6|RB _PG3_01_|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_AND_G|I_A1|B _PG3_01_|_AND_G|A1 _PG3_01_|_AND_G|I_A1|MID  2e-12
I_PG3_01_|_AND_G|I_A1|B 0 _PG3_01_|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_AND_G|I_B1|B _PG3_01_|_AND_G|B1 _PG3_01_|_AND_G|I_B1|MID  2e-12
I_PG3_01_|_AND_G|I_B1|B 0 _PG3_01_|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_AND_G|I_Q3|B _PG3_01_|_AND_G|Q3 _PG3_01_|_AND_G|I_Q3|MID  2e-12
I_PG3_01_|_AND_G|I_Q3|B 0 _PG3_01_|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01_|_AND_G|I_Q2|B _PG3_01_|_AND_G|Q2 _PG3_01_|_AND_G|I_Q2|MID  2e-12
I_PG3_01_|_AND_G|I_Q2|B 0 _PG3_01_|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_AND_G|I_Q1|B _PG3_01_|_AND_G|Q1 _PG3_01_|_AND_G|I_Q1|MID  2e-12
I_PG3_01_|_AND_G|I_Q1|B 0 _PG3_01_|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_AND_G|A1|1 _PG3_01_|_AND_G|A1 _PG3_01_|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_G|A1|P _PG3_01_|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01_|_AND_G|A1|B _PG3_01_|_AND_G|A1 _PG3_01_|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_G|A1|RB _PG3_01_|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_G|A2|1 _PG3_01_|_AND_G|A2 _PG3_01_|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_G|A2|P _PG3_01_|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01_|_AND_G|A2|B _PG3_01_|_AND_G|A2 _PG3_01_|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_G|A2|RB _PG3_01_|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_G|A12|1 _PG3_01_|_AND_G|A2 _PG3_01_|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_AND_G|A12|B _PG3_01_|_AND_G|A2 _PG3_01_|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01_|_AND_G|A12|RB _PG3_01_|_AND_G|A12|MID_SHUNT _PG3_01_|_AND_G|A3  2.1704737578552e-12
B_PG3_01_|_AND_G|B1|1 _PG3_01_|_AND_G|B1 _PG3_01_|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_G|B1|P _PG3_01_|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01_|_AND_G|B1|B _PG3_01_|_AND_G|B1 _PG3_01_|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_G|B1|RB _PG3_01_|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_G|B2|1 _PG3_01_|_AND_G|B2 _PG3_01_|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_G|B2|P _PG3_01_|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01_|_AND_G|B2|B _PG3_01_|_AND_G|B2 _PG3_01_|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_G|B2|RB _PG3_01_|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_G|B12|1 _PG3_01_|_AND_G|B2 _PG3_01_|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_AND_G|B12|B _PG3_01_|_AND_G|B2 _PG3_01_|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01_|_AND_G|B12|RB _PG3_01_|_AND_G|B12|MID_SHUNT _PG3_01_|_AND_G|B3  2.1704737578552e-12
B_PG3_01_|_AND_G|Q2|1 _PG3_01_|_AND_G|Q2 _PG3_01_|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_G|Q2|P _PG3_01_|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01_|_AND_G|Q2|B _PG3_01_|_AND_G|Q2 _PG3_01_|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_G|Q2|RB _PG3_01_|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_G|Q1|1 _PG3_01_|_AND_G|Q1 _PG3_01_|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_G|Q1|P _PG3_01_|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01_|_AND_G|Q1|B _PG3_01_|_AND_G|Q1 _PG3_01_|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_G|Q1|RB _PG3_01_|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01_|_AND_P|I_A1|B _PG3_01_|_AND_P|A1 _PG3_01_|_AND_P|I_A1|MID  2e-12
I_PG3_01_|_AND_P|I_A1|B 0 _PG3_01_|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_AND_P|I_B1|B _PG3_01_|_AND_P|B1 _PG3_01_|_AND_P|I_B1|MID  2e-12
I_PG3_01_|_AND_P|I_B1|B 0 _PG3_01_|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_AND_P|I_Q3|B _PG3_01_|_AND_P|Q3 _PG3_01_|_AND_P|I_Q3|MID  2e-12
I_PG3_01_|_AND_P|I_Q3|B 0 _PG3_01_|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01_|_AND_P|I_Q2|B _PG3_01_|_AND_P|Q2 _PG3_01_|_AND_P|I_Q2|MID  2e-12
I_PG3_01_|_AND_P|I_Q2|B 0 _PG3_01_|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01_|_AND_P|I_Q1|B _PG3_01_|_AND_P|Q1 _PG3_01_|_AND_P|I_Q1|MID  2e-12
I_PG3_01_|_AND_P|I_Q1|B 0 _PG3_01_|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01_|_AND_P|A1|1 _PG3_01_|_AND_P|A1 _PG3_01_|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_P|A1|P _PG3_01_|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01_|_AND_P|A1|B _PG3_01_|_AND_P|A1 _PG3_01_|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_P|A1|RB _PG3_01_|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_P|A2|1 _PG3_01_|_AND_P|A2 _PG3_01_|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_P|A2|P _PG3_01_|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01_|_AND_P|A2|B _PG3_01_|_AND_P|A2 _PG3_01_|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_P|A2|RB _PG3_01_|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_P|A12|1 _PG3_01_|_AND_P|A2 _PG3_01_|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_AND_P|A12|B _PG3_01_|_AND_P|A2 _PG3_01_|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01_|_AND_P|A12|RB _PG3_01_|_AND_P|A12|MID_SHUNT _PG3_01_|_AND_P|A3  2.1704737578552e-12
B_PG3_01_|_AND_P|B1|1 _PG3_01_|_AND_P|B1 _PG3_01_|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_P|B1|P _PG3_01_|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01_|_AND_P|B1|B _PG3_01_|_AND_P|B1 _PG3_01_|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_P|B1|RB _PG3_01_|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_P|B2|1 _PG3_01_|_AND_P|B2 _PG3_01_|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_P|B2|P _PG3_01_|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01_|_AND_P|B2|B _PG3_01_|_AND_P|B2 _PG3_01_|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_P|B2|RB _PG3_01_|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_P|B12|1 _PG3_01_|_AND_P|B2 _PG3_01_|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01_|_AND_P|B12|B _PG3_01_|_AND_P|B2 _PG3_01_|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01_|_AND_P|B12|RB _PG3_01_|_AND_P|B12|MID_SHUNT _PG3_01_|_AND_P|B3  2.1704737578552e-12
B_PG3_01_|_AND_P|Q2|1 _PG3_01_|_AND_P|Q2 _PG3_01_|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_P|Q2|P _PG3_01_|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01_|_AND_P|Q2|B _PG3_01_|_AND_P|Q2 _PG3_01_|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_P|Q2|RB _PG3_01_|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01_|_AND_P|Q1|1 _PG3_01_|_AND_P|Q1 _PG3_01_|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01_|_AND_P|Q1|P _PG3_01_|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01_|_AND_P|Q1|B _PG3_01_|_AND_P|Q1 _PG3_01_|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01_|_AND_P|Q1|RB _PG3_01_|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1_|SPL1|I_D1|B SPL_G1_1_|SPL1|D1 SPL_G1_1_|SPL1|I_D1|MID  2e-12
ISPL_G1_1_|SPL1|I_D1|B 0 SPL_G1_1_|SPL1|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1_|SPL1|I_D2|B SPL_G1_1_|SPL1|D2 SPL_G1_1_|SPL1|I_D2|MID  2e-12
ISPL_G1_1_|SPL1|I_D2|B 0 SPL_G1_1_|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_G1_1_|SPL1|I_Q1|B SPL_G1_1_|SPL1|QA1 SPL_G1_1_|SPL1|I_Q1|MID  2e-12
ISPL_G1_1_|SPL1|I_Q1|B 0 SPL_G1_1_|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1_|SPL1|I_Q2|B SPL_G1_1_|SPL1|QB1 SPL_G1_1_|SPL1|I_Q2|MID  2e-12
ISPL_G1_1_|SPL1|I_Q2|B 0 SPL_G1_1_|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_G1_1_|SPL1|1|1 SPL_G1_1_|SPL1|D1 SPL_G1_1_|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL1|1|P SPL_G1_1_|SPL1|1|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL1|1|B SPL_G1_1_|SPL1|D1 SPL_G1_1_|SPL1|1|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL1|1|RB SPL_G1_1_|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1_|SPL1|2|1 SPL_G1_1_|SPL1|D2 SPL_G1_1_|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL1|2|P SPL_G1_1_|SPL1|2|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL1|2|B SPL_G1_1_|SPL1|D2 SPL_G1_1_|SPL1|2|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL1|2|RB SPL_G1_1_|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1_|SPL1|A|1 SPL_G1_1_|SPL1|QA1 SPL_G1_1_|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL1|A|P SPL_G1_1_|SPL1|A|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL1|A|B SPL_G1_1_|SPL1|QA1 SPL_G1_1_|SPL1|A|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL1|A|RB SPL_G1_1_|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1_|SPL1|B|1 SPL_G1_1_|SPL1|QB1 SPL_G1_1_|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL1|B|P SPL_G1_1_|SPL1|B|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL1|B|B SPL_G1_1_|SPL1|QB1 SPL_G1_1_|SPL1|B|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL1|B|RB SPL_G1_1_|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1_|SPL2|I_D1|B SPL_G1_1_|SPL2|D1 SPL_G1_1_|SPL2|I_D1|MID  2e-12
ISPL_G1_1_|SPL2|I_D1|B 0 SPL_G1_1_|SPL2|I_D1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1_|SPL2|I_D2|B SPL_G1_1_|SPL2|D2 SPL_G1_1_|SPL2|I_D2|MID  2e-12
ISPL_G1_1_|SPL2|I_D2|B 0 SPL_G1_1_|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000245)
LSPL_G1_1_|SPL2|I_Q1|B SPL_G1_1_|SPL2|QA1 SPL_G1_1_|SPL2|I_Q1|MID  2e-12
ISPL_G1_1_|SPL2|I_Q1|B 0 SPL_G1_1_|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
LSPL_G1_1_|SPL2|I_Q2|B SPL_G1_1_|SPL2|QB1 SPL_G1_1_|SPL2|I_Q2|MID  2e-12
ISPL_G1_1_|SPL2|I_Q2|B 0 SPL_G1_1_|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
BSPL_G1_1_|SPL2|1|1 SPL_G1_1_|SPL2|D1 SPL_G1_1_|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL2|1|P SPL_G1_1_|SPL2|1|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL2|1|B SPL_G1_1_|SPL2|D1 SPL_G1_1_|SPL2|1|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL2|1|RB SPL_G1_1_|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1_|SPL2|2|1 SPL_G1_1_|SPL2|D2 SPL_G1_1_|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL2|2|P SPL_G1_1_|SPL2|2|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL2|2|B SPL_G1_1_|SPL2|D2 SPL_G1_1_|SPL2|2|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL2|2|RB SPL_G1_1_|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1_|SPL2|A|1 SPL_G1_1_|SPL2|QA1 SPL_G1_1_|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL2|A|P SPL_G1_1_|SPL2|A|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL2|A|B SPL_G1_1_|SPL2|QA1 SPL_G1_1_|SPL2|A|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL2|A|RB SPL_G1_1_|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1_|SPL2|B|1 SPL_G1_1_|SPL2|QB1 SPL_G1_1_|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1_|SPL2|B|P SPL_G1_1_|SPL2|B|MID_SERIES 0  2e-13
RSPL_G1_1_|SPL2|B|B SPL_G1_1_|SPL2|QB1 SPL_G1_1_|SPL2|B|MID_SHUNT  2.7439617672
LSPL_G1_1_|SPL2|B|RB SPL_G1_1_|SPL2|B|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_P0_1
.print DEVI R_G0_1
.print DEVI R_P1_1_TO1
.print DEVI R_P1_1_TO2
.print DEVI R_P1_1_TO3
.print DEVI R_G1_1_TO1
.print DEVI R_G1_1_TO2
.print DEVI R_G1_1_TO3
.print DEVI R_P2_1
.print DEVI R_G2_1
.print DEVI R_P3_1
.print DEVI R_G3_1
.print DEVI R_IP1_1
.print DEVI R_IP2_1
.print DEVI R_IP3_1
.print DEVI IA0_|A
.print DEVI IB0_|B
.print DEVI IA1_|C
.print DEVI IB1_|D
.print DEVI IA2_|E
.print DEVI IB2_|F
.print DEVI IA3_|G
.print DEVI IB3_|H
.print DEVI IT00_|T
.print DEVI IT01_|T
.print DEVI IT02_|T
.print DEVI IT03_|T
.print DEVI LSPL_IG0_0_|1
.print DEVI LSPL_IG0_0_|2
.print DEVI LSPL_IG0_0_|3
.print DEVI LSPL_IG0_0_|4
.print DEVI LSPL_IG0_0_|5
.print DEVI LSPL_IG0_0_|6
.print DEVI LSPL_IG0_0_|7
.print DEVI LSPL_IP1_0_|1
.print DEVI LSPL_IP1_0_|2
.print DEVI LSPL_IP1_0_|3
.print DEVI LSPL_IP1_0_|4
.print DEVI LSPL_IP1_0_|5
.print DEVI LSPL_IP1_0_|6
.print DEVI LSPL_IP1_0_|7
.print DEVI LSPL_IG2_0_|1
.print DEVI LSPL_IG2_0_|2
.print DEVI LSPL_IG2_0_|3
.print DEVI LSPL_IG2_0_|4
.print DEVI LSPL_IG2_0_|5
.print DEVI LSPL_IG2_0_|6
.print DEVI LSPL_IG2_0_|7
.print DEVI LSPL_IP3_0_|1
.print DEVI LSPL_IP3_0_|2
.print DEVI LSPL_IP3_0_|3
.print DEVI LSPL_IP3_0_|4
.print DEVI LSPL_IP3_0_|5
.print DEVI LSPL_IP3_0_|6
.print DEVI LSPL_IP3_0_|7
.print DEVI IT04_|T
.print DEVI IT05_|T
.print DEVI IT06_|T
.print DEVI IT07_|T
.print DEVI ID01_|T
.print DEVI L_DFF_IP1_01_|1
.print DEVI L_DFF_IP1_01_|2
.print DEVI L_DFF_IP1_01_|3
.print DEVI L_DFF_IP1_01_|T
.print DEVI L_DFF_IP1_01_|4
.print DEVI L_DFF_IP1_01_|5
.print DEVI L_DFF_IP1_01_|6
.print DEVI ID02_|T
.print DEVI L_DFF_IP2_01_|1
.print DEVI L_DFF_IP2_01_|2
.print DEVI L_DFF_IP2_01_|3
.print DEVI L_DFF_IP2_01_|T
.print DEVI L_DFF_IP2_01_|4
.print DEVI L_DFF_IP2_01_|5
.print DEVI L_DFF_IP2_01_|6
.print DEVI ID03_|T
.print DEVI L_DFF_IP3_01_|1
.print DEVI L_DFF_IP3_01_|2
.print DEVI L_DFF_IP3_01_|3
.print DEVI L_DFF_IP3_01_|T
.print DEVI L_DFF_IP3_01_|4
.print DEVI L_DFF_IP3_01_|5
.print DEVI L_DFF_IP3_01_|6
.print DEVI LI0_|_SPL_A|1
.print DEVI LI0_|_SPL_A|2
.print DEVI LI0_|_SPL_A|3
.print DEVI LI0_|_SPL_A|4
.print DEVI LI0_|_SPL_A|5
.print DEVI LI0_|_SPL_A|6
.print DEVI LI0_|_SPL_A|7
.print DEVI LI0_|_SPL_B|1
.print DEVI LI0_|_SPL_B|2
.print DEVI LI0_|_SPL_B|3
.print DEVI LI0_|_SPL_B|4
.print DEVI LI0_|_SPL_B|5
.print DEVI LI0_|_SPL_B|6
.print DEVI LI0_|_SPL_B|7
.print DEVI LI0_|_DFF_A|1
.print DEVI LI0_|_DFF_A|2
.print DEVI LI0_|_DFF_A|3
.print DEVI LI0_|_DFF_A|T
.print DEVI LI0_|_DFF_A|4
.print DEVI LI0_|_DFF_A|5
.print DEVI LI0_|_DFF_A|6
.print DEVI LI0_|_DFF_B|1
.print DEVI LI0_|_DFF_B|2
.print DEVI LI0_|_DFF_B|3
.print DEVI LI0_|_DFF_B|T
.print DEVI LI0_|_DFF_B|4
.print DEVI LI0_|_DFF_B|5
.print DEVI LI0_|_DFF_B|6
.print DEVI LI0_|_XOR|A1
.print DEVI LI0_|_XOR|A2
.print DEVI LI0_|_XOR|A3
.print DEVI LI0_|_XOR|B1
.print DEVI LI0_|_XOR|B2
.print DEVI LI0_|_XOR|B3
.print DEVI LI0_|_XOR|T1
.print DEVI LI0_|_XOR|T2
.print DEVI LI0_|_XOR|Q2
.print DEVI LI0_|_XOR|Q1
.print DEVI LI0_|_AND|A1
.print DEVI LI0_|_AND|A2
.print DEVI LI0_|_AND|A3
.print DEVI LI0_|_AND|B1
.print DEVI LI0_|_AND|B2
.print DEVI LI0_|_AND|B3
.print DEVI LI0_|_AND|Q3
.print DEVI LI0_|_AND|Q2
.print DEVI LI0_|_AND|Q1
.print DEVI LI1_|_SPL_A|1
.print DEVI LI1_|_SPL_A|2
.print DEVI LI1_|_SPL_A|3
.print DEVI LI1_|_SPL_A|4
.print DEVI LI1_|_SPL_A|5
.print DEVI LI1_|_SPL_A|6
.print DEVI LI1_|_SPL_A|7
.print DEVI LI1_|_SPL_B|1
.print DEVI LI1_|_SPL_B|2
.print DEVI LI1_|_SPL_B|3
.print DEVI LI1_|_SPL_B|4
.print DEVI LI1_|_SPL_B|5
.print DEVI LI1_|_SPL_B|6
.print DEVI LI1_|_SPL_B|7
.print DEVI LI1_|_DFF_A|1
.print DEVI LI1_|_DFF_A|2
.print DEVI LI1_|_DFF_A|3
.print DEVI LI1_|_DFF_A|T
.print DEVI LI1_|_DFF_A|4
.print DEVI LI1_|_DFF_A|5
.print DEVI LI1_|_DFF_A|6
.print DEVI LI1_|_DFF_B|1
.print DEVI LI1_|_DFF_B|2
.print DEVI LI1_|_DFF_B|3
.print DEVI LI1_|_DFF_B|T
.print DEVI LI1_|_DFF_B|4
.print DEVI LI1_|_DFF_B|5
.print DEVI LI1_|_DFF_B|6
.print DEVI LI1_|_XOR|A1
.print DEVI LI1_|_XOR|A2
.print DEVI LI1_|_XOR|A3
.print DEVI LI1_|_XOR|B1
.print DEVI LI1_|_XOR|B2
.print DEVI LI1_|_XOR|B3
.print DEVI LI1_|_XOR|T1
.print DEVI LI1_|_XOR|T2
.print DEVI LI1_|_XOR|Q2
.print DEVI LI1_|_XOR|Q1
.print DEVI LI1_|_AND|A1
.print DEVI LI1_|_AND|A2
.print DEVI LI1_|_AND|A3
.print DEVI LI1_|_AND|B1
.print DEVI LI1_|_AND|B2
.print DEVI LI1_|_AND|B3
.print DEVI LI1_|_AND|Q3
.print DEVI LI1_|_AND|Q2
.print DEVI LI1_|_AND|Q1
.print DEVI LI2_|_SPL_A|1
.print DEVI LI2_|_SPL_A|2
.print DEVI LI2_|_SPL_A|3
.print DEVI LI2_|_SPL_A|4
.print DEVI LI2_|_SPL_A|5
.print DEVI LI2_|_SPL_A|6
.print DEVI LI2_|_SPL_A|7
.print DEVI LI2_|_SPL_B|1
.print DEVI LI2_|_SPL_B|2
.print DEVI LI2_|_SPL_B|3
.print DEVI LI2_|_SPL_B|4
.print DEVI LI2_|_SPL_B|5
.print DEVI LI2_|_SPL_B|6
.print DEVI LI2_|_SPL_B|7
.print DEVI LI2_|_DFF_A|1
.print DEVI LI2_|_DFF_A|2
.print DEVI LI2_|_DFF_A|3
.print DEVI LI2_|_DFF_A|T
.print DEVI LI2_|_DFF_A|4
.print DEVI LI2_|_DFF_A|5
.print DEVI LI2_|_DFF_A|6
.print DEVI LI2_|_DFF_B|1
.print DEVI LI2_|_DFF_B|2
.print DEVI LI2_|_DFF_B|3
.print DEVI LI2_|_DFF_B|T
.print DEVI LI2_|_DFF_B|4
.print DEVI LI2_|_DFF_B|5
.print DEVI LI2_|_DFF_B|6
.print DEVI LI2_|_XOR|A1
.print DEVI LI2_|_XOR|A2
.print DEVI LI2_|_XOR|A3
.print DEVI LI2_|_XOR|B1
.print DEVI LI2_|_XOR|B2
.print DEVI LI2_|_XOR|B3
.print DEVI LI2_|_XOR|T1
.print DEVI LI2_|_XOR|T2
.print DEVI LI2_|_XOR|Q2
.print DEVI LI2_|_XOR|Q1
.print DEVI LI2_|_AND|A1
.print DEVI LI2_|_AND|A2
.print DEVI LI2_|_AND|A3
.print DEVI LI2_|_AND|B1
.print DEVI LI2_|_AND|B2
.print DEVI LI2_|_AND|B3
.print DEVI LI2_|_AND|Q3
.print DEVI LI2_|_AND|Q2
.print DEVI LI2_|_AND|Q1
.print DEVI LI3_|_SPL_A|1
.print DEVI LI3_|_SPL_A|2
.print DEVI LI3_|_SPL_A|3
.print DEVI LI3_|_SPL_A|4
.print DEVI LI3_|_SPL_A|5
.print DEVI LI3_|_SPL_A|6
.print DEVI LI3_|_SPL_A|7
.print DEVI LI3_|_SPL_B|1
.print DEVI LI3_|_SPL_B|2
.print DEVI LI3_|_SPL_B|3
.print DEVI LI3_|_SPL_B|4
.print DEVI LI3_|_SPL_B|5
.print DEVI LI3_|_SPL_B|6
.print DEVI LI3_|_SPL_B|7
.print DEVI LI3_|_DFF_A|1
.print DEVI LI3_|_DFF_A|2
.print DEVI LI3_|_DFF_A|3
.print DEVI LI3_|_DFF_A|T
.print DEVI LI3_|_DFF_A|4
.print DEVI LI3_|_DFF_A|5
.print DEVI LI3_|_DFF_A|6
.print DEVI LI3_|_DFF_B|1
.print DEVI LI3_|_DFF_B|2
.print DEVI LI3_|_DFF_B|3
.print DEVI LI3_|_DFF_B|T
.print DEVI LI3_|_DFF_B|4
.print DEVI LI3_|_DFF_B|5
.print DEVI LI3_|_DFF_B|6
.print DEVI LI3_|_XOR|A1
.print DEVI LI3_|_XOR|A2
.print DEVI LI3_|_XOR|A3
.print DEVI LI3_|_XOR|B1
.print DEVI LI3_|_XOR|B2
.print DEVI LI3_|_XOR|B3
.print DEVI LI3_|_XOR|T1
.print DEVI LI3_|_XOR|T2
.print DEVI LI3_|_XOR|Q2
.print DEVI LI3_|_XOR|Q1
.print DEVI LI3_|_AND|A1
.print DEVI LI3_|_AND|A2
.print DEVI LI3_|_AND|A3
.print DEVI LI3_|_AND|B1
.print DEVI LI3_|_AND|B2
.print DEVI LI3_|_AND|B3
.print DEVI LI3_|_AND|Q3
.print DEVI LI3_|_AND|Q2
.print DEVI LI3_|_AND|Q1
.print DEVI LSPL_IG0_0_|I_D1|B
.print DEVI ISPL_IG0_0_|I_D1|B
.print DEVI LSPL_IG0_0_|I_D2|B
.print DEVI ISPL_IG0_0_|I_D2|B
.print DEVI LSPL_IG0_0_|I_Q1|B
.print DEVI ISPL_IG0_0_|I_Q1|B
.print DEVI LSPL_IG0_0_|I_Q2|B
.print DEVI ISPL_IG0_0_|I_Q2|B
.print DEVI BSPL_IG0_0_|1|1
.print DEVI LSPL_IG0_0_|1|P
.print DEVI RSPL_IG0_0_|1|B
.print DEVI LSPL_IG0_0_|1|RB
.print DEVI BSPL_IG0_0_|2|1
.print DEVI LSPL_IG0_0_|2|P
.print DEVI RSPL_IG0_0_|2|B
.print DEVI LSPL_IG0_0_|2|RB
.print DEVI BSPL_IG0_0_|A|1
.print DEVI LSPL_IG0_0_|A|P
.print DEVI RSPL_IG0_0_|A|B
.print DEVI LSPL_IG0_0_|A|RB
.print DEVI BSPL_IG0_0_|B|1
.print DEVI LSPL_IG0_0_|B|P
.print DEVI RSPL_IG0_0_|B|B
.print DEVI LSPL_IG0_0_|B|RB
.print DEVI LSPL_IP1_0_|I_D1|B
.print DEVI ISPL_IP1_0_|I_D1|B
.print DEVI LSPL_IP1_0_|I_D2|B
.print DEVI ISPL_IP1_0_|I_D2|B
.print DEVI LSPL_IP1_0_|I_Q1|B
.print DEVI ISPL_IP1_0_|I_Q1|B
.print DEVI LSPL_IP1_0_|I_Q2|B
.print DEVI ISPL_IP1_0_|I_Q2|B
.print DEVI BSPL_IP1_0_|1|1
.print DEVI LSPL_IP1_0_|1|P
.print DEVI RSPL_IP1_0_|1|B
.print DEVI LSPL_IP1_0_|1|RB
.print DEVI BSPL_IP1_0_|2|1
.print DEVI LSPL_IP1_0_|2|P
.print DEVI RSPL_IP1_0_|2|B
.print DEVI LSPL_IP1_0_|2|RB
.print DEVI BSPL_IP1_0_|A|1
.print DEVI LSPL_IP1_0_|A|P
.print DEVI RSPL_IP1_0_|A|B
.print DEVI LSPL_IP1_0_|A|RB
.print DEVI BSPL_IP1_0_|B|1
.print DEVI LSPL_IP1_0_|B|P
.print DEVI RSPL_IP1_0_|B|B
.print DEVI LSPL_IP1_0_|B|RB
.print DEVI LSPL_IP2_0_|SPL1|1
.print DEVI LSPL_IP2_0_|SPL1|2
.print DEVI LSPL_IP2_0_|SPL1|3
.print DEVI LSPL_IP2_0_|SPL1|4
.print DEVI LSPL_IP2_0_|SPL1|5
.print DEVI LSPL_IP2_0_|SPL1|6
.print DEVI LSPL_IP2_0_|SPL1|7
.print DEVI LSPL_IP2_0_|SPL2|1
.print DEVI LSPL_IP2_0_|SPL2|2
.print DEVI LSPL_IP2_0_|SPL2|3
.print DEVI LSPL_IP2_0_|SPL2|4
.print DEVI LSPL_IP2_0_|SPL2|5
.print DEVI LSPL_IP2_0_|SPL2|6
.print DEVI LSPL_IP2_0_|SPL2|7
.print DEVI LSPL_IG2_0_|I_D1|B
.print DEVI ISPL_IG2_0_|I_D1|B
.print DEVI LSPL_IG2_0_|I_D2|B
.print DEVI ISPL_IG2_0_|I_D2|B
.print DEVI LSPL_IG2_0_|I_Q1|B
.print DEVI ISPL_IG2_0_|I_Q1|B
.print DEVI LSPL_IG2_0_|I_Q2|B
.print DEVI ISPL_IG2_0_|I_Q2|B
.print DEVI BSPL_IG2_0_|1|1
.print DEVI LSPL_IG2_0_|1|P
.print DEVI RSPL_IG2_0_|1|B
.print DEVI LSPL_IG2_0_|1|RB
.print DEVI BSPL_IG2_0_|2|1
.print DEVI LSPL_IG2_0_|2|P
.print DEVI RSPL_IG2_0_|2|B
.print DEVI LSPL_IG2_0_|2|RB
.print DEVI BSPL_IG2_0_|A|1
.print DEVI LSPL_IG2_0_|A|P
.print DEVI RSPL_IG2_0_|A|B
.print DEVI LSPL_IG2_0_|A|RB
.print DEVI BSPL_IG2_0_|B|1
.print DEVI LSPL_IG2_0_|B|P
.print DEVI RSPL_IG2_0_|B|B
.print DEVI LSPL_IG2_0_|B|RB
.print DEVI LSPL_IP3_0_|I_D1|B
.print DEVI ISPL_IP3_0_|I_D1|B
.print DEVI LSPL_IP3_0_|I_D2|B
.print DEVI ISPL_IP3_0_|I_D2|B
.print DEVI LSPL_IP3_0_|I_Q1|B
.print DEVI ISPL_IP3_0_|I_Q1|B
.print DEVI LSPL_IP3_0_|I_Q2|B
.print DEVI ISPL_IP3_0_|I_Q2|B
.print DEVI BSPL_IP3_0_|1|1
.print DEVI LSPL_IP3_0_|1|P
.print DEVI RSPL_IP3_0_|1|B
.print DEVI LSPL_IP3_0_|1|RB
.print DEVI BSPL_IP3_0_|2|1
.print DEVI LSPL_IP3_0_|2|P
.print DEVI RSPL_IP3_0_|2|B
.print DEVI LSPL_IP3_0_|2|RB
.print DEVI BSPL_IP3_0_|A|1
.print DEVI LSPL_IP3_0_|A|P
.print DEVI RSPL_IP3_0_|A|B
.print DEVI LSPL_IP3_0_|A|RB
.print DEVI BSPL_IP3_0_|B|1
.print DEVI LSPL_IP3_0_|B|P
.print DEVI RSPL_IP3_0_|B|B
.print DEVI LSPL_IP3_0_|B|RB
.print DEVI L_PG0_01_|P|1
.print DEVI L_PG0_01_|P|2
.print DEVI L_PG0_01_|P|3
.print DEVI L_PG0_01_|P|T
.print DEVI L_PG0_01_|P|4
.print DEVI L_PG0_01_|P|5
.print DEVI L_PG0_01_|P|6
.print DEVI L_PG0_01_|G|1
.print DEVI L_PG0_01_|G|2
.print DEVI L_PG0_01_|G|3
.print DEVI L_PG0_01_|G|T
.print DEVI L_PG0_01_|G|4
.print DEVI L_PG0_01_|G|5
.print DEVI L_PG0_01_|G|6
.print DEVI L_PG1_01_|_SPL_G1|1
.print DEVI L_PG1_01_|_SPL_G1|2
.print DEVI L_PG1_01_|_SPL_G1|3
.print DEVI L_PG1_01_|_SPL_G1|4
.print DEVI L_PG1_01_|_SPL_G1|5
.print DEVI L_PG1_01_|_SPL_G1|6
.print DEVI L_PG1_01_|_SPL_G1|7
.print DEVI L_PG1_01_|_PG|A1
.print DEVI L_PG1_01_|_PG|A2
.print DEVI L_PG1_01_|_PG|A3
.print DEVI L_PG1_01_|_PG|B1
.print DEVI L_PG1_01_|_PG|B2
.print DEVI L_PG1_01_|_PG|B3
.print DEVI L_PG1_01_|_PG|Q3
.print DEVI L_PG1_01_|_PG|Q2
.print DEVI L_PG1_01_|_PG|Q1
.print DEVI L_PG1_01_|_GG|A1
.print DEVI L_PG1_01_|_GG|A2
.print DEVI L_PG1_01_|_GG|A3
.print DEVI L_PG1_01_|_GG|B1
.print DEVI L_PG1_01_|_GG|B2
.print DEVI L_PG1_01_|_GG|B3
.print DEVI L_PG1_01_|_GG|Q3
.print DEVI L_PG1_01_|_GG|Q2
.print DEVI L_PG1_01_|_GG|Q1
.print DEVI L_PG1_01_|_DFF_PG|1
.print DEVI L_PG1_01_|_DFF_PG|2
.print DEVI L_PG1_01_|_DFF_PG|3
.print DEVI L_PG1_01_|_DFF_PG|T
.print DEVI L_PG1_01_|_DFF_PG|4
.print DEVI L_PG1_01_|_DFF_PG|5
.print DEVI L_PG1_01_|_DFF_PG|6
.print DEVI L_PG1_01_|_DFF_GG|1
.print DEVI L_PG1_01_|_DFF_GG|2
.print DEVI L_PG1_01_|_DFF_GG|3
.print DEVI L_PG1_01_|_DFF_GG|T
.print DEVI L_PG1_01_|_DFF_GG|4
.print DEVI L_PG1_01_|_DFF_GG|5
.print DEVI L_PG1_01_|_DFF_GG|6
.print DEVI L_PG1_01_|_AND_G|A1
.print DEVI L_PG1_01_|_AND_G|A2
.print DEVI L_PG1_01_|_AND_G|A3
.print DEVI L_PG1_01_|_AND_G|B1
.print DEVI L_PG1_01_|_AND_G|B2
.print DEVI L_PG1_01_|_AND_G|B3
.print DEVI L_PG1_01_|_AND_G|Q3
.print DEVI L_PG1_01_|_AND_G|Q2
.print DEVI L_PG1_01_|_AND_G|Q1
.print DEVI L_PG2_01_|P|1
.print DEVI L_PG2_01_|P|2
.print DEVI L_PG2_01_|P|3
.print DEVI L_PG2_01_|P|T
.print DEVI L_PG2_01_|P|4
.print DEVI L_PG2_01_|P|5
.print DEVI L_PG2_01_|P|6
.print DEVI L_PG2_01_|G|1
.print DEVI L_PG2_01_|G|2
.print DEVI L_PG2_01_|G|3
.print DEVI L_PG2_01_|G|T
.print DEVI L_PG2_01_|G|4
.print DEVI L_PG2_01_|G|5
.print DEVI L_PG2_01_|G|6
.print DEVI L_PG3_01_|_SPL_G1|1
.print DEVI L_PG3_01_|_SPL_G1|2
.print DEVI L_PG3_01_|_SPL_G1|3
.print DEVI L_PG3_01_|_SPL_G1|4
.print DEVI L_PG3_01_|_SPL_G1|5
.print DEVI L_PG3_01_|_SPL_G1|6
.print DEVI L_PG3_01_|_SPL_G1|7
.print DEVI L_PG3_01_|_SPL_P1|1
.print DEVI L_PG3_01_|_SPL_P1|2
.print DEVI L_PG3_01_|_SPL_P1|3
.print DEVI L_PG3_01_|_SPL_P1|4
.print DEVI L_PG3_01_|_SPL_P1|5
.print DEVI L_PG3_01_|_SPL_P1|6
.print DEVI L_PG3_01_|_SPL_P1|7
.print DEVI L_PG3_01_|_PG|A1
.print DEVI L_PG3_01_|_PG|A2
.print DEVI L_PG3_01_|_PG|A3
.print DEVI L_PG3_01_|_PG|B1
.print DEVI L_PG3_01_|_PG|B2
.print DEVI L_PG3_01_|_PG|B3
.print DEVI L_PG3_01_|_PG|Q3
.print DEVI L_PG3_01_|_PG|Q2
.print DEVI L_PG3_01_|_PG|Q1
.print DEVI L_PG3_01_|_GG|A1
.print DEVI L_PG3_01_|_GG|A2
.print DEVI L_PG3_01_|_GG|A3
.print DEVI L_PG3_01_|_GG|B1
.print DEVI L_PG3_01_|_GG|B2
.print DEVI L_PG3_01_|_GG|B3
.print DEVI L_PG3_01_|_GG|Q3
.print DEVI L_PG3_01_|_GG|Q2
.print DEVI L_PG3_01_|_GG|Q1
.print DEVI L_PG3_01_|_DFF_P0|1
.print DEVI L_PG3_01_|_DFF_P0|2
.print DEVI L_PG3_01_|_DFF_P0|3
.print DEVI L_PG3_01_|_DFF_P0|T
.print DEVI L_PG3_01_|_DFF_P0|4
.print DEVI L_PG3_01_|_DFF_P0|5
.print DEVI L_PG3_01_|_DFF_P0|6
.print DEVI L_PG3_01_|_DFF_P1|1
.print DEVI L_PG3_01_|_DFF_P1|2
.print DEVI L_PG3_01_|_DFF_P1|3
.print DEVI L_PG3_01_|_DFF_P1|T
.print DEVI L_PG3_01_|_DFF_P1|4
.print DEVI L_PG3_01_|_DFF_P1|5
.print DEVI L_PG3_01_|_DFF_P1|6
.print DEVI L_PG3_01_|_DFF_PG|1
.print DEVI L_PG3_01_|_DFF_PG|2
.print DEVI L_PG3_01_|_DFF_PG|3
.print DEVI L_PG3_01_|_DFF_PG|T
.print DEVI L_PG3_01_|_DFF_PG|4
.print DEVI L_PG3_01_|_DFF_PG|5
.print DEVI L_PG3_01_|_DFF_PG|6
.print DEVI L_PG3_01_|_DFF_GG|1
.print DEVI L_PG3_01_|_DFF_GG|2
.print DEVI L_PG3_01_|_DFF_GG|3
.print DEVI L_PG3_01_|_DFF_GG|T
.print DEVI L_PG3_01_|_DFF_GG|4
.print DEVI L_PG3_01_|_DFF_GG|5
.print DEVI L_PG3_01_|_DFF_GG|6
.print DEVI L_PG3_01_|_AND_G|A1
.print DEVI L_PG3_01_|_AND_G|A2
.print DEVI L_PG3_01_|_AND_G|A3
.print DEVI L_PG3_01_|_AND_G|B1
.print DEVI L_PG3_01_|_AND_G|B2
.print DEVI L_PG3_01_|_AND_G|B3
.print DEVI L_PG3_01_|_AND_G|Q3
.print DEVI L_PG3_01_|_AND_G|Q2
.print DEVI L_PG3_01_|_AND_G|Q1
.print DEVI L_PG3_01_|_AND_P|A1
.print DEVI L_PG3_01_|_AND_P|A2
.print DEVI L_PG3_01_|_AND_P|A3
.print DEVI L_PG3_01_|_AND_P|B1
.print DEVI L_PG3_01_|_AND_P|B2
.print DEVI L_PG3_01_|_AND_P|B3
.print DEVI L_PG3_01_|_AND_P|Q3
.print DEVI L_PG3_01_|_AND_P|Q2
.print DEVI L_PG3_01_|_AND_P|Q1
.print DEVI L_DFF_IP1_01_|I_1|B
.print DEVI I_DFF_IP1_01_|I_1|B
.print DEVI L_DFF_IP1_01_|I_3|B
.print DEVI I_DFF_IP1_01_|I_3|B
.print DEVI L_DFF_IP1_01_|I_T|B
.print DEVI I_DFF_IP1_01_|I_T|B
.print DEVI L_DFF_IP1_01_|I_6|B
.print DEVI I_DFF_IP1_01_|I_6|B
.print DEVI B_DFF_IP1_01_|1|1
.print DEVI L_DFF_IP1_01_|1|P
.print DEVI R_DFF_IP1_01_|1|B
.print DEVI L_DFF_IP1_01_|1|RB
.print DEVI B_DFF_IP1_01_|23|1
.print DEVI R_DFF_IP1_01_|23|B
.print DEVI L_DFF_IP1_01_|23|RB
.print DEVI B_DFF_IP1_01_|3|1
.print DEVI L_DFF_IP1_01_|3|P
.print DEVI R_DFF_IP1_01_|3|B
.print DEVI L_DFF_IP1_01_|3|RB
.print DEVI B_DFF_IP1_01_|4|1
.print DEVI L_DFF_IP1_01_|4|P
.print DEVI R_DFF_IP1_01_|4|B
.print DEVI L_DFF_IP1_01_|4|RB
.print DEVI B_DFF_IP1_01_|T|1
.print DEVI L_DFF_IP1_01_|T|P
.print DEVI R_DFF_IP1_01_|T|B
.print DEVI L_DFF_IP1_01_|T|RB
.print DEVI B_DFF_IP1_01_|45|1
.print DEVI R_DFF_IP1_01_|45|B
.print DEVI L_DFF_IP1_01_|45|RB
.print DEVI B_DFF_IP1_01_|6|1
.print DEVI L_DFF_IP1_01_|6|P
.print DEVI R_DFF_IP1_01_|6|B
.print DEVI L_DFF_IP1_01_|6|RB
.print DEVI L_DFF_IP2_01_|I_1|B
.print DEVI I_DFF_IP2_01_|I_1|B
.print DEVI L_DFF_IP2_01_|I_3|B
.print DEVI I_DFF_IP2_01_|I_3|B
.print DEVI L_DFF_IP2_01_|I_T|B
.print DEVI I_DFF_IP2_01_|I_T|B
.print DEVI L_DFF_IP2_01_|I_6|B
.print DEVI I_DFF_IP2_01_|I_6|B
.print DEVI B_DFF_IP2_01_|1|1
.print DEVI L_DFF_IP2_01_|1|P
.print DEVI R_DFF_IP2_01_|1|B
.print DEVI L_DFF_IP2_01_|1|RB
.print DEVI B_DFF_IP2_01_|23|1
.print DEVI R_DFF_IP2_01_|23|B
.print DEVI L_DFF_IP2_01_|23|RB
.print DEVI B_DFF_IP2_01_|3|1
.print DEVI L_DFF_IP2_01_|3|P
.print DEVI R_DFF_IP2_01_|3|B
.print DEVI L_DFF_IP2_01_|3|RB
.print DEVI B_DFF_IP2_01_|4|1
.print DEVI L_DFF_IP2_01_|4|P
.print DEVI R_DFF_IP2_01_|4|B
.print DEVI L_DFF_IP2_01_|4|RB
.print DEVI B_DFF_IP2_01_|T|1
.print DEVI L_DFF_IP2_01_|T|P
.print DEVI R_DFF_IP2_01_|T|B
.print DEVI L_DFF_IP2_01_|T|RB
.print DEVI B_DFF_IP2_01_|45|1
.print DEVI R_DFF_IP2_01_|45|B
.print DEVI L_DFF_IP2_01_|45|RB
.print DEVI B_DFF_IP2_01_|6|1
.print DEVI L_DFF_IP2_01_|6|P
.print DEVI R_DFF_IP2_01_|6|B
.print DEVI L_DFF_IP2_01_|6|RB
.print DEVI L_DFF_IP3_01_|I_1|B
.print DEVI I_DFF_IP3_01_|I_1|B
.print DEVI L_DFF_IP3_01_|I_3|B
.print DEVI I_DFF_IP3_01_|I_3|B
.print DEVI L_DFF_IP3_01_|I_T|B
.print DEVI I_DFF_IP3_01_|I_T|B
.print DEVI L_DFF_IP3_01_|I_6|B
.print DEVI I_DFF_IP3_01_|I_6|B
.print DEVI B_DFF_IP3_01_|1|1
.print DEVI L_DFF_IP3_01_|1|P
.print DEVI R_DFF_IP3_01_|1|B
.print DEVI L_DFF_IP3_01_|1|RB
.print DEVI B_DFF_IP3_01_|23|1
.print DEVI R_DFF_IP3_01_|23|B
.print DEVI L_DFF_IP3_01_|23|RB
.print DEVI B_DFF_IP3_01_|3|1
.print DEVI L_DFF_IP3_01_|3|P
.print DEVI R_DFF_IP3_01_|3|B
.print DEVI L_DFF_IP3_01_|3|RB
.print DEVI B_DFF_IP3_01_|4|1
.print DEVI L_DFF_IP3_01_|4|P
.print DEVI R_DFF_IP3_01_|4|B
.print DEVI L_DFF_IP3_01_|4|RB
.print DEVI B_DFF_IP3_01_|T|1
.print DEVI L_DFF_IP3_01_|T|P
.print DEVI R_DFF_IP3_01_|T|B
.print DEVI L_DFF_IP3_01_|T|RB
.print DEVI B_DFF_IP3_01_|45|1
.print DEVI R_DFF_IP3_01_|45|B
.print DEVI L_DFF_IP3_01_|45|RB
.print DEVI B_DFF_IP3_01_|6|1
.print DEVI L_DFF_IP3_01_|6|P
.print DEVI R_DFF_IP3_01_|6|B
.print DEVI L_DFF_IP3_01_|6|RB
.print DEVI LSPL_G1_1_|SPL1|1
.print DEVI LSPL_G1_1_|SPL1|2
.print DEVI LSPL_G1_1_|SPL1|3
.print DEVI LSPL_G1_1_|SPL1|4
.print DEVI LSPL_G1_1_|SPL1|5
.print DEVI LSPL_G1_1_|SPL1|6
.print DEVI LSPL_G1_1_|SPL1|7
.print DEVI LSPL_G1_1_|SPL2|1
.print DEVI LSPL_G1_1_|SPL2|2
.print DEVI LSPL_G1_1_|SPL2|3
.print DEVI LSPL_G1_1_|SPL2|4
.print DEVI LSPL_G1_1_|SPL2|5
.print DEVI LSPL_G1_1_|SPL2|6
.print DEVI LSPL_G1_1_|SPL2|7
.print V I1_|_XOR|Q1
.print V _PG3_01_|_DFF_GG|A2
.print V I1_|_SPL_B|D1
.print V T02_
.print V _DFF_IP2_01_|4|MID_SERIES
.print V I0_|_DFF_A|T1
.print V _PG3_01_|_DFF_GG|A3
.print V I0_|_AND|A2
.print V _PG1_01_|_SPL_G1|JCT
.print V I1_|_AND|B2
.print V G1_1_TO1_
.print V _PG2_01_|G|T1
.print V _DFF_IP3_01_|23|MID_SHUNT
.print V I3_|_XOR|ABTQ
.print V IP1_0_
.print V _PG3_01_|_AND_P|Q1
.print V I3_|_DFF_A|A2
.print V SPL_IP3_0_|2|MID_SERIES
.print V SPL_IP1_0_|I_Q1|MID
.print V _PG3_01_|GG_SYNC
.print V I2_|_XOR|T2
.print V I1_|_AND|Q1
.print V _PG1_01_|_PG|B3
.print V _PG3_01_|_DFF_P0|A4
.print V I0_|_DFF_B|Q1
.print V _PG3_01_|_DFF_P1|T2
.print V I0_|_DFF_A|A3
.print V SPL_G1_1_|SPL1|D1
.print V I2_|A1
.print V SPL_IP2_0_|SPL1|D2
.print V _PG3_01_|_DFF_GG|Q1
.print V _PG3_01_|_AND_G|Q2
.print V SPL_IP3_0_|1|MID_SHUNT
.print V SPL_IG2_0_|I_D2|MID
.print V I0_|_SPL_A|QA1
.print V I1_|_XOR|A2
.print V _DFF_IP1_01_|4|MID_SERIES
.print V _DFF_IP2_01_|4|MID_SHUNT
.print V I2_|_DFF_A|A3
.print V _PG3_01_|_DFF_PG|A1
.print V _DFF_IP3_01_|45|MID_SHUNT
.print V _PG1_01_|_PG|B2
.print V _PG3_01_|_SPL_P1|QB1
.print V SPL_IG2_0_|2|MID_SERIES
.print V _DFF_IP1_01_|T|MID_SERIES
.print V _PG3_01_|_DFF_P0|Q1
.print V I3_|_AND|A1
.print V I0_|B1
.print V _DFF_IP1_01_|I_T|MID
.print V _PG1_01_|_DFF_GG|T2
.print V _PG3_01_|_AND_P|B3
.print V SPL_IP1_0_|2|MID_SHUNT
.print V I0_|_XOR|A1
.print V _DFF_IP1_01_|6|MID_SHUNT
.print V I1_|_DFF_B|A4
.print V _DFF_IP2_01_|A3
.print V I2_|_XOR|Q1
.print V _PG0_01_|P|T2
.print V _PG3_01_|P1_COPY_2
.print V _DFF_IP2_01_|T|MID_SHUNT
.print V I0_|_SPL_B|JCT
.print V I1_|_XOR|ABTQ
.print V _PG3_01_|_PG|B2
.print V SPL_IP2_0_|SPL1|D1
.print V I0_|_AND|A3
.print V _PG3_01_|_DFF_P0|A3
.print V I3_|_XOR|A1
.print V P3_1
.print V _DFF_IP1_01_|1|MID_SHUNT
.print V _PG2_01_|G|T2
.print V SPL_IP3_0_|JCT
.print V _PG3_01_|_DFF_PG|A4
.print V I0_|_AND|Q1
.print V _DFF_IP2_01_|T2
.print V _PG3_01_|GG
.print V IP2_0_TO2_
.print V SPL_IG0_0_|QA1
.print V I1_|_AND|A1
.print V _PG2_01_|G|A3
.print V I1_|_SPL_A|QA1
.print V I1_|B2
.print V _PG3_01_|_AND_G|A2
.print V _DFF_IP3_01_|A1
.print V IG0_0_
.print V _DFF_IP1_01_|1|MID_SERIES
.print V I1_|_DFF_A|A1
.print V _PG3_01_|_SPL_G1|QB1
.print V _PG3_01_|_GG|A2
.print V I3_|_DFF_B|A3
.print V _DFF_IP3_01_|T2
.print V I1_|_DFF_A|A3
.print V SPL_IG2_0_|A|MID_SERIES
.print V _DFF_IP3_01_|3|MID_SHUNT
.print V _PG3_01_|_DFF_GG|A4
.print V I3_|_SPL_B|D1
.print V I2_|B2
.print V SPL_IP1_0_|I_D2|MID
.print V IP2_0_OUT_
.print V I0_|_XOR|Q1
.print V _PG3_01_|_AND_P|B1
.print V _PG3_01_|_GG|B2
.print V I0_|_AND|B2
.print V I3_|A2
.print V _PG1_01_|_SPL_G1|D1
.print V I3_|_SPL_B|QA1
.print V _PG3_01_|_SPL_P1|QA1
.print V _DFF_IP1_01_|T|MID_SHUNT
.print V P0_1
.print V SPL_IG2_0_|I_D1|MID
.print V G1_1_
.print V _PG0_01_|P|A1
.print V I1_|B1_SYNC
.print V I3_|_XOR|T2
.print V _DFF_IP1_01_|A4
.print V SPL_IP3_0_|B|MID_SERIES
.print V _PG0_01_|G|A3
.print V _PG3_01_|_GG|Q2
.print V _PG1_01_|_GG|Q2
.print V _PG1_01_|PG_SYNC
.print V P1_1_TO2
.print V SPL_IP3_0_|I_D2|MID
.print V _PG0_01_|P|A3
.print V SPL_IP2_0_|SPL2|QB1
.print V _PG0_01_|G|A1
.print V I1_|_SPL_A|JCT
.print V I0_|_SPL_A|D1
.print V _PG3_01_|_PG|A2
.print V _DFF_IP2_01_|A2
.print V G1_1_TO1
.print V I2_|_AND|A3
.print V SPL_IP1_0_|D2
.print V I2_|_AND|B2
.print V _PG3_01_|_AND_G|B1
.print V _PG1_01_|_DFF_PG|Q1
.print V _PG3_01_|_AND_P|Q2
.print V SPL_IP1_0_|B|MID_SERIES
.print V I3_|_DFF_B|A2
.print V I3_|_SPL_A|QB1
.print V I3_|_XOR|Q1
.print V I2_|_DFF_B|A3
.print V SPL_IP2_0_|SPL2|QA1
.print V I3_|_SPL_A|QA1
.print V I3_|A1_SYNC
.print V I1_|_AND|B3
.print V IP2_0_
.print V I1_|_SPL_A|D1
.print V _PG3_01_|_AND_G|Q1
.print V SPL_IG2_0_|1|MID_SERIES
.print V G0_1
.print V I2_|_AND|A2
.print V I2_|_AND|Q2
.print V I0_|_DFF_B|T2
.print V _PG1_01_|_DFF_PG|A4
.print V SPL_IG0_0_|2|MID_SERIES
.print V A0_
.print V I3_|_DFF_A|A4
.print V _PG1_01_|_DFF_GG|A3
.print V SPL_IG0_0_|I_Q1|MID
.print V I3_|_DFF_A|A1
.print V SPL_IG0_0_|2|MID_SHUNT
.print V B0_
.print V I3_|_DFF_A|T2
.print V _PG3_01_|_DFF_GG|T1
.print V _DFF_IP2_01_|T|MID_SERIES
.print V _DFF_IP1_01_|6|MID_SERIES
.print V _PG3_01_|_PG|B1
.print V I2_|_XOR|B2
.print V _PG0_01_|P|Q1
.print V _DFF_IP2_01_|3|MID_SHUNT
.print V SPL_IG0_0_|JCT
.print V I2_|_SPL_A|QB1
.print V _DFF_IP2_01_|A4
.print V I1_|_XOR|AB
.print V I3_|_SPL_A|D2
.print V I1_|_XOR|B2
.print V I3_|_DFF_B|T1
.print V _PG3_01_|_SPL_G1|JCT
.print V _PG3_01_|_PG|Q3
.print V _DFF_IP3_01_|T|MID_SERIES
.print V I2_|_DFF_A|T2
.print V _DFF_IP1_01_|A1
.print V _DFF_IP3_01_|Q1
.print V SPL_IP3_0_|QA1
.print V SPL_IG0_0_|1|MID_SERIES
.print V I3_|_XOR|B1
.print V I2_|_DFF_B|A2
.print V I3_|_DFF_B|A4
.print V SPL_IG0_0_|QB1
.print V _PG2_01_|P|A4
.print V _PG1_01_|_SPL_G1|QA1
.print V SPL_IP3_0_|I_D1|MID
.print V SPL_IP2_0_|SPL2|JCT
.print V SPL_IG2_0_|A|MID_SHUNT
.print V IP2_0_TO3_
.print V I2_|_AND|B1
.print V SPL_IP1_0_|B|MID_SHUNT
.print V I2_|_SPL_A|D1
.print V SPL_IP1_0_|QA1
.print V I1_|_SPL_A|D2
.print V D03_
.print V _DFF_IP1_01_|T1
.print V _PG3_01_|_DFF_GG|A1
.print V I2_|B1
.print V I3_|_DFF_A|A3
.print V I0_|_AND|Q2
.print V SPL_IG2_0_|1|MID_SHUNT
.print V IP3_0_
.print V SPL_IP2_0_|SPL2|D1
.print V _PG3_01_|_PG|A3
.print V _DFF_IP3_01_|A2
.print V _PG0_01_|G|A2
.print V D02_
.print V G1_1_TO2
.print V I1_|_AND|A2
.print V I0_|_XOR|A2
.print V P1_1_TO1
.print V SPL_IG0_0_|I_D1|MID
.print V I1_|_AND|B1
.print V SPL_IP3_0_|D1
.print V SPL_IG2_0_|B|MID_SERIES
.print V IP2_1_OUT
.print V _PG0_01_|P|A4
.print V _PG1_01_|_AND_G|Q2
.print V _PG3_01_|_DFF_P0|T2
.print V _DFF_IP1_01_|I_1|MID
.print V _DFF_IP1_01_|45|MID_SHUNT
.print V I0_|_XOR|ABTQ
.print V I2_|_XOR|A2
.print V _DFF_IP3_01_|6|MID_SERIES
.print V _DFF_IP2_01_|1|MID_SERIES
.print V SPL_IG2_0_|JCT
.print V SPL_IP1_0_|D1
.print V G0_1_
.print V I2_|_DFF_B|A4
.print V I0_|_SPL_A|QB1
.print V T07_
.print V G1_1_TO3_
.print V I2_|_XOR|B1
.print V SPL_IG2_0_|QB1
.print V _DFF_IP3_01_|4|MID_SHUNT
.print V I2_|B1_SYNC
.print V _PG1_01_|G1_COPY_2
.print V _DFF_IP3_01_|3|MID_SERIES
.print V SPL_G1_1_|SPL1|QA1
.print V _DFF_IP3_01_|I_3|MID
.print V _PG3_01_|_PG|B3
.print V I0_|_SPL_A|JCT
.print V _PG2_01_|G|A4
.print V _DFF_IP3_01_|I_6|MID
.print V I0_|_DFF_A|A1
.print V _DFF_IP2_01_|A1
.print V _DFF_IP3_01_|6|MID_SHUNT
.print V I3_|_XOR|B2
.print V SPL_G1_1_|SPL2|JCT
.print V _DFF_IP1_01_|I_6|MID
.print V I1_|A1
.print V I1_|_XOR|A3
.print V _PG3_01_|P0_SYNC
.print V I1_|_SPL_A|QB1
.print V _PG3_01_|_PG|Q2
.print V _DFF_IP1_01_|T2
.print V I2_|_XOR|AB
.print V I1_|_SPL_B|D2
.print V _PG1_01_|PG
.print V _DFF_IP3_01_|T|MID_SHUNT
.print V SPL_IP2_0_|SPL2|D2
.print V I0_|_XOR|AB
.print V _PG1_01_|_GG|Q3
.print V _PG1_01_|_GG|A3
.print V _PG1_01_|_PG|A2
.print V IP0_0_
.print V I0_|_XOR|A3
.print V P2_1_
.print V I2_|_DFF_B|A1
.print V _DFF_IP2_01_|I_T|MID
.print V IG3_0_
.print V T01_
.print V SPL_IG2_0_|I_Q1|MID
.print V _PG1_01_|_DFF_GG|Q1
.print V SPL_IP3_0_|A|MID_SHUNT
.print V SPL_IP3_0_|2|MID_SHUNT
.print V _PG3_01_|_DFF_P1|A1
.print V SPL_G1_1_|SPL1|JCT
.print V _PG1_01_|_AND_G|A1
.print V I0_|_XOR|B3
.print V I2_|_DFF_A|Q1
.print V I0_|_DFF_B|A1
.print V SPL_IG0_0_|D1
.print V B2_
.print V SPL_IG2_0_|D1
.print V IP3_0_OUT_
.print V _PG3_01_|G1_COPY_2
.print V _PG3_01_|_DFF_PG|T1
.print V _PG3_01_|_GG|Q1
.print V SPL_IP2_0_|QTMP
.print V _PG1_01_|_AND_G|Q3
.print V _PG2_01_|P|A3
.print V _PG3_01_|_DFF_P1|Q1
.print V I3_|_XOR|A3
.print V IP3_0_TO1_
.print V I2_|_DFF_A|T1
.print V SPL_G1_1_|SPL1|D2
.print V I1_|_DFF_B|T2
.print V I0_|_XOR|B2
.print V I3_|_DFF_B|Q1
.print V G2_1
.print V P3_1_
.print V I3_|_AND|B2
.print V I3_|_DFF_A|Q1
.print V _DFF_IP3_01_|1|MID_SERIES
.print V I0_|_AND|Q3
.print V I3_|_AND|A2
.print V _PG3_01_|_DFF_PG|T2
.print V SPL_IG0_0_|B|MID_SHUNT
.print V _DFF_IP1_01_|3|MID_SERIES
.print V B1_
.print V IP1_0_OUT_
.print V _PG2_01_|P|Q1
.print V _DFF_IP2_01_|23|MID_SHUNT
.print V A2_
.print V A1_
.print V I1_|_AND|Q3
.print V SPL_IP2_0_|SPL1|JCT
.print V I3_|_AND|B1
.print V I3_|_DFF_A|T1
.print V I0_|_SPL_B|D2
.print V _PG3_01_|_GG|Q3
.print V I3_|_SPL_B|D2
.print V _PG1_01_|_SPL_G1|QB1
.print V I2_|_SPL_B|JCT
.print V _PG0_01_|G|T1
.print V _PG3_01_|_AND_G|Q3
.print V _PG1_01_|_PG|A1
.print V _PG3_01_|_AND_P|A1
.print V I0_|A2
.print V I1_|_DFF_B|A3
.print V _PG3_01_|_DFF_PG|Q1
.print V I2_|_XOR|T1
.print V _DFF_IP2_01_|Q1
.print V G3_1
.print V I3_|_AND|A3
.print V _PG3_01_|_DFF_P1|A4
.print V SPL_IG2_0_|I_Q2|MID
.print V IP3_1_OUT
.print V _PG1_01_|GG_SYNC
.print V _DFF_IP2_01_|3|MID_SERIES
.print V _DFF_IP3_01_|A4
.print V _PG0_01_|G|Q1
.print V _PG2_01_|P|A2
.print V SPL_IP3_0_|I_Q2|MID
.print V _PG3_01_|_DFF_PG|A2
.print V SPL_IP2_0_|SPL1|QB1
.print V _PG3_01_|_DFF_P0|A2
.print V _PG3_01_|G1_COPY_1
.print V IP3_1_OUT_
.print V _PG3_01_|PG
.print V SPL_IG0_0_|A|MID_SHUNT
.print V _PG3_01_|_SPL_G1|QA1
.print V _DFF_IP1_01_|A2
.print V SPL_IP3_0_|I_Q1|MID
.print V SPL_IP1_0_|1|MID_SERIES
.print V I3_|_SPL_A|D1
.print V SPL_G1_1_|SPL2|D1
.print V IG0_0_TO0_
.print V _PG1_01_|_DFF_PG|A2
.print V SPL_G1_1_|SPL2|D2
.print V _PG1_01_|_DFF_PG|A3
.print V T04_
.print V _PG3_01_|_PG|A1
.print V I0_|_DFF_B|A3
.print V I3_|_AND|B3
.print V I2_|_AND|B3
.print V I1_|_DFF_B|Q1
.print V _DFF_IP2_01_|I_3|MID
.print V T05_
.print V _DFF_IP2_01_|T1
.print V IP1_1_OUT_
.print V _PG1_01_|_GG|Q1
.print V I2_|_SPL_B|D2
.print V T00_
.print V I1_|_DFF_A|T2
.print V SPL_IP1_0_|1|MID_SHUNT
.print V I1_|_DFF_A|A4
.print V I1_|_DFF_A|A2
.print V _DFF_IP3_01_|1|MID_SHUNT
.print V I0_|B1_SYNC
.print V _PG1_01_|_AND_G|A2
.print V _DFF_IP1_01_|Q1
.print V I3_|_DFF_B|T2
.print V _PG1_01_|_DFF_GG|T1
.print V SPL_IP3_0_|D2
.print V I0_|_SPL_B|QA1
.print V I1_|_XOR|B3
.print V IP1_0_TO1_
.print V I2_|_DFF_A|A1
.print V SPL_IP1_0_|QB1
.print V SPL_IP3_0_|A|MID_SERIES
.print V _PG3_01_|P1_SYNC
.print V SPL_IP3_0_|B|MID_SHUNT
.print V SPL_IP1_0_|JCT
.print V _DFF_IP2_01_|6|MID_SERIES
.print V _PG3_01_|_SPL_P1|D2
.print V I0_|_SPL_B|QB1
.print V _PG2_01_|P|T1
.print V _DFF_IP3_01_|A3
.print V I0_|_DFF_A|Q1
.print V G1_1_TO3
.print V _PG3_01_|_AND_G|A3
.print V SPL_IG2_0_|2|MID_SHUNT
.print V I1_|_AND|Q2
.print V G2_1_
.print V I1_|_XOR|A1
.print V IG0_0_TO1_
.print V I0_|_DFF_A|T2
.print V I0_|_XOR|T2
.print V I2_|_XOR|B3
.print V _DFF_IP3_01_|I_T|MID
.print V _PG2_01_|G|A1
.print V _PG3_01_|_AND_P|A2
.print V _PG3_01_|_DFF_P1|T1
.print V I0_|_DFF_B|A4
.print V _PG0_01_|G|A4
.print V _PG1_01_|_DFF_GG|A4
.print V I1_|_XOR|T1
.print V I3_|_AND|Q1
.print V _PG2_01_|P|T2
.print V _PG3_01_|_SPL_P1|JCT
.print V _DFF_IP2_01_|I_6|MID
.print V I2_|_DFF_A|A4
.print V _PG1_01_|_DFF_PG|T1
.print V _PG3_01_|_DFF_P1|A2
.print V I2_|_AND|Q3
.print V _PG3_01_|_AND_P|B2
.print V I1_|B1
.print V _PG3_01_|_AND_G|B3
.print V _PG0_01_|P|A2
.print V I1_|_DFF_B|T1
.print V T06_
.print V I2_|_DFF_B|Q1
.print V _PG3_01_|_DFF_PG|A3
.print V IG2_0_
.print V I1_|_DFF_B|A1
.print V _PG1_01_|_GG|A2
.print V _PG1_01_|_PG|A3
.print V I0_|_SPL_B|D1
.print V I2_|A1_SYNC
.print V _PG1_01_|_DFF_GG|A2
.print V SPL_G1_1_|SPL1|QB1
.print V _PG1_01_|_AND_G|A3
.print V I3_|_XOR|T1
.print V I2_|_AND|A1
.print V SPL_G1_1_|QTMP
.print V _DFF_IP1_01_|4|MID_SHUNT
.print V SPL_IG0_0_|A|MID_SERIES
.print V I2_|_DFF_B|T2
.print V I2_|_DFF_B|T1
.print V I3_|B2
.print V _PG3_01_|_DFF_P0|A1
.print V _PG1_01_|_PG|B1
.print V _DFF_IP2_01_|45|MID_SHUNT
.print V _DFF_IP2_01_|I_1|MID
.print V _DFF_IP2_01_|6|MID_SHUNT
.print V I0_|B2
.print V I2_|_SPL_B|QA1
.print V _PG1_01_|_DFF_PG|T2
.print V _DFF_IP3_01_|4|MID_SERIES
.print V _PG0_01_|P|T1
.print V SPL_IP3_0_|1|MID_SERIES
.print V SPL_G1_1_|SPL2|QA1
.print V _PG1_01_|_AND_G|B2
.print V SPL_IG2_0_|B|MID_SHUNT
.print V _PG1_01_|_DFF_PG|A1
.print V I0_|_AND|B1
.print V _PG3_01_|_GG|B1
.print V I0_|_DFF_A|A4
.print V _PG3_01_|_PG|Q1
.print V _PG2_01_|G|Q1
.print V I2_|_SPL_A|QA1
.print V _PG3_01_|_SPL_G1|D1
.print V SPL_IP1_0_|A|MID_SERIES
.print V _PG3_01_|_SPL_G1|D2
.print V I3_|_AND|Q3
.print V I1_|_SPL_B|JCT
.print V _PG1_01_|_AND_G|B3
.print V SPL_IG0_0_|I_D2|MID
.print V I1_|A2
.print V IP2_1_OUT_
.print V I2_|_XOR|A3
.print V _PG1_01_|_PG|Q3
.print V I3_|_XOR|A2
.print V B3_
.print V _PG0_01_|G|T2
.print V IG1_0_
.print V _PG2_01_|P|A1
.print V I1_|A1_SYNC
.print V I3_|_AND|Q2
.print V I0_|_AND|A1
.print V _PG3_01_|_DFF_P1|A3
.print V I0_|_DFF_B|T1
.print V SPL_IP1_0_|I_Q2|MID
.print V _DFF_IP3_01_|I_1|MID
.print V _PG3_01_|_GG|A3
.print V I1_|_SPL_B|QB1
.print V _DFF_IP1_01_|A3
.print V G1_1_TO2_
.print V _PG3_01_|_AND_G|B2
.print V I1_|_DFF_B|A2
.print V P1_1_TO3
.print V _PG1_01_|_GG|B1
.print V _DFF_IP3_01_|T1
.print V I2_|_SPL_A|JCT
.print V _PG1_01_|_PG|Q1
.print V I1_|_DFF_A|T1
.print V I2_|_AND|Q1
.print V SPL_IG0_0_|B|MID_SERIES
.print V _DFF_IP2_01_|1|MID_SHUNT
.print V I0_|_AND|B3
.print V SPL_IP2_0_|SPL1|QA1
.print V I2_|_XOR|A1
.print V SPL_IG0_0_|I_Q2|MID
.print V I1_|_AND|A3
.print V _PG1_01_|_SPL_G1|D2
.print V _PG3_01_|_DFF_GG|T2
.print V I2_|_SPL_B|D1
.print V I3_|_DFF_B|A1
.print V G3_1_
.print V _DFF_IP1_01_|I_3|MID
.print V I2_|A2
.print V _PG3_01_|_DFF_P0|T1
.print V _PG1_01_|_GG|B2
.print V I0_|_XOR|T1
.print V I3_|B1
.print V IG2_0_TO2_
.print V I0_|_XOR|B1
.print V I0_|A1_SYNC
.print V I3_|_XOR|B3
.print V _PG1_01_|_GG|A1
.print V P2_1
.print V I2_|_SPL_A|D2
.print V _PG1_01_|GG
.print V I3_|_XOR|AB
.print V SPL_IP1_0_|2|MID_SERIES
.print V I1_|_SPL_B|QA1
.print V T03_
.print V _PG3_01_|_GG|B3
.print V SPL_IG2_0_|QA1
.print V I0_|_DFF_B|A2
.print V I1_|_XOR|B1
.print V SPL_IP1_0_|I_D1|MID
.print V I2_|_SPL_B|QB1
.print V IP1_1_OUT
.print V D01_
.print V I1_|_DFF_A|Q1
.print V _PG3_01_|PG_SYNC
.print V _PG1_01_|_PG|Q2
.print V I2_|_DFF_A|A2
.print V P0_1_
.print V _PG1_01_|_DFF_GG|A1
.print V IG2_0_TO3_
.print V SPL_G1_1_|SPL2|QB1
.print V SPL_IP1_0_|A|MID_SHUNT
.print V SPL_IG0_0_|D2
.print V _PG1_01_|_GG|B3
.print V _PG3_01_|_SPL_P1|D1
.print V I1_|_XOR|T2
.print V _PG3_01_|P1_COPY_1
.print V _PG1_01_|_AND_G|Q1
.print V I3_|_SPL_B|QB1
.print V SPL_IG0_0_|1|MID_SHUNT
.print V _PG3_01_|_AND_P|A3
.print V SPL_IG2_0_|D2
.print V A3_
.print V _PG2_01_|G|A2
.print V _PG3_01_|_AND_G|A1
.print V _PG3_01_|_GG|A1
.print V _PG3_01_|_AND_P|Q3
.print V I3_|B1_SYNC
.print V I2_|_XOR|ABTQ
.print V I3_|A1
.print V SPL_IP3_0_|QB1
.print V I0_|_SPL_A|D2
.print V I0_|_DFF_A|A2
.print V _DFF_IP1_01_|23|MID_SHUNT
.print V I3_|_SPL_A|JCT
.print V _PG1_01_|G1_COPY_1
.print V I3_|_SPL_B|JCT
.print V I0_|A1
.print V _DFF_IP1_01_|3|MID_SHUNT
.print V _PG1_01_|_AND_G|B1
.print DEVP BSPL_IG0_0_|1|1
.print DEVP BSPL_IG0_0_|2|1
.print DEVP BSPL_IG0_0_|A|1
.print DEVP BSPL_IG0_0_|B|1
.print DEVP BSPL_IP1_0_|1|1
.print DEVP BSPL_IP1_0_|2|1
.print DEVP BSPL_IP1_0_|A|1
.print DEVP BSPL_IP1_0_|B|1
.print DEVP BSPL_IG2_0_|1|1
.print DEVP BSPL_IG2_0_|2|1
.print DEVP BSPL_IG2_0_|A|1
.print DEVP BSPL_IG2_0_|B|1
.print DEVP BSPL_IP3_0_|1|1
.print DEVP BSPL_IP3_0_|2|1
.print DEVP BSPL_IP3_0_|A|1
.print DEVP BSPL_IP3_0_|B|1
.print DEVP B_DFF_IP1_01_|1|1
.print DEVP B_DFF_IP1_01_|23|1
.print DEVP B_DFF_IP1_01_|3|1
.print DEVP B_DFF_IP1_01_|4|1
.print DEVP B_DFF_IP1_01_|T|1
.print DEVP B_DFF_IP1_01_|45|1
.print DEVP B_DFF_IP1_01_|6|1
.print DEVP B_DFF_IP2_01_|1|1
.print DEVP B_DFF_IP2_01_|23|1
.print DEVP B_DFF_IP2_01_|3|1
.print DEVP B_DFF_IP2_01_|4|1
.print DEVP B_DFF_IP2_01_|T|1
.print DEVP B_DFF_IP2_01_|45|1
.print DEVP B_DFF_IP2_01_|6|1
.print DEVP B_DFF_IP3_01_|1|1
.print DEVP B_DFF_IP3_01_|23|1
.print DEVP B_DFF_IP3_01_|3|1
.print DEVP B_DFF_IP3_01_|4|1
.print DEVP B_DFF_IP3_01_|T|1
.print DEVP B_DFF_IP3_01_|45|1
.print DEVP B_DFF_IP3_01_|6|1
