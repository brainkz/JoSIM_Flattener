*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=5e-11
.PARAM TCLOCK=1e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.1E-12 1E-09
L1 Q0 Q1  PHI0/(4*IC*IC0)
ROUT Q 0  1
IT1|T 0 CLK  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 1.47e-10 0 1.5e-10 0.0007 1.53e-10 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 3.47e-10 0 3.5e-10 0.0007 3.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 5.47e-10 0 5.5e-10 0.0007 5.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 7.47e-10 0 7.5e-10 0.0007 7.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 9.47e-10 0 9.5e-10 0.0007 9.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.147e-09 0 1.15e-09 0.0007 1.153e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.347e-09 0 1.35e-09 0.0007 1.353e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.547e-09 0 1.55e-09 0.0007 1.553e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.747e-09 0 1.75e-09 0.0007 1.753e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 1.947e-09 0 1.95e-09 0.0007 1.953e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.147e-09 0 2.15e-09 0.0007 2.153e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.347e-09 0 2.35e-09 0.0007 2.353e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.547e-09 0 2.55e-09 0.0007 2.553e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.747e-09 0 2.75e-09 0.0007 2.753e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 2.947e-09 0 2.95e-09 0.0007 2.953e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.147e-09 0 3.15e-09 0.0007 3.153e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.347e-09 0 3.35e-09 0.0007 3.353e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.547e-09 0 3.55e-09 0.0007 3.553e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.747e-09 0 3.75e-09 0.0007 3.753e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 3.947e-09 0 3.95e-09 0.0007 3.953e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.147e-09 0 4.15e-09 0.0007 4.153e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.347e-09 0 4.35e-09 0.0007 4.353e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.547e-09 0 4.55e-09 0.0007 4.553e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.747e-09 0 4.75e-09 0.0007 4.753e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 4.947e-09 0 4.95e-09 0.0007 4.953e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.147e-09 0 5.15e-09 0.0007 5.153e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.347e-09 0 5.35e-09 0.0007 5.353e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.547e-09 0 5.55e-09 0.0007 5.553e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.747e-09 0 5.75e-09 0.0007 5.753e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 5.947e-09 0 5.95e-09 0.0007 5.953e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.147e-09 0 6.15e-09 0.0007 6.153e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.347e-09 0 6.35e-09 0.0007 6.353e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.547e-09 0 6.55e-09 0.0007 6.553e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.747e-09 0 6.75e-09 0.0007 6.753e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 6.947e-09 0 6.95e-09 0.0007 6.953e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.147e-09 0 7.15e-09 0.0007 7.153e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.347e-09 0 7.35e-09 0.0007 7.353e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.547e-09 0 7.55e-09 0.0007 7.553e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.747e-09 0 7.75e-09 0.0007 7.753e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 7.947e-09 0 7.95e-09 0.0007 7.953e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.147e-09 0 8.15e-09 0.0007 8.153e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.347e-09 0 8.35e-09 0.0007 8.353e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.547e-09 0 8.55e-09 0.0007 8.553e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.747e-09 0 8.75e-09 0.0007 8.753e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 8.947e-09 0 8.95e-09 0.0007 8.953e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.147e-09 0 9.15e-09 0.0007 9.153e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.347e-09 0 9.35e-09 0.0007 9.353e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.547e-09 0 9.55e-09 0.0007 9.553e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.747e-09 0 9.75e-09 0.0007 9.753e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 9.947e-09 0 9.95e-09 0.0007 9.953e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0147e-08 0 1.015e-08 0.0007 1.0153e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0347e-08 0 1.035e-08 0.0007 1.0353e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0547e-08 0 1.055e-08 0.0007 1.0553e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0747e-08 0 1.075e-08 0.0007 1.0753e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.0947e-08 0 1.095e-08 0.0007 1.0953e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1147e-08 0 1.115e-08 0.0007 1.1153e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1347e-08 0 1.135e-08 0.0007 1.1353e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1547e-08 0 1.155e-08 0.0007 1.1553e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1747e-08 0 1.175e-08 0.0007 1.1753e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.1947e-08 0 1.195e-08 0.0007 1.1953e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2147e-08 0 1.215e-08 0.0007 1.2153e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2347e-08 0 1.235e-08 0.0007 1.2353e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2547e-08 0 1.255e-08 0.0007 1.2553e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2747e-08 0 1.275e-08 0.0007 1.2753e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.2947e-08 0 1.295e-08 0.0007 1.2953e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3147e-08 0 1.315e-08 0.0007 1.3153e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3347e-08 0 1.335e-08 0.0007 1.3353e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3547e-08 0 1.355e-08 0.0007 1.3553e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3747e-08 0 1.375e-08 0.0007 1.3753e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.3947e-08 0 1.395e-08 0.0007 1.3953e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4147e-08 0 1.415e-08 0.0007 1.4153e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4347e-08 0 1.435e-08 0.0007 1.4353e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4547e-08 0 1.455e-08 0.0007 1.4553e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4747e-08 0 1.475e-08 0.0007 1.4753e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.4947e-08 0 1.495e-08 0.0007 1.4953e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5147e-08 0 1.515e-08 0.0007 1.5153e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5347e-08 0 1.535e-08 0.0007 1.5353e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5547e-08 0 1.555e-08 0.0007 1.5553e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5747e-08 0 1.575e-08 0.0007 1.5753e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.5947e-08 0 1.595e-08 0.0007 1.5953e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6147e-08 0 1.615e-08 0.0007 1.6153e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6347e-08 0 1.635e-08 0.0007 1.6353e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6547e-08 0 1.655e-08 0.0007 1.6553e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6747e-08 0 1.675e-08 0.0007 1.6753e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.6947e-08 0 1.695e-08 0.0007 1.6953e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7147e-08 0 1.715e-08 0.0007 1.7153e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7347e-08 0 1.735e-08 0.0007 1.7353e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7547e-08 0 1.755e-08 0.0007 1.7553e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7747e-08 0 1.775e-08 0.0007 1.7753e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.7947e-08 0 1.795e-08 0.0007 1.7953e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8147e-08 0 1.815e-08 0.0007 1.8153e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8347e-08 0 1.835e-08 0.0007 1.8353e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8547e-08 0 1.855e-08 0.0007 1.8553e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8747e-08 0 1.875e-08 0.0007 1.8753e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.8947e-08 0 1.895e-08 0.0007 1.8953e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9147e-08 0 1.915e-08 0.0007 1.9153e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9347e-08 0 1.935e-08 0.0007 1.9353e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9547e-08 0 1.955e-08 0.0007 1.9553e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9747e-08 0 1.975e-08 0.0007 1.9753e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 1.9947e-08 0 1.995e-08 0.0007 1.9953e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0147e-08 0 2.015e-08 0.0007 2.0153e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0347e-08 0 2.035e-08 0.0007 2.0353e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0547e-08 0 2.055e-08 0.0007 2.0553e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0747e-08 0 2.075e-08 0.0007 2.0753e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.0947e-08 0 2.095e-08 0.0007 2.0953e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1147e-08 0 2.115e-08 0.0007 2.1153e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1347e-08 0 2.135e-08 0.0007 2.1353e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1547e-08 0 2.155e-08 0.0007 2.1553e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1747e-08 0 2.175e-08 0.0007 2.1753e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.1947e-08 0 2.195e-08 0.0007 2.1953e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2147e-08 0 2.215e-08 0.0007 2.2153e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2347e-08 0 2.235e-08 0.0007 2.2353e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2547e-08 0 2.255e-08 0.0007 2.2553e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2747e-08 0 2.275e-08 0.0007 2.2753e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.2947e-08 0 2.295e-08 0.0007 2.2953e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3147e-08 0 2.315e-08 0.0007 2.3153e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3347e-08 0 2.335e-08 0.0007 2.3353e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3547e-08 0 2.355e-08 0.0007 2.3553e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3747e-08 0 2.375e-08 0.0007 2.3753e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.3947e-08 0 2.395e-08 0.0007 2.3953e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4147e-08 0 2.415e-08 0.0007 2.4153e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4347e-08 0 2.435e-08 0.0007 2.4353e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4547e-08 0 2.455e-08 0.0007 2.4553e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4747e-08 0 2.475e-08 0.0007 2.4753e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.4947e-08 0 2.495e-08 0.0007 2.4953e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5147e-08 0 2.515e-08 0.0007 2.5153e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5347e-08 0 2.535e-08 0.0007 2.5353e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5547e-08 0 2.555e-08 0.0007 2.5553e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5747e-08 0 2.575e-08 0.0007 2.5753e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.5947e-08 0 2.595e-08 0.0007 2.5953e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6147e-08 0 2.615e-08 0.0007 2.6153e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6347e-08 0 2.635e-08 0.0007 2.6353e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6547e-08 0 2.655e-08 0.0007 2.6553e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6747e-08 0 2.675e-08 0.0007 2.6753e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.6947e-08 0 2.695e-08 0.0007 2.6953e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7147e-08 0 2.715e-08 0.0007 2.7153e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7347e-08 0 2.735e-08 0.0007 2.7353e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7547e-08 0 2.755e-08 0.0007 2.7553e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7747e-08 0 2.775e-08 0.0007 2.7753e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.7947e-08 0 2.795e-08 0.0007 2.7953e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8147e-08 0 2.815e-08 0.0007 2.8153e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8347e-08 0 2.835e-08 0.0007 2.8353e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8547e-08 0 2.855e-08 0.0007 2.8553e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8747e-08 0 2.875e-08 0.0007 2.8753e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.8947e-08 0 2.895e-08 0.0007 2.8953e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9147e-08 0 2.915e-08 0.0007 2.9153e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9347e-08 0 2.935e-08 0.0007 2.9353e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9547e-08 0 2.955e-08 0.0007 2.9553e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9747e-08 0 2.975e-08 0.0007 2.9753e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 2.9947e-08 0 2.995e-08 0.0007 2.9953e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0147e-08 0 3.015e-08 0.0007 3.0153e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0347e-08 0 3.035e-08 0.0007 3.0353e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0547e-08 0 3.055e-08 0.0007 3.0553e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0747e-08 0 3.075e-08 0.0007 3.0753e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.0947e-08 0 3.095e-08 0.0007 3.0953e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1147e-08 0 3.115e-08 0.0007 3.1153e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1347e-08 0 3.135e-08 0.0007 3.1353e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1547e-08 0 3.155e-08 0.0007 3.1553e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1747e-08 0 3.175e-08 0.0007 3.1753e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.1947e-08 0 3.195e-08 0.0007 3.1953e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2147e-08 0 3.215e-08 0.0007 3.2153e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2347e-08 0 3.235e-08 0.0007 3.2353e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2547e-08 0 3.255e-08 0.0007 3.2553e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2747e-08 0 3.275e-08 0.0007 3.2753e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.2947e-08 0 3.295e-08 0.0007 3.2953e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3147e-08 0 3.315e-08 0.0007 3.3153e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3347e-08 0 3.335e-08 0.0007 3.3353e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3547e-08 0 3.355e-08 0.0007 3.3553e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3747e-08 0 3.375e-08 0.0007 3.3753e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.3947e-08 0 3.395e-08 0.0007 3.3953e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4147e-08 0 3.415e-08 0.0007 3.4153e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4347e-08 0 3.435e-08 0.0007 3.4353e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4547e-08 0 3.455e-08 0.0007 3.4553e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4747e-08 0 3.475e-08 0.0007 3.4753e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.4947e-08 0 3.495e-08 0.0007 3.4953e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5147e-08 0 3.515e-08 0.0007 3.5153e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5347e-08 0 3.535e-08 0.0007 3.5353e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5547e-08 0 3.555e-08 0.0007 3.5553e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5747e-08 0 3.575e-08 0.0007 3.5753e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.5947e-08 0 3.595e-08 0.0007 3.5953e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6147e-08 0 3.615e-08 0.0007 3.6153e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6347e-08 0 3.635e-08 0.0007 3.6353e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6547e-08 0 3.655e-08 0.0007 3.6553e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6747e-08 0 3.675e-08 0.0007 3.6753e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.6947e-08 0 3.695e-08 0.0007 3.6953e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7147e-08 0 3.715e-08 0.0007 3.7153e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7347e-08 0 3.735e-08 0.0007 3.7353e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7547e-08 0 3.755e-08 0.0007 3.7553e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7747e-08 0 3.775e-08 0.0007 3.7753e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.7947e-08 0 3.795e-08 0.0007 3.7953e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8147e-08 0 3.815e-08 0.0007 3.8153e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8347e-08 0 3.835e-08 0.0007 3.8353e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8547e-08 0 3.855e-08 0.0007 3.8553e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8747e-08 0 3.875e-08 0.0007 3.8753e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.8947e-08 0 3.895e-08 0.0007 3.8953e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9147e-08 0 3.915e-08 0.0007 3.9153e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9347e-08 0 3.935e-08 0.0007 3.9353e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9547e-08 0 3.955e-08 0.0007 3.9553e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9747e-08 0 3.975e-08 0.0007 3.9753e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0)
L_TFF|A1 CLK _TFF|A1  2.067833848e-12
L_TFF|JCT _TFF|A1 _TFF|JCT  2.067833848e-12
L_TFF|U1 _TFF|JCT _TFF|U1  4.135667696e-12
L_TFF|UQ _TFF|U2 _TFF|Q1  2.067833848e-12
L_TFF|L1 _TFF|JCT _TFF|L1  8.271335392e-12
L_TFF|L2 _TFF|L2 _TFF|L3  2.067833848e-12
L_TFF|LQ _TFF|L3 _TFF|Q1  2.2746172328000002e-11
L_TFF|Q _TFF|Q1 Q0  4.135667696e-12
B_BUF|1 _BUF|1 _BUF|2 JJMIT AREA=2.5
B_BUF|2 _BUF|4 _BUF|5 JJMIT AREA=2.5
B_BUF|3 _BUF|7 _BUF|8 JJMIT AREA=2.5
B_BUF|4 _BUF|10 _BUF|11 JJMIT AREA=2.5
I_BUF|B1 0 _BUF|3  PWL(0 0 5e-12 0.000175)
I_BUF|B2 0 _BUF|6  PWL(0 0 5e-12 0.0002375)
I_BUF|B3 0 _BUF|9  PWL(0 0 5e-12 0.0002375)
I_BUF|B4 0 _BUF|12  PWL(0 0 5e-12 0.000175)
L_BUF|1 Q1 _BUF|1  2.067833848e-12
L_BUF|2 _BUF|1 _BUF|4  4.135667696e-12
L_BUF|3 _BUF|4 _BUF|7  4.135667696e-12
L_BUF|4 _BUF|7 _BUF|10  4.135667696e-12
L_BUF|5 _BUF|10 Q  2.067833848e-12
L_BUF|P1 _BUF|2 0  5e-13
L_BUF|P2 _BUF|5 0  5e-13
L_BUF|P3 _BUF|8 0  5e-13
L_BUF|P4 _BUF|11 0  5e-13
L_BUF|B1 _BUF|1 _BUF|3  2e-12
L_BUF|B2 _BUF|4 _BUF|6  2e-12
L_BUF|B3 _BUF|7 _BUF|9  2e-12
L_BUF|B4 _BUF|10 _BUF|12  2e-12
R_BUF|B1 _BUF|1 _BUF|101  2.7439617672
R_BUF|B2 _BUF|4 _BUF|104  2.7439617672
R_BUF|B3 _BUF|7 _BUF|107  2.7439617672
R_BUF|B4 _BUF|10 _BUF|110  2.7439617672
L_BUF|RB1 _BUF|101 0  2.050338398468e-12
L_BUF|RB2 _BUF|104 0  2.050338398468e-12
L_BUF|RB3 _BUF|107 0  2.050338398468e-12
L_BUF|RB4 _BUF|110 0  2.050338398468e-12
L_TFF|I_A1|B _TFF|A1 _TFF|I_A1|MID  2e-12
I_TFF|I_A1|B 0 _TFF|I_A1|MID  PWL(0 0 5e-12 0.0003675)
L_TFF|I_L3|B _TFF|L3 _TFF|I_L3|MID  2e-12
I_TFF|I_L3|B 0 _TFF|I_L3|MID  PWL(0 0 5e-12 3.5e-05)
L_TFF|I_U2|B _TFF|U2 _TFF|I_U2|MID  2e-12
I_TFF|I_U2|B _TFF|I_U2|MID 0  PWL(0 0 5e-12 8.75e-05)
B_TFF|A1|1 _TFF|A1 _TFF|A1|MID_SERIES JJMIT AREA=2.5
L_TFF|A1|P _TFF|A1|MID_SERIES 0  2e-13
R_TFF|A1|B _TFF|A1 _TFF|A1|MID_SHUNT  2.7439617672
L_TFF|A1|RB _TFF|A1|MID_SHUNT 0  1.550338398468e-12
B_TFF|U1|1 _TFF|U1 _TFF|U1|MID_SERIES JJMIT AREA=2.5
L_TFF|U1|P _TFF|U1|MID_SERIES _TFF|U2  2e-13
R_TFF|U1|B _TFF|U1 _TFF|U1|MID_SHUNT  2.7439617672
L_TFF|U1|RB _TFF|U1|MID_SHUNT _TFF|U2  1.550338398468e-12
B_TFF|U2|1 _TFF|U2 _TFF|U2|MID_SERIES JJMIT AREA=2.5
L_TFF|U2|P _TFF|U2|MID_SERIES 0  2e-13
R_TFF|U2|B _TFF|U2 _TFF|U2|MID_SHUNT  2.7439617672
L_TFF|U2|RB _TFF|U2|MID_SHUNT 0  1.550338398468e-12
B_TFF|L1|1 _TFF|L1 _TFF|L1|MID_SERIES JJMIT AREA=2.5
L_TFF|L1|P _TFF|L1|MID_SERIES _TFF|L2  2e-13
R_TFF|L1|B _TFF|L1 _TFF|L1|MID_SHUNT  2.7439617672
L_TFF|L1|RB _TFF|L1|MID_SHUNT _TFF|L2  1.550338398468e-12
B_TFF|L2|1 _TFF|L2 _TFF|L2|MID_SERIES JJMIT AREA=2.5
L_TFF|L2|P _TFF|L2|MID_SERIES 0  2e-13
R_TFF|L2|B _TFF|L2 _TFF|L2|MID_SHUNT  2.7439617672
L_TFF|L2|RB _TFF|L2|MID_SHUNT 0  1.550338398468e-12
.print DEVI L1
.print DEVI ROUT
.print DEVI IT1|T
.print DEVI L_TFF|A1
.print DEVI L_TFF|JCT
.print DEVI L_TFF|U1
.print DEVI L_TFF|UQ
.print DEVI L_TFF|L1
.print DEVI L_TFF|L2
.print DEVI L_TFF|LQ
.print DEVI L_TFF|Q
.print DEVI B_BUF|1
.print DEVI B_BUF|2
.print DEVI B_BUF|3
.print DEVI B_BUF|4
.print DEVI I_BUF|B1
.print DEVI I_BUF|B2
.print DEVI I_BUF|B3
.print DEVI I_BUF|B4
.print DEVI L_BUF|1
.print DEVI L_BUF|2
.print DEVI L_BUF|3
.print DEVI L_BUF|4
.print DEVI L_BUF|5
.print DEVI L_BUF|P1
.print DEVI L_BUF|P2
.print DEVI L_BUF|P3
.print DEVI L_BUF|P4
.print DEVI L_BUF|B1
.print DEVI L_BUF|B2
.print DEVI L_BUF|B3
.print DEVI L_BUF|B4
.print DEVI R_BUF|B1
.print DEVI R_BUF|B2
.print DEVI R_BUF|B3
.print DEVI R_BUF|B4
.print DEVI L_BUF|RB1
.print DEVI L_BUF|RB2
.print DEVI L_BUF|RB3
.print DEVI L_BUF|RB4
.print V _BUF|9
.print V _TFF|L2
.print V CLK
.print V _BUF|4
.print V _BUF|110
.print V _BUF|107
.print V _BUF|10
.print V _BUF|11
.print V _TFF|Q1
.print V Q0
.print V _TFF|A1
.print V _BUF|6
.print V _BUF|5
.print V _TFF|JCT
.print V _BUF|12
.print V _BUF|3
.print V _BUF|1
.print V _BUF|7
.print V _BUF|101
.print V _BUF|104
.print V _TFF|U2
.print V Q
.print V Q1
.print V _TFF|L1
.print V _TFF|U1
.print V _BUF|2
.print V _TFF|L3
.print V _BUF|8
.print DEVP B_BUF|1
.print DEVP B_BUF|2
.print DEVP B_BUF|3
.print DEVP B_BUF|4
.print DEVP B_TFF|A1|1
.print DEVP B_TFF|U1|1
.print DEVP B_TFF|U2|1
.print DEVP B_TFF|L1|1
.print DEVP B_TFF|L2|1
