*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=1e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.1E-12 4E-10
ROUT A_AND_B 0  1
IDATA_A1|A 0 A  PWL(0 0 1.52e-10 0 1.55e-10 0.0005 1.58e-10 0 2.52e-10 0 2.55e-10 0.0005 2.58e-10 0 3.52e-10 0 3.55e-10 0.0005 3.58e-10 0 4.52e-10 0 4.55e-10 0.0005 4.58e-10 0 5.52e-10 0 5.55e-10 0.0005 5.58e-10 0 6.52e-10 0 6.55e-10 0.0005 6.58e-10 0 7.52e-10 0 7.55e-10 0.0005 7.58e-10 0 8.52e-10 0 8.55e-10 0.0005 8.58e-10 0 9.52e-10 0 9.55e-10 0.0005 9.58e-10 0 1.052e-09 0 1.055e-09 0.0005 1.058e-09 0 1.152e-09 0 1.155e-09 0.0005 1.158e-09 0 1.252e-09 0 1.255e-09 0.0005 1.258e-09 0 1.352e-09 0 1.355e-09 0.0005 1.358e-09 0 1.452e-09 0 1.455e-09 0.0005 1.458e-09 0 1.552e-09 0 1.555e-09 0.0005 1.558e-09 0 1.652e-09 0 1.655e-09 0.0005 1.658e-09 0 1.752e-09 0 1.755e-09 0.0005 1.758e-09 0 1.852e-09 0 1.855e-09 0.0005 1.858e-09 0 1.952e-09 0 1.955e-09 0.0005 1.958e-09 0)
IDATA_B1|B 0 B  PWL(0 0 2.02e-10 0 2.05e-10 0.0005 2.08e-10 0 2.52e-10 0 2.55e-10 0.0005 2.58e-10 0 4.02e-10 0 4.05e-10 0.0005 4.08e-10 0 4.52e-10 0 4.55e-10 0.0005 4.58e-10 0 6.02e-10 0 6.05e-10 0.0005 6.08e-10 0 6.52e-10 0 6.55e-10 0.0005 6.58e-10 0 8.02e-10 0 8.05e-10 0.0005 8.08e-10 0 8.52e-10 0 8.55e-10 0.0005 8.58e-10 0 1.002e-09 0 1.005e-09 0.0005 1.008e-09 0 1.052e-09 0 1.055e-09 0.0005 1.058e-09 0 1.202e-09 0 1.205e-09 0.0005 1.208e-09 0 1.252e-09 0 1.255e-09 0.0005 1.258e-09 0 1.402e-09 0 1.405e-09 0.0005 1.408e-09 0 1.452e-09 0 1.455e-09 0.0005 1.458e-09 0 1.602e-09 0 1.605e-09 0.0005 1.608e-09 0 1.652e-09 0 1.655e-09 0.0005 1.658e-09 0 1.802e-09 0 1.805e-09 0.0005 1.808e-09 0 1.852e-09 0 1.855e-09 0.0005 1.858e-09 0 2.002e-09 0 2.005e-09 0.0005 2.008e-09 0)
L_JTL1|1 B _JTL1|1  2.067833848e-12
L_JTL1|2 _JTL1|1 _JTL1|4  2.067833848e-12
L_JTL1|3 _JTL1|4 _JTL1|6  2.067833848e-12
L_JTL1|4 _JTL1|6 1  2.067833848e-12
L_JTL2|1 1 _JTL2|1  2.067833848e-12
L_JTL2|2 _JTL2|1 _JTL2|4  2.067833848e-12
L_JTL2|3 _JTL2|4 _JTL2|6  2.067833848e-12
L_JTL2|4 _JTL2|6 2  2.067833848e-12
L_JTL3|1 2 _JTL3|1  2.067833848e-12
L_JTL3|2 _JTL3|1 _JTL3|4  2.067833848e-12
L_JTL3|3 _JTL3|4 _JTL3|6  2.067833848e-12
L_JTL3|4 _JTL3|6 3  2.067833848e-12
L_JTL5|1 3 _JTL5|1  2.067833848e-12
L_JTL5|2 _JTL5|1 _JTL5|4  2.067833848e-12
L_JTL5|3 _JTL5|4 _JTL5|6  2.067833848e-12
L_JTL5|4 _JTL5|6 B1  2.067833848e-12
L_MERGE|A1 A _MERGE|A1  2.067833848e-12
L_MERGE|A2 _MERGE|A1 _MERGE|A2  4.135667696e-12
L_MERGE|A3 _MERGE|A3 _MERGE|Q3  1.2e-12
L_MERGE|B1 B1 _MERGE|B1  2.067833848e-12
L_MERGE|B2 _MERGE|B1 _MERGE|B2  4.135667696e-12
L_MERGE|B3 _MERGE|B3 _MERGE|Q3  1.2e-12
L_MERGE|Q3 _MERGE|Q3 _MERGE|Q2  4.135667696e-12
L_MERGE|Q2 _MERGE|Q2 _MERGE|Q1  4.135667696e-12
L_MERGE|Q1 _MERGE|Q1 A_AND_B  2.067833848e-12
B_JTL1|1|1 _JTL1|1 _JTL1|1|MID_SERIES JJMIT AREA=2.5
L_JTL1|1|P _JTL1|1|MID_SERIES 0  2e-13
R_JTL1|1|B _JTL1|1 _JTL1|1|MID_SHUNT  2.7439617672
L_JTL1|1|RB _JTL1|1|MID_SHUNT 0  1.750338398468e-12
L_JTL1|B|B _JTL1|4 _JTL1|B|MID  2e-12
I_JTL1|B|B 0 _JTL1|B|MID  0.0005
B_JTL1|2|1 _JTL1|6 _JTL1|2|MID_SERIES JJMIT AREA=2.5
L_JTL1|2|P _JTL1|2|MID_SERIES 0  2e-13
R_JTL1|2|B _JTL1|6 _JTL1|2|MID_SHUNT  2.7439617672
L_JTL1|2|RB _JTL1|2|MID_SHUNT 0  1.750338398468e-12
B_JTL2|1|1 _JTL2|1 _JTL2|1|MID_SERIES JJMIT AREA=2.5
L_JTL2|1|P _JTL2|1|MID_SERIES 0  2e-13
R_JTL2|1|B _JTL2|1 _JTL2|1|MID_SHUNT  2.7439617672
L_JTL2|1|RB _JTL2|1|MID_SHUNT 0  1.750338398468e-12
L_JTL2|B|B _JTL2|4 _JTL2|B|MID  2e-12
I_JTL2|B|B 0 _JTL2|B|MID  0.0005
B_JTL2|2|1 _JTL2|6 _JTL2|2|MID_SERIES JJMIT AREA=2.5
L_JTL2|2|P _JTL2|2|MID_SERIES 0  2e-13
R_JTL2|2|B _JTL2|6 _JTL2|2|MID_SHUNT  2.7439617672
L_JTL2|2|RB _JTL2|2|MID_SHUNT 0  1.750338398468e-12
B_JTL3|1|1 _JTL3|1 _JTL3|1|MID_SERIES JJMIT AREA=2.5
L_JTL3|1|P _JTL3|1|MID_SERIES 0  2e-13
R_JTL3|1|B _JTL3|1 _JTL3|1|MID_SHUNT  2.7439617672
L_JTL3|1|RB _JTL3|1|MID_SHUNT 0  1.750338398468e-12
L_JTL3|B|B _JTL3|4 _JTL3|B|MID  2e-12
I_JTL3|B|B 0 _JTL3|B|MID  0.0005
B_JTL3|2|1 _JTL3|6 _JTL3|2|MID_SERIES JJMIT AREA=2.5
L_JTL3|2|P _JTL3|2|MID_SERIES 0  2e-13
R_JTL3|2|B _JTL3|6 _JTL3|2|MID_SHUNT  2.7439617672
L_JTL3|2|RB _JTL3|2|MID_SHUNT 0  1.750338398468e-12
B_JTL5|1|1 _JTL5|1 _JTL5|1|MID_SERIES JJMIT AREA=2.5
L_JTL5|1|P _JTL5|1|MID_SERIES 0  2e-13
R_JTL5|1|B _JTL5|1 _JTL5|1|MID_SHUNT  2.7439617672
L_JTL5|1|RB _JTL5|1|MID_SHUNT 0  1.750338398468e-12
L_JTL5|B|B _JTL5|4 _JTL5|B|MID  2e-12
I_JTL5|B|B 0 _JTL5|B|MID  0.0005
B_JTL5|2|1 _JTL5|6 _JTL5|2|MID_SERIES JJMIT AREA=2.5
L_JTL5|2|P _JTL5|2|MID_SERIES 0  2e-13
R_JTL5|2|B _JTL5|6 _JTL5|2|MID_SHUNT  2.7439617672
L_JTL5|2|RB _JTL5|2|MID_SHUNT 0  1.750338398468e-12
L_MERGE|I_A1|B _MERGE|A1 _MERGE|I_A1|MID  2e-12
I_MERGE|I_A1|B 0 _MERGE|I_A1|MID  0.000175
L_MERGE|I_B1|B _MERGE|B1 _MERGE|I_B1|MID  2e-12
I_MERGE|I_B1|B 0 _MERGE|I_B1|MID  0.000175
L_MERGE|I_Q3|B _MERGE|Q3 _MERGE|I_Q3|MID  2e-12
I_MERGE|I_Q3|B 0 _MERGE|I_Q3|MID  7.5e-05
L_MERGE|I_Q2|B _MERGE|Q2 _MERGE|I_Q2|MID  2e-12
I_MERGE|I_Q2|B 0 _MERGE|I_Q2|MID  0.000175
L_MERGE|I_Q1|B _MERGE|Q1 _MERGE|I_Q1|MID  2e-12
I_MERGE|I_Q1|B 0 _MERGE|I_Q1|MID  0.000175
B_MERGE|A1|1 _MERGE|A1 _MERGE|A1|MID_SERIES JJMIT AREA=2.5
L_MERGE|A1|P _MERGE|A1|MID_SERIES 0  2e-13
R_MERGE|A1|B _MERGE|A1 _MERGE|A1|MID_SHUNT  2.7439617672
L_MERGE|A1|RB _MERGE|A1|MID_SHUNT 0  1.550338398468e-12
B_MERGE|A2|1 _MERGE|A2 _MERGE|A2|MID_SERIES JJMIT AREA=2.5
L_MERGE|A2|P _MERGE|A2|MID_SERIES 0  2e-13
R_MERGE|A2|B _MERGE|A2 _MERGE|A2|MID_SHUNT  2.7439617672
L_MERGE|A2|RB _MERGE|A2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|A12|1 _MERGE|A2 _MERGE|A3 JJMIT AREA=1.7857142857142858
R_MERGE|A12|B _MERGE|A2 _MERGE|A12|MID_SHUNT  3.84154647408
L_MERGE|A12|RB _MERGE|A12|MID_SHUNT _MERGE|A3  2.1704737578552e-12
B_MERGE|B1|1 _MERGE|B1 _MERGE|B1|MID_SERIES JJMIT AREA=2.5
L_MERGE|B1|P _MERGE|B1|MID_SERIES 0  2e-13
R_MERGE|B1|B _MERGE|B1 _MERGE|B1|MID_SHUNT  2.7439617672
L_MERGE|B1|RB _MERGE|B1|MID_SHUNT 0  1.550338398468e-12
B_MERGE|B2|1 _MERGE|B2 _MERGE|B2|MID_SERIES JJMIT AREA=2.5
L_MERGE|B2|P _MERGE|B2|MID_SERIES 0  2e-13
R_MERGE|B2|B _MERGE|B2 _MERGE|B2|MID_SHUNT  2.7439617672
L_MERGE|B2|RB _MERGE|B2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|B12|1 _MERGE|B2 _MERGE|B3 JJMIT AREA=1.7857142857142858
R_MERGE|B12|B _MERGE|B2 _MERGE|B12|MID_SHUNT  3.84154647408
L_MERGE|B12|RB _MERGE|B12|MID_SHUNT _MERGE|B3  2.1704737578552e-12
B_MERGE|Q2|1 _MERGE|Q2 _MERGE|Q2|MID_SERIES JJMIT AREA=2.5
L_MERGE|Q2|P _MERGE|Q2|MID_SERIES 0  2e-13
R_MERGE|Q2|B _MERGE|Q2 _MERGE|Q2|MID_SHUNT  2.7439617672
L_MERGE|Q2|RB _MERGE|Q2|MID_SHUNT 0  1.550338398468e-12
B_MERGE|Q1|1 _MERGE|Q1 _MERGE|Q1|MID_SERIES JJMIT AREA=2.5
L_MERGE|Q1|P _MERGE|Q1|MID_SERIES 0  2e-13
R_MERGE|Q1|B _MERGE|Q1 _MERGE|Q1|MID_SHUNT  2.7439617672
L_MERGE|Q1|RB _MERGE|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI ROUT
.print DEVI IDATA_A1|A
.print DEVI IDATA_B1|B
.print DEVI L_JTL1|1
.print DEVI L_JTL1|2
.print DEVI L_JTL1|3
.print DEVI L_JTL1|4
.print DEVI L_JTL2|1
.print DEVI L_JTL2|2
.print DEVI L_JTL2|3
.print DEVI L_JTL2|4
.print DEVI L_JTL3|1
.print DEVI L_JTL3|2
.print DEVI L_JTL3|3
.print DEVI L_JTL3|4
.print DEVI L_JTL5|1
.print DEVI L_JTL5|2
.print DEVI L_JTL5|3
.print DEVI L_JTL5|4
.print DEVI L_MERGE|A1
.print DEVI L_MERGE|A2
.print DEVI L_MERGE|A3
.print DEVI L_MERGE|B1
.print DEVI L_MERGE|B2
.print DEVI L_MERGE|B3
.print DEVI L_MERGE|Q3
.print DEVI L_MERGE|Q2
.print DEVI L_MERGE|Q1
.print DEVI B_JTL1|1|1
.print DEVI L_JTL1|1|P
.print DEVI R_JTL1|1|B
.print DEVI L_JTL1|1|RB
.print DEVI L_JTL1|B|B
.print DEVI I_JTL1|B|B
.print DEVI B_JTL1|2|1
.print DEVI L_JTL1|2|P
.print DEVI R_JTL1|2|B
.print DEVI L_JTL1|2|RB
.print DEVI B_JTL2|1|1
.print DEVI L_JTL2|1|P
.print DEVI R_JTL2|1|B
.print DEVI L_JTL2|1|RB
.print DEVI L_JTL2|B|B
.print DEVI I_JTL2|B|B
.print DEVI B_JTL2|2|1
.print DEVI L_JTL2|2|P
.print DEVI R_JTL2|2|B
.print DEVI L_JTL2|2|RB
.print DEVI B_JTL3|1|1
.print DEVI L_JTL3|1|P
.print DEVI R_JTL3|1|B
.print DEVI L_JTL3|1|RB
.print DEVI L_JTL3|B|B
.print DEVI I_JTL3|B|B
.print DEVI B_JTL3|2|1
.print DEVI L_JTL3|2|P
.print DEVI R_JTL3|2|B
.print DEVI L_JTL3|2|RB
.print DEVI B_JTL5|1|1
.print DEVI L_JTL5|1|P
.print DEVI R_JTL5|1|B
.print DEVI L_JTL5|1|RB
.print DEVI L_JTL5|B|B
.print DEVI I_JTL5|B|B
.print DEVI B_JTL5|2|1
.print DEVI L_JTL5|2|P
.print DEVI R_JTL5|2|B
.print DEVI L_JTL5|2|RB
.print DEVI L_MERGE|I_A1|B
.print DEVI I_MERGE|I_A1|B
.print DEVI L_MERGE|I_B1|B
.print DEVI I_MERGE|I_B1|B
.print DEVI L_MERGE|I_Q3|B
.print DEVI I_MERGE|I_Q3|B
.print DEVI L_MERGE|I_Q2|B
.print DEVI I_MERGE|I_Q2|B
.print DEVI L_MERGE|I_Q1|B
.print DEVI I_MERGE|I_Q1|B
.print DEVI B_MERGE|A1|1
.print DEVI L_MERGE|A1|P
.print DEVI R_MERGE|A1|B
.print DEVI L_MERGE|A1|RB
.print DEVI B_MERGE|A2|1
.print DEVI L_MERGE|A2|P
.print DEVI R_MERGE|A2|B
.print DEVI L_MERGE|A2|RB
.print DEVI B_MERGE|A12|1
.print DEVI R_MERGE|A12|B
.print DEVI L_MERGE|A12|RB
.print DEVI B_MERGE|B1|1
.print DEVI L_MERGE|B1|P
.print DEVI R_MERGE|B1|B
.print DEVI L_MERGE|B1|RB
.print DEVI B_MERGE|B2|1
.print DEVI L_MERGE|B2|P
.print DEVI R_MERGE|B2|B
.print DEVI L_MERGE|B2|RB
.print DEVI B_MERGE|B12|1
.print DEVI R_MERGE|B12|B
.print DEVI L_MERGE|B12|RB
.print DEVI B_MERGE|Q2|1
.print DEVI L_MERGE|Q2|P
.print DEVI R_MERGE|Q2|B
.print DEVI L_MERGE|Q2|RB
.print DEVI B_MERGE|Q1|1
.print DEVI L_MERGE|Q1|P
.print DEVI R_MERGE|Q1|B
.print DEVI L_MERGE|Q1|RB
.print V _JTL1|B|MID
.print V A
.print V _MERGE|A1|MID_SERIES
.print V _MERGE|B12|MID_SHUNT
.print V _MERGE|Q1
.print V _JTL5|2|MID_SHUNT
.print V B1
.print V _MERGE|B3
.print V _MERGE|A3
.print V _MERGE|A2
.print V _MERGE|Q2|MID_SHUNT
.print V _MERGE|Q2
.print V _MERGE|A1|MID_SHUNT
.print V _JTL5|4
.print V _MERGE|Q1|MID_SERIES
.print V _MERGE|A2|MID_SHUNT
.print V B
.print V _JTL3|4
.print V A_AND_B
.print V _MERGE|I_B1|MID
.print V _JTL1|6
.print V _JTL5|1
.print V _JTL3|2|MID_SERIES
.print V _MERGE|A12|MID_SHUNT
.print V _MERGE|B1
.print V _JTL3|6
.print V _MERGE|A1
.print V _JTL3|B|MID
.print V _JTL2|B|MID
.print V _MERGE|I_Q2|MID
.print V _MERGE|Q3
.print V _JTL1|1|MID_SHUNT
.print V _JTL2|2|MID_SERIES
.print V _JTL3|1|MID_SHUNT
.print V _JTL1|4
.print V _JTL5|B|MID
.print V _MERGE|B1|MID_SHUNT
.print V _JTL5|1|MID_SERIES
.print V _JTL5|2|MID_SERIES
.print V _JTL3|1
.print V _JTL2|2|MID_SHUNT
.print V _MERGE|B2
.print V _MERGE|I_Q1|MID
.print V _MERGE|B1|MID_SERIES
.print V _JTL2|6
.print V 2
.print V _MERGE|B2|MID_SHUNT
.print V _MERGE|I_A1|MID
.print V _JTL2|1|MID_SERIES
.print V _MERGE|Q1|MID_SHUNT
.print V _JTL5|1|MID_SHUNT
.print V _MERGE|I_Q3|MID
.print V _MERGE|Q2|MID_SERIES
.print V _JTL2|4
.print V _JTL3|1|MID_SERIES
.print V 3
.print V 1
.print V _JTL2|1|MID_SHUNT
.print V _MERGE|A2|MID_SERIES
.print V _JTL1|2|MID_SERIES
.print V _JTL3|2|MID_SHUNT
.print V _JTL1|1
.print V _JTL2|1
.print V _JTL5|6
.print V _JTL1|1|MID_SERIES
.print V _MERGE|B2|MID_SERIES
.print V _JTL1|2|MID_SHUNT
.print DEVP B_JTL1|1|1
.print DEVP B_JTL1|2|1
.print DEVP B_JTL2|1|1
.print DEVP B_JTL2|2|1
.print DEVP B_JTL3|1|1
.print DEVP B_JTL3|2|1
.print DEVP B_JTL5|1|1
.print DEVP B_JTL5|2|1
.print DEVP B_MERGE|A1|1
.print DEVP B_MERGE|A2|1
.print DEVP B_MERGE|A12|1
.print DEVP B_MERGE|B1|1
.print DEVP B_MERGE|B2|1
.print DEVP B_MERGE|B12|1
.print DEVP B_MERGE|Q2|1
.print DEVP B_MERGE|Q1|1
