*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM GLOBAL_SCALE=1.0
.PARAM TCLOCK=1.2e-10
.PARAM OS=6e-12
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 2000E-12
R_S0 S0 0  1
R_S1 S1 0  1
R_S2 S2 0  1
R_S3 S3 0  1
R_S4 S4 0  1
I_VEC|A0 0 A0  PWL(0 0 3.06e-11 0 3.36e-11 0.0007 3.66e-11 0 2.706e-10 0 2.736e-10 0.0007 2.766e-10 0 3.906e-10 0 3.936e-10 0.0007 3.966e-10 0 5.106e-10 0 5.136e-10 0.0007 5.166e-10 0 6.306e-10 0 6.336e-10 0.0007 6.366e-10 0 8.706e-10 0 8.736e-10 0.0007 8.766e-10 0 9.906e-10 0 9.936e-10 0.0007 9.966e-10 0 1.2306e-09 0 1.2336e-09 0.0007 1.2366e-09 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|A1 0 A1  PWL(0 0 3.906e-10 0 3.936e-10 0.0007 3.966e-10 0 5.106e-10 0 5.136e-10 0.0007 5.166e-10 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|A2 0 A2  PWL(0 0 1.506e-10 0 1.536e-10 0.0007 1.566e-10 0 5.106e-10 0 5.136e-10 0.0007 5.166e-10 0 7.506e-10 0 7.536e-10 0.0007 7.566e-10 0 9.906e-10 0 9.936e-10 0.0007 9.966e-10 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|A3 0 A3  PWL(0 0 7.506e-10 0 7.536e-10 0.0007 7.566e-10 0 9.906e-10 0 9.936e-10 0.0007 9.966e-10 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|B0 0 B0  PWL(0 0 3.06e-11 0 3.36e-11 0.0007 3.66e-11 0 2.706e-10 0 2.736e-10 0.0007 2.766e-10 0 6.306e-10 0 6.336e-10 0.0007 6.366e-10 0 8.706e-10 0 8.736e-10 0.0007 8.766e-10 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|B1 0 B1  PWL(0 0 3.06e-11 0 3.36e-11 0.0007 3.66e-11 0 2.706e-10 0 2.736e-10 0.0007 2.766e-10 0 3.906e-10 0 3.936e-10 0.0007 3.966e-10 0 5.106e-10 0 5.136e-10 0.0007 5.166e-10 0 1.1106e-09 0 1.1136e-09 0.0007 1.1166e-09 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|B2 0 B2  PWL(0 0 3.06e-11 0 3.36e-11 0.0007 3.66e-11 0 1.506e-10 0 1.536e-10 0.0007 1.566e-10 0 2.706e-10 0 2.736e-10 0.0007 2.766e-10 0 5.106e-10 0 5.136e-10 0.0007 5.166e-10 0 6.306e-10 0 6.336e-10 0.0007 6.366e-10 0 8.706e-10 0 8.736e-10 0.0007 8.766e-10 0 9.906e-10 0 9.936e-10 0.0007 9.966e-10 0 1.1106e-09 0 1.1136e-09 0.0007 1.1166e-09 0 1.2306e-09 0 1.2336e-09 0.0007 1.2366e-09 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
I_VEC|B3 0 B3  PWL(0 0 3.06e-11 0 3.36e-11 0.0007 3.66e-11 0 1.506e-10 0 1.536e-10 0.0007 1.566e-10 0 3.906e-10 0 3.936e-10 0.0007 3.966e-10 0 8.706e-10 0 8.736e-10 0.0007 8.766e-10 0 1.2306e-09 0 1.2336e-09 0.0007 1.2366e-09 0 1.3506e-09 0 1.3536e-09 0.0007 1.3566e-09 0)
IT00|T 0 T00  PWL(0 0 2.1e-11 0 2.4e-11 0.0021 2.7e-11 0 1.41e-10 0 1.44e-10 0.0021 1.47e-10 0 2.61e-10 0 2.64e-10 0.0021 2.67e-10 0 3.81e-10 0 3.84e-10 0.0021 3.87e-10 0 5.01e-10 0 5.04e-10 0.0021 5.07e-10 0 6.21e-10 0 6.24e-10 0.0021 6.27e-10 0 7.41e-10 0 7.44e-10 0.0021 7.47e-10 0 8.61e-10 0 8.64e-10 0.0021 8.67e-10 0 9.81e-10 0 9.84e-10 0.0021 9.87e-10 0 1.101e-09 0 1.104e-09 0.0021 1.107e-09 0 1.221e-09 0 1.224e-09 0.0021 1.227e-09 0 1.341e-09 0 1.344e-09 0.0021 1.347e-09 0 1.461e-09 0 1.464e-09 0.0021 1.467e-09 0 1.581e-09 0 1.584e-09 0.0021 1.587e-09 0 1.701e-09 0 1.704e-09 0.0021 1.707e-09 0 1.821e-09 0 1.824e-09 0.0021 1.827e-09 0 1.941e-09 0 1.944e-09 0.0021 1.947e-09 0 2.061e-09 0 2.064e-09 0.0021 2.067e-09 0 2.181e-09 0 2.184e-09 0.0021 2.187e-09 0 2.301e-09 0 2.304e-09 0.0021 2.307e-09 0 2.421e-09 0 2.424e-09 0.0021 2.427e-09 0 2.541e-09 0 2.544e-09 0.0021 2.547e-09 0 2.661e-09 0 2.664e-09 0.0021 2.667e-09 0 2.781e-09 0 2.784e-09 0.0021 2.787e-09 0 2.901e-09 0 2.904e-09 0.0021 2.907e-09 0 3.021e-09 0 3.024e-09 0.0021 3.027e-09 0 3.141e-09 0 3.144e-09 0.0021 3.147e-09 0 3.261e-09 0 3.264e-09 0.0021 3.267e-09 0 3.381e-09 0 3.384e-09 0.0021 3.387e-09 0 3.501e-09 0 3.504e-09 0.0021 3.507e-09 0 3.621e-09 0 3.624e-09 0.0021 3.627e-09 0 3.741e-09 0 3.744e-09 0.0021 3.747e-09 0 3.861e-09 0 3.864e-09 0.0021 3.867e-09 0 3.981e-09 0 3.984e-09 0.0021 3.987e-09 0 4.101e-09 0 4.104e-09 0.0021 4.107e-09 0 4.221e-09 0 4.224e-09 0.0021 4.227e-09 0 4.341e-09 0 4.344e-09 0.0021 4.347e-09 0 4.461e-09 0 4.464e-09 0.0021 4.467e-09 0 4.581e-09 0 4.584e-09 0.0021 4.587e-09 0 4.701e-09 0 4.704e-09 0.0021 4.707e-09 0 4.821e-09 0 4.824e-09 0.0021 4.827e-09 0 4.941e-09 0 4.944e-09 0.0021 4.947e-09 0 5.061e-09 0 5.064e-09 0.0021 5.067e-09 0 5.181e-09 0 5.184e-09 0.0021 5.187e-09 0 5.301e-09 0 5.304e-09 0.0021 5.307e-09 0 5.421e-09 0 5.424e-09 0.0021 5.427e-09 0 5.541e-09 0 5.544e-09 0.0021 5.547e-09 0 5.661e-09 0 5.664e-09 0.0021 5.667e-09 0 5.781e-09 0 5.784e-09 0.0021 5.787e-09 0 5.901e-09 0 5.904e-09 0.0021 5.907e-09 0 6.021e-09 0 6.024e-09 0.0021 6.027e-09 0 6.141e-09 0 6.144e-09 0.0021 6.147e-09 0 6.261e-09 0 6.264e-09 0.0021 6.267e-09 0 6.381e-09 0 6.384e-09 0.0021 6.387e-09 0 6.501e-09 0 6.504e-09 0.0021 6.507e-09 0 6.621e-09 0 6.624e-09 0.0021 6.627e-09 0 6.741e-09 0 6.744e-09 0.0021 6.747e-09 0 6.861e-09 0 6.864e-09 0.0021 6.867e-09 0 6.981e-09 0 6.984e-09 0.0021 6.987e-09 0 7.101e-09 0 7.104e-09 0.0021 7.107e-09 0 7.221e-09 0 7.224e-09 0.0021 7.227e-09 0 7.341e-09 0 7.344e-09 0.0021 7.347e-09 0 7.461e-09 0 7.464e-09 0.0021 7.467e-09 0 7.581e-09 0 7.584e-09 0.0021 7.587e-09 0 7.701e-09 0 7.704e-09 0.0021 7.707e-09 0 7.821e-09 0 7.824e-09 0.0021 7.827e-09 0 7.941e-09 0 7.944e-09 0.0021 7.947e-09 0 8.061e-09 0 8.064e-09 0.0021 8.067e-09 0 8.181e-09 0 8.184e-09 0.0021 8.187e-09 0 8.301e-09 0 8.304e-09 0.0021 8.307e-09 0 8.421e-09 0 8.424e-09 0.0021 8.427e-09 0 8.541e-09 0 8.544e-09 0.0021 8.547e-09 0 8.661e-09 0 8.664e-09 0.0021 8.667e-09 0 8.781e-09 0 8.784e-09 0.0021 8.787e-09 0 8.901e-09 0 8.904e-09 0.0021 8.907e-09 0 9.021e-09 0 9.024e-09 0.0021 9.027e-09 0 9.141e-09 0 9.144e-09 0.0021 9.147e-09 0 9.261e-09 0 9.264e-09 0.0021 9.267e-09 0 9.381e-09 0 9.384e-09 0.0021 9.387e-09 0 9.501e-09 0 9.504e-09 0.0021 9.507e-09 0 9.621e-09 0 9.624e-09 0.0021 9.627e-09 0 9.741e-09 0 9.744e-09 0.0021 9.747e-09 0 9.861e-09 0 9.864e-09 0.0021 9.867e-09 0 9.981e-09 0 9.984e-09 0.0021 9.987e-09 0 1.0101e-08 0 1.0104e-08 0.0021 1.0107e-08 0 1.0221e-08 0 1.0224e-08 0.0021 1.0227e-08 0 1.0341e-08 0 1.0344e-08 0.0021 1.0347e-08 0 1.0461e-08 0 1.0464e-08 0.0021 1.0467e-08 0 1.0581e-08 0 1.0584e-08 0.0021 1.0587e-08 0 1.0701e-08 0 1.0704e-08 0.0021 1.0707e-08 0 1.0821e-08 0 1.0824e-08 0.0021 1.0827e-08 0 1.0941e-08 0 1.0944e-08 0.0021 1.0947e-08 0 1.1061e-08 0 1.1064e-08 0.0021 1.1067e-08 0 1.1181e-08 0 1.1184e-08 0.0021 1.1187e-08 0 1.1301e-08 0 1.1304e-08 0.0021 1.1307e-08 0 1.1421e-08 0 1.1424e-08 0.0021 1.1427e-08 0 1.1541e-08 0 1.1544e-08 0.0021 1.1547e-08 0 1.1661e-08 0 1.1664e-08 0.0021 1.1667e-08 0 1.1781e-08 0 1.1784e-08 0.0021 1.1787e-08 0 1.1901e-08 0 1.1904e-08 0.0021 1.1907e-08 0 1.2021e-08 0 1.2024e-08 0.0021 1.2027e-08 0 1.2141e-08 0 1.2144e-08 0.0021 1.2147e-08 0 1.2261e-08 0 1.2264e-08 0.0021 1.2267e-08 0 1.2381e-08 0 1.2384e-08 0.0021 1.2387e-08 0 1.2501e-08 0 1.2504e-08 0.0021 1.2507e-08 0 1.2621e-08 0 1.2624e-08 0.0021 1.2627e-08 0 1.2741e-08 0 1.2744e-08 0.0021 1.2747e-08 0 1.2861e-08 0 1.2864e-08 0.0021 1.2867e-08 0 1.2981e-08 0 1.2984e-08 0.0021 1.2987e-08 0 1.3101e-08 0 1.3104e-08 0.0021 1.3107e-08 0 1.3221e-08 0 1.3224e-08 0.0021 1.3227e-08 0 1.3341e-08 0 1.3344e-08 0.0021 1.3347e-08 0 1.3461e-08 0 1.3464e-08 0.0021 1.3467e-08 0 1.3581e-08 0 1.3584e-08 0.0021 1.3587e-08 0 1.3701e-08 0 1.3704e-08 0.0021 1.3707e-08 0 1.3821e-08 0 1.3824e-08 0.0021 1.3827e-08 0 1.3941e-08 0 1.3944e-08 0.0021 1.3947e-08 0 1.4061e-08 0 1.4064e-08 0.0021 1.4067e-08 0 1.4181e-08 0 1.4184e-08 0.0021 1.4187e-08 0 1.4301e-08 0 1.4304e-08 0.0021 1.4307e-08 0 1.4421e-08 0 1.4424e-08 0.0021 1.4427e-08 0 1.4541e-08 0 1.4544e-08 0.0021 1.4547e-08 0 1.4661e-08 0 1.4664e-08 0.0021 1.4667e-08 0 1.4781e-08 0 1.4784e-08 0.0021 1.4787e-08 0 1.4901e-08 0 1.4904e-08 0.0021 1.4907e-08 0 1.5021e-08 0 1.5024e-08 0.0021 1.5027e-08 0 1.5141e-08 0 1.5144e-08 0.0021 1.5147e-08 0 1.5261e-08 0 1.5264e-08 0.0021 1.5267e-08 0 1.5381e-08 0 1.5384e-08 0.0021 1.5387e-08 0 1.5501e-08 0 1.5504e-08 0.0021 1.5507e-08 0 1.5621e-08 0 1.5624e-08 0.0021 1.5627e-08 0 1.5741e-08 0 1.5744e-08 0.0021 1.5747e-08 0 1.5861e-08 0 1.5864e-08 0.0021 1.5867e-08 0 1.5981e-08 0 1.5984e-08 0.0021 1.5987e-08 0 1.6101e-08 0 1.6104e-08 0.0021 1.6107e-08 0 1.6221e-08 0 1.6224e-08 0.0021 1.6227e-08 0 1.6341e-08 0 1.6344e-08 0.0021 1.6347e-08 0 1.6461e-08 0 1.6464e-08 0.0021 1.6467e-08 0 1.6581e-08 0 1.6584e-08 0.0021 1.6587e-08 0 1.6701e-08 0 1.6704e-08 0.0021 1.6707e-08 0 1.6821e-08 0 1.6824e-08 0.0021 1.6827e-08 0 1.6941e-08 0 1.6944e-08 0.0021 1.6947e-08 0 1.7061e-08 0 1.7064e-08 0.0021 1.7067e-08 0 1.7181e-08 0 1.7184e-08 0.0021 1.7187e-08 0 1.7301e-08 0 1.7304e-08 0.0021 1.7307e-08 0 1.7421e-08 0 1.7424e-08 0.0021 1.7427e-08 0 1.7541e-08 0 1.7544e-08 0.0021 1.7547e-08 0 1.7661e-08 0 1.7664e-08 0.0021 1.7667e-08 0 1.7781e-08 0 1.7784e-08 0.0021 1.7787e-08 0 1.7901e-08 0 1.7904e-08 0.0021 1.7907e-08 0 1.8021e-08 0 1.8024e-08 0.0021 1.8027e-08 0 1.8141e-08 0 1.8144e-08 0.0021 1.8147e-08 0 1.8261e-08 0 1.8264e-08 0.0021 1.8267e-08 0 1.8381e-08 0 1.8384e-08 0.0021 1.8387e-08 0 1.8501e-08 0 1.8504e-08 0.0021 1.8507e-08 0 1.8621e-08 0 1.8624e-08 0.0021 1.8627e-08 0 1.8741e-08 0 1.8744e-08 0.0021 1.8747e-08 0 1.8861e-08 0 1.8864e-08 0.0021 1.8867e-08 0 1.8981e-08 0 1.8984e-08 0.0021 1.8987e-08 0 1.9101e-08 0 1.9104e-08 0.0021 1.9107e-08 0 1.9221e-08 0 1.9224e-08 0.0021 1.9227e-08 0 1.9341e-08 0 1.9344e-08 0.0021 1.9347e-08 0 1.9461e-08 0 1.9464e-08 0.0021 1.9467e-08 0 1.9581e-08 0 1.9584e-08 0.0021 1.9587e-08 0 1.9701e-08 0 1.9704e-08 0.0021 1.9707e-08 0 1.9821e-08 0 1.9824e-08 0.0021 1.9827e-08 0 1.9941e-08 0 1.9944e-08 0.0021 1.9947e-08 0 2.0061e-08 0 2.0064e-08 0.0021 2.0067e-08 0 2.0181e-08 0 2.0184e-08 0.0021 2.0187e-08 0 2.0301e-08 0 2.0304e-08 0.0021 2.0307e-08 0 2.0421e-08 0 2.0424e-08 0.0021 2.0427e-08 0 2.0541e-08 0 2.0544e-08 0.0021 2.0547e-08 0 2.0661e-08 0 2.0664e-08 0.0021 2.0667e-08 0 2.0781e-08 0 2.0784e-08 0.0021 2.0787e-08 0 2.0901e-08 0 2.0904e-08 0.0021 2.0907e-08 0 2.1021e-08 0 2.1024e-08 0.0021 2.1027e-08 0 2.1141e-08 0 2.1144e-08 0.0021 2.1147e-08 0 2.1261e-08 0 2.1264e-08 0.0021 2.1267e-08 0 2.1381e-08 0 2.1384e-08 0.0021 2.1387e-08 0 2.1501e-08 0 2.1504e-08 0.0021 2.1507e-08 0 2.1621e-08 0 2.1624e-08 0.0021 2.1627e-08 0 2.1741e-08 0 2.1744e-08 0.0021 2.1747e-08 0 2.1861e-08 0 2.1864e-08 0.0021 2.1867e-08 0 2.1981e-08 0 2.1984e-08 0.0021 2.1987e-08 0 2.2101e-08 0 2.2104e-08 0.0021 2.2107e-08 0 2.2221e-08 0 2.2224e-08 0.0021 2.2227e-08 0 2.2341e-08 0 2.2344e-08 0.0021 2.2347e-08 0 2.2461e-08 0 2.2464e-08 0.0021 2.2467e-08 0 2.2581e-08 0 2.2584e-08 0.0021 2.2587e-08 0 2.2701e-08 0 2.2704e-08 0.0021 2.2707e-08 0 2.2821e-08 0 2.2824e-08 0.0021 2.2827e-08 0 2.2941e-08 0 2.2944e-08 0.0021 2.2947e-08 0 2.3061e-08 0 2.3064e-08 0.0021 2.3067e-08 0 2.3181e-08 0 2.3184e-08 0.0021 2.3187e-08 0 2.3301e-08 0 2.3304e-08 0.0021 2.3307e-08 0 2.3421e-08 0 2.3424e-08 0.0021 2.3427e-08 0 2.3541e-08 0 2.3544e-08 0.0021 2.3547e-08 0 2.3661e-08 0 2.3664e-08 0.0021 2.3667e-08 0 2.3781e-08 0 2.3784e-08 0.0021 2.3787e-08 0 2.3901e-08 0 2.3904e-08 0.0021 2.3907e-08 0 2.4021e-08 0 2.4024e-08 0.0021 2.4027e-08 0 2.4141e-08 0 2.4144e-08 0.0021 2.4147e-08 0 2.4261e-08 0 2.4264e-08 0.0021 2.4267e-08 0 2.4381e-08 0 2.4384e-08 0.0021 2.4387e-08 0 2.4501e-08 0 2.4504e-08 0.0021 2.4507e-08 0 2.4621e-08 0 2.4624e-08 0.0021 2.4627e-08 0 2.4741e-08 0 2.4744e-08 0.0021 2.4747e-08 0 2.4861e-08 0 2.4864e-08 0.0021 2.4867e-08 0 2.4981e-08 0 2.4984e-08 0.0021 2.4987e-08 0 2.5101e-08 0 2.5104e-08 0.0021 2.5107e-08 0 2.5221e-08 0 2.5224e-08 0.0021 2.5227e-08 0 2.5341e-08 0 2.5344e-08 0.0021 2.5347e-08 0 2.5461e-08 0 2.5464e-08 0.0021 2.5467e-08 0 2.5581e-08 0 2.5584e-08 0.0021 2.5587e-08 0 2.5701e-08 0 2.5704e-08 0.0021 2.5707e-08 0 2.5821e-08 0 2.5824e-08 0.0021 2.5827e-08 0 2.5941e-08 0 2.5944e-08 0.0021 2.5947e-08 0 2.6061e-08 0 2.6064e-08 0.0021 2.6067e-08 0 2.6181e-08 0 2.6184e-08 0.0021 2.6187e-08 0 2.6301e-08 0 2.6304e-08 0.0021 2.6307e-08 0 2.6421e-08 0 2.6424e-08 0.0021 2.6427e-08 0 2.6541e-08 0 2.6544e-08 0.0021 2.6547e-08 0 2.6661e-08 0 2.6664e-08 0.0021 2.6667e-08 0 2.6781e-08 0 2.6784e-08 0.0021 2.6787e-08 0 2.6901e-08 0 2.6904e-08 0.0021 2.6907e-08 0 2.7021e-08 0 2.7024e-08 0.0021 2.7027e-08 0 2.7141e-08 0 2.7144e-08 0.0021 2.7147e-08 0 2.7261e-08 0 2.7264e-08 0.0021 2.7267e-08 0 2.7381e-08 0 2.7384e-08 0.0021 2.7387e-08 0 2.7501e-08 0 2.7504e-08 0.0021 2.7507e-08 0 2.7621e-08 0 2.7624e-08 0.0021 2.7627e-08 0 2.7741e-08 0 2.7744e-08 0.0021 2.7747e-08 0 2.7861e-08 0 2.7864e-08 0.0021 2.7867e-08 0 2.7981e-08 0 2.7984e-08 0.0021 2.7987e-08 0 2.8101e-08 0 2.8104e-08 0.0021 2.8107e-08 0 2.8221e-08 0 2.8224e-08 0.0021 2.8227e-08 0 2.8341e-08 0 2.8344e-08 0.0021 2.8347e-08 0 2.8461e-08 0 2.8464e-08 0.0021 2.8467e-08 0 2.8581e-08 0 2.8584e-08 0.0021 2.8587e-08 0 2.8701e-08 0 2.8704e-08 0.0021 2.8707e-08 0 2.8821e-08 0 2.8824e-08 0.0021 2.8827e-08 0 2.8941e-08 0 2.8944e-08 0.0021 2.8947e-08 0 2.9061e-08 0 2.9064e-08 0.0021 2.9067e-08 0 2.9181e-08 0 2.9184e-08 0.0021 2.9187e-08 0 2.9301e-08 0 2.9304e-08 0.0021 2.9307e-08 0 2.9421e-08 0 2.9424e-08 0.0021 2.9427e-08 0 2.9541e-08 0 2.9544e-08 0.0021 2.9547e-08 0 2.9661e-08 0 2.9664e-08 0.0021 2.9667e-08 0 2.9781e-08 0 2.9784e-08 0.0021 2.9787e-08 0 2.9901e-08 0 2.9904e-08 0.0021 2.9907e-08 0 3.0021e-08 0 3.0024e-08 0.0021 3.0027e-08 0 3.0141e-08 0 3.0144e-08 0.0021 3.0147e-08 0 3.0261e-08 0 3.0264e-08 0.0021 3.0267e-08 0 3.0381e-08 0 3.0384e-08 0.0021 3.0387e-08 0 3.0501e-08 0 3.0504e-08 0.0021 3.0507e-08 0 3.0621e-08 0 3.0624e-08 0.0021 3.0627e-08 0 3.0741e-08 0 3.0744e-08 0.0021 3.0747e-08 0 3.0861e-08 0 3.0864e-08 0.0021 3.0867e-08 0 3.0981e-08 0 3.0984e-08 0.0021 3.0987e-08 0 3.1101e-08 0 3.1104e-08 0.0021 3.1107e-08 0 3.1221e-08 0 3.1224e-08 0.0021 3.1227e-08 0 3.1341e-08 0 3.1344e-08 0.0021 3.1347e-08 0 3.1461e-08 0 3.1464e-08 0.0021 3.1467e-08 0 3.1581e-08 0 3.1584e-08 0.0021 3.1587e-08 0 3.1701e-08 0 3.1704e-08 0.0021 3.1707e-08 0 3.1821e-08 0 3.1824e-08 0.0021 3.1827e-08 0 3.1941e-08 0 3.1944e-08 0.0021 3.1947e-08 0 3.2061e-08 0 3.2064e-08 0.0021 3.2067e-08 0 3.2181e-08 0 3.2184e-08 0.0021 3.2187e-08 0 3.2301e-08 0 3.2304e-08 0.0021 3.2307e-08 0 3.2421e-08 0 3.2424e-08 0.0021 3.2427e-08 0 3.2541e-08 0 3.2544e-08 0.0021 3.2547e-08 0 3.2661e-08 0 3.2664e-08 0.0021 3.2667e-08 0 3.2781e-08 0 3.2784e-08 0.0021 3.2787e-08 0 3.2901e-08 0 3.2904e-08 0.0021 3.2907e-08 0 3.3021e-08 0 3.3024e-08 0.0021 3.3027e-08 0 3.3141e-08 0 3.3144e-08 0.0021 3.3147e-08 0 3.3261e-08 0 3.3264e-08 0.0021 3.3267e-08 0 3.3381e-08 0 3.3384e-08 0.0021 3.3387e-08 0 3.3501e-08 0 3.3504e-08 0.0021 3.3507e-08 0 3.3621e-08 0 3.3624e-08 0.0021 3.3627e-08 0 3.3741e-08 0 3.3744e-08 0.0021 3.3747e-08 0 3.3861e-08 0 3.3864e-08 0.0021 3.3867e-08 0 3.3981e-08 0 3.3984e-08 0.0021 3.3987e-08 0 3.4101e-08 0 3.4104e-08 0.0021 3.4107e-08 0 3.4221e-08 0 3.4224e-08 0.0021 3.4227e-08 0 3.4341e-08 0 3.4344e-08 0.0021 3.4347e-08 0 3.4461e-08 0 3.4464e-08 0.0021 3.4467e-08 0 3.4581e-08 0 3.4584e-08 0.0021 3.4587e-08 0 3.4701e-08 0 3.4704e-08 0.0021 3.4707e-08 0 3.4821e-08 0 3.4824e-08 0.0021 3.4827e-08 0 3.4941e-08 0 3.4944e-08 0.0021 3.4947e-08 0 3.5061e-08 0 3.5064e-08 0.0021 3.5067e-08 0 3.5181e-08 0 3.5184e-08 0.0021 3.5187e-08 0 3.5301e-08 0 3.5304e-08 0.0021 3.5307e-08 0 3.5421e-08 0 3.5424e-08 0.0021 3.5427e-08 0 3.5541e-08 0 3.5544e-08 0.0021 3.5547e-08 0 3.5661e-08 0 3.5664e-08 0.0021 3.5667e-08 0 3.5781e-08 0 3.5784e-08 0.0021 3.5787e-08 0 3.5901e-08 0 3.5904e-08 0.0021 3.5907e-08 0 3.6021e-08 0 3.6024e-08 0.0021 3.6027e-08 0 3.6141e-08 0 3.6144e-08 0.0021 3.6147e-08 0 3.6261e-08 0 3.6264e-08 0.0021 3.6267e-08 0 3.6381e-08 0 3.6384e-08 0.0021 3.6387e-08 0 3.6501e-08 0 3.6504e-08 0.0021 3.6507e-08 0 3.6621e-08 0 3.6624e-08 0.0021 3.6627e-08 0 3.6741e-08 0 3.6744e-08 0.0021 3.6747e-08 0 3.6861e-08 0 3.6864e-08 0.0021 3.6867e-08 0 3.6981e-08 0 3.6984e-08 0.0021 3.6987e-08 0 3.7101e-08 0 3.7104e-08 0.0021 3.7107e-08 0 3.7221e-08 0 3.7224e-08 0.0021 3.7227e-08 0 3.7341e-08 0 3.7344e-08 0.0021 3.7347e-08 0 3.7461e-08 0 3.7464e-08 0.0021 3.7467e-08 0 3.7581e-08 0 3.7584e-08 0.0021 3.7587e-08 0 3.7701e-08 0 3.7704e-08 0.0021 3.7707e-08 0 3.7821e-08 0 3.7824e-08 0.0021 3.7827e-08 0 3.7941e-08 0 3.7944e-08 0.0021 3.7947e-08 0 3.8061e-08 0 3.8064e-08 0.0021 3.8067e-08 0 3.8181e-08 0 3.8184e-08 0.0021 3.8187e-08 0 3.8301e-08 0 3.8304e-08 0.0021 3.8307e-08 0 3.8421e-08 0 3.8424e-08 0.0021 3.8427e-08 0 3.8541e-08 0 3.8544e-08 0.0021 3.8547e-08 0 3.8661e-08 0 3.8664e-08 0.0021 3.8667e-08 0 3.8781e-08 0 3.8784e-08 0.0021 3.8787e-08 0 3.8901e-08 0 3.8904e-08 0.0021 3.8907e-08 0 3.9021e-08 0 3.9024e-08 0.0021 3.9027e-08 0 3.9141e-08 0 3.9144e-08 0.0021 3.9147e-08 0 3.9261e-08 0 3.9264e-08 0.0021 3.9267e-08 0 3.9381e-08 0 3.9384e-08 0.0021 3.9387e-08 0 3.9501e-08 0 3.9504e-08 0.0021 3.9507e-08 0 3.9621e-08 0 3.9624e-08 0.0021 3.9627e-08 0 3.9741e-08 0 3.9744e-08 0.0021 3.9747e-08 0 3.9861e-08 0 3.9864e-08 0.0021 3.9867e-08 0 3.9981e-08 0 3.9984e-08 0.0021 3.9987e-08 0 4.0101e-08 0 4.0104e-08 0.0021 4.0107e-08 0 4.0221e-08 0 4.0224e-08 0.0021 4.0227e-08 0 4.0341e-08 0 4.0344e-08 0.0021 4.0347e-08 0 4.0461e-08 0 4.0464e-08 0.0021 4.0467e-08 0 4.0581e-08 0 4.0584e-08 0.0021 4.0587e-08 0 4.0701e-08 0 4.0704e-08 0.0021 4.0707e-08 0 4.0821e-08 0 4.0824e-08 0.0021 4.0827e-08 0 4.0941e-08 0 4.0944e-08 0.0021 4.0947e-08 0 4.1061e-08 0 4.1064e-08 0.0021 4.1067e-08 0 4.1181e-08 0 4.1184e-08 0.0021 4.1187e-08 0 4.1301e-08 0 4.1304e-08 0.0021 4.1307e-08 0 4.1421e-08 0 4.1424e-08 0.0021 4.1427e-08 0 4.1541e-08 0 4.1544e-08 0.0021 4.1547e-08 0 4.1661e-08 0 4.1664e-08 0.0021 4.1667e-08 0 4.1781e-08 0 4.1784e-08 0.0021 4.1787e-08 0 4.1901e-08 0 4.1904e-08 0.0021 4.1907e-08 0 4.2021e-08 0 4.2024e-08 0.0021 4.2027e-08 0 4.2141e-08 0 4.2144e-08 0.0021 4.2147e-08 0 4.2261e-08 0 4.2264e-08 0.0021 4.2267e-08 0 4.2381e-08 0 4.2384e-08 0.0021 4.2387e-08 0 4.2501e-08 0 4.2504e-08 0.0021 4.2507e-08 0 4.2621e-08 0 4.2624e-08 0.0021 4.2627e-08 0 4.2741e-08 0 4.2744e-08 0.0021 4.2747e-08 0 4.2861e-08 0 4.2864e-08 0.0021 4.2867e-08 0 4.2981e-08 0 4.2984e-08 0.0021 4.2987e-08 0 4.3101e-08 0 4.3104e-08 0.0021 4.3107e-08 0 4.3221e-08 0 4.3224e-08 0.0021 4.3227e-08 0 4.3341e-08 0 4.3344e-08 0.0021 4.3347e-08 0 4.3461e-08 0 4.3464e-08 0.0021 4.3467e-08 0 4.3581e-08 0 4.3584e-08 0.0021 4.3587e-08 0 4.3701e-08 0 4.3704e-08 0.0021 4.3707e-08 0 4.3821e-08 0 4.3824e-08 0.0021 4.3827e-08 0 4.3941e-08 0 4.3944e-08 0.0021 4.3947e-08 0 4.4061e-08 0 4.4064e-08 0.0021 4.4067e-08 0 4.4181e-08 0 4.4184e-08 0.0021 4.4187e-08 0 4.4301e-08 0 4.4304e-08 0.0021 4.4307e-08 0 4.4421e-08 0 4.4424e-08 0.0021 4.4427e-08 0 4.4541e-08 0 4.4544e-08 0.0021 4.4547e-08 0 4.4661e-08 0 4.4664e-08 0.0021 4.4667e-08 0 4.4781e-08 0 4.4784e-08 0.0021 4.4787e-08 0 4.4901e-08 0 4.4904e-08 0.0021 4.4907e-08 0 4.5021e-08 0 4.5024e-08 0.0021 4.5027e-08 0 4.5141e-08 0 4.5144e-08 0.0021 4.5147e-08 0 4.5261e-08 0 4.5264e-08 0.0021 4.5267e-08 0 4.5381e-08 0 4.5384e-08 0.0021 4.5387e-08 0 4.5501e-08 0 4.5504e-08 0.0021 4.5507e-08 0 4.5621e-08 0 4.5624e-08 0.0021 4.5627e-08 0 4.5741e-08 0 4.5744e-08 0.0021 4.5747e-08 0 4.5861e-08 0 4.5864e-08 0.0021 4.5867e-08 0 4.5981e-08 0 4.5984e-08 0.0021 4.5987e-08 0 4.6101e-08 0 4.6104e-08 0.0021 4.6107e-08 0 4.6221e-08 0 4.6224e-08 0.0021 4.6227e-08 0 4.6341e-08 0 4.6344e-08 0.0021 4.6347e-08 0 4.6461e-08 0 4.6464e-08 0.0021 4.6467e-08 0 4.6581e-08 0 4.6584e-08 0.0021 4.6587e-08 0 4.6701e-08 0 4.6704e-08 0.0021 4.6707e-08 0 4.6821e-08 0 4.6824e-08 0.0021 4.6827e-08 0 4.6941e-08 0 4.6944e-08 0.0021 4.6947e-08 0 4.7061e-08 0 4.7064e-08 0.0021 4.7067e-08 0 4.7181e-08 0 4.7184e-08 0.0021 4.7187e-08 0 4.7301e-08 0 4.7304e-08 0.0021 4.7307e-08 0 4.7421e-08 0 4.7424e-08 0.0021 4.7427e-08 0 4.7541e-08 0 4.7544e-08 0.0021 4.7547e-08 0 4.7661e-08 0 4.7664e-08 0.0021 4.7667e-08 0 4.7781e-08 0 4.7784e-08 0.0021 4.7787e-08 0)
IT01|T 0 T01  PWL(0 0 2.1e-11 0 2.4e-11 0.0021 2.7e-11 0 1.41e-10 0 1.44e-10 0.0021 1.47e-10 0 2.61e-10 0 2.64e-10 0.0021 2.67e-10 0 3.81e-10 0 3.84e-10 0.0021 3.87e-10 0 5.01e-10 0 5.04e-10 0.0021 5.07e-10 0 6.21e-10 0 6.24e-10 0.0021 6.27e-10 0 7.41e-10 0 7.44e-10 0.0021 7.47e-10 0 8.61e-10 0 8.64e-10 0.0021 8.67e-10 0 9.81e-10 0 9.84e-10 0.0021 9.87e-10 0 1.101e-09 0 1.104e-09 0.0021 1.107e-09 0 1.221e-09 0 1.224e-09 0.0021 1.227e-09 0 1.341e-09 0 1.344e-09 0.0021 1.347e-09 0 1.461e-09 0 1.464e-09 0.0021 1.467e-09 0 1.581e-09 0 1.584e-09 0.0021 1.587e-09 0 1.701e-09 0 1.704e-09 0.0021 1.707e-09 0 1.821e-09 0 1.824e-09 0.0021 1.827e-09 0 1.941e-09 0 1.944e-09 0.0021 1.947e-09 0 2.061e-09 0 2.064e-09 0.0021 2.067e-09 0 2.181e-09 0 2.184e-09 0.0021 2.187e-09 0 2.301e-09 0 2.304e-09 0.0021 2.307e-09 0 2.421e-09 0 2.424e-09 0.0021 2.427e-09 0 2.541e-09 0 2.544e-09 0.0021 2.547e-09 0 2.661e-09 0 2.664e-09 0.0021 2.667e-09 0 2.781e-09 0 2.784e-09 0.0021 2.787e-09 0 2.901e-09 0 2.904e-09 0.0021 2.907e-09 0 3.021e-09 0 3.024e-09 0.0021 3.027e-09 0 3.141e-09 0 3.144e-09 0.0021 3.147e-09 0 3.261e-09 0 3.264e-09 0.0021 3.267e-09 0 3.381e-09 0 3.384e-09 0.0021 3.387e-09 0 3.501e-09 0 3.504e-09 0.0021 3.507e-09 0 3.621e-09 0 3.624e-09 0.0021 3.627e-09 0 3.741e-09 0 3.744e-09 0.0021 3.747e-09 0 3.861e-09 0 3.864e-09 0.0021 3.867e-09 0 3.981e-09 0 3.984e-09 0.0021 3.987e-09 0 4.101e-09 0 4.104e-09 0.0021 4.107e-09 0 4.221e-09 0 4.224e-09 0.0021 4.227e-09 0 4.341e-09 0 4.344e-09 0.0021 4.347e-09 0 4.461e-09 0 4.464e-09 0.0021 4.467e-09 0 4.581e-09 0 4.584e-09 0.0021 4.587e-09 0 4.701e-09 0 4.704e-09 0.0021 4.707e-09 0 4.821e-09 0 4.824e-09 0.0021 4.827e-09 0 4.941e-09 0 4.944e-09 0.0021 4.947e-09 0 5.061e-09 0 5.064e-09 0.0021 5.067e-09 0 5.181e-09 0 5.184e-09 0.0021 5.187e-09 0 5.301e-09 0 5.304e-09 0.0021 5.307e-09 0 5.421e-09 0 5.424e-09 0.0021 5.427e-09 0 5.541e-09 0 5.544e-09 0.0021 5.547e-09 0 5.661e-09 0 5.664e-09 0.0021 5.667e-09 0 5.781e-09 0 5.784e-09 0.0021 5.787e-09 0 5.901e-09 0 5.904e-09 0.0021 5.907e-09 0 6.021e-09 0 6.024e-09 0.0021 6.027e-09 0 6.141e-09 0 6.144e-09 0.0021 6.147e-09 0 6.261e-09 0 6.264e-09 0.0021 6.267e-09 0 6.381e-09 0 6.384e-09 0.0021 6.387e-09 0 6.501e-09 0 6.504e-09 0.0021 6.507e-09 0 6.621e-09 0 6.624e-09 0.0021 6.627e-09 0 6.741e-09 0 6.744e-09 0.0021 6.747e-09 0 6.861e-09 0 6.864e-09 0.0021 6.867e-09 0 6.981e-09 0 6.984e-09 0.0021 6.987e-09 0 7.101e-09 0 7.104e-09 0.0021 7.107e-09 0 7.221e-09 0 7.224e-09 0.0021 7.227e-09 0 7.341e-09 0 7.344e-09 0.0021 7.347e-09 0 7.461e-09 0 7.464e-09 0.0021 7.467e-09 0 7.581e-09 0 7.584e-09 0.0021 7.587e-09 0 7.701e-09 0 7.704e-09 0.0021 7.707e-09 0 7.821e-09 0 7.824e-09 0.0021 7.827e-09 0 7.941e-09 0 7.944e-09 0.0021 7.947e-09 0 8.061e-09 0 8.064e-09 0.0021 8.067e-09 0 8.181e-09 0 8.184e-09 0.0021 8.187e-09 0 8.301e-09 0 8.304e-09 0.0021 8.307e-09 0 8.421e-09 0 8.424e-09 0.0021 8.427e-09 0 8.541e-09 0 8.544e-09 0.0021 8.547e-09 0 8.661e-09 0 8.664e-09 0.0021 8.667e-09 0 8.781e-09 0 8.784e-09 0.0021 8.787e-09 0 8.901e-09 0 8.904e-09 0.0021 8.907e-09 0 9.021e-09 0 9.024e-09 0.0021 9.027e-09 0 9.141e-09 0 9.144e-09 0.0021 9.147e-09 0 9.261e-09 0 9.264e-09 0.0021 9.267e-09 0 9.381e-09 0 9.384e-09 0.0021 9.387e-09 0 9.501e-09 0 9.504e-09 0.0021 9.507e-09 0 9.621e-09 0 9.624e-09 0.0021 9.627e-09 0 9.741e-09 0 9.744e-09 0.0021 9.747e-09 0 9.861e-09 0 9.864e-09 0.0021 9.867e-09 0 9.981e-09 0 9.984e-09 0.0021 9.987e-09 0 1.0101e-08 0 1.0104e-08 0.0021 1.0107e-08 0 1.0221e-08 0 1.0224e-08 0.0021 1.0227e-08 0 1.0341e-08 0 1.0344e-08 0.0021 1.0347e-08 0 1.0461e-08 0 1.0464e-08 0.0021 1.0467e-08 0 1.0581e-08 0 1.0584e-08 0.0021 1.0587e-08 0 1.0701e-08 0 1.0704e-08 0.0021 1.0707e-08 0 1.0821e-08 0 1.0824e-08 0.0021 1.0827e-08 0 1.0941e-08 0 1.0944e-08 0.0021 1.0947e-08 0 1.1061e-08 0 1.1064e-08 0.0021 1.1067e-08 0 1.1181e-08 0 1.1184e-08 0.0021 1.1187e-08 0 1.1301e-08 0 1.1304e-08 0.0021 1.1307e-08 0 1.1421e-08 0 1.1424e-08 0.0021 1.1427e-08 0 1.1541e-08 0 1.1544e-08 0.0021 1.1547e-08 0 1.1661e-08 0 1.1664e-08 0.0021 1.1667e-08 0 1.1781e-08 0 1.1784e-08 0.0021 1.1787e-08 0 1.1901e-08 0 1.1904e-08 0.0021 1.1907e-08 0 1.2021e-08 0 1.2024e-08 0.0021 1.2027e-08 0 1.2141e-08 0 1.2144e-08 0.0021 1.2147e-08 0 1.2261e-08 0 1.2264e-08 0.0021 1.2267e-08 0 1.2381e-08 0 1.2384e-08 0.0021 1.2387e-08 0 1.2501e-08 0 1.2504e-08 0.0021 1.2507e-08 0 1.2621e-08 0 1.2624e-08 0.0021 1.2627e-08 0 1.2741e-08 0 1.2744e-08 0.0021 1.2747e-08 0 1.2861e-08 0 1.2864e-08 0.0021 1.2867e-08 0 1.2981e-08 0 1.2984e-08 0.0021 1.2987e-08 0 1.3101e-08 0 1.3104e-08 0.0021 1.3107e-08 0 1.3221e-08 0 1.3224e-08 0.0021 1.3227e-08 0 1.3341e-08 0 1.3344e-08 0.0021 1.3347e-08 0 1.3461e-08 0 1.3464e-08 0.0021 1.3467e-08 0 1.3581e-08 0 1.3584e-08 0.0021 1.3587e-08 0 1.3701e-08 0 1.3704e-08 0.0021 1.3707e-08 0 1.3821e-08 0 1.3824e-08 0.0021 1.3827e-08 0 1.3941e-08 0 1.3944e-08 0.0021 1.3947e-08 0 1.4061e-08 0 1.4064e-08 0.0021 1.4067e-08 0 1.4181e-08 0 1.4184e-08 0.0021 1.4187e-08 0 1.4301e-08 0 1.4304e-08 0.0021 1.4307e-08 0 1.4421e-08 0 1.4424e-08 0.0021 1.4427e-08 0 1.4541e-08 0 1.4544e-08 0.0021 1.4547e-08 0 1.4661e-08 0 1.4664e-08 0.0021 1.4667e-08 0 1.4781e-08 0 1.4784e-08 0.0021 1.4787e-08 0 1.4901e-08 0 1.4904e-08 0.0021 1.4907e-08 0 1.5021e-08 0 1.5024e-08 0.0021 1.5027e-08 0 1.5141e-08 0 1.5144e-08 0.0021 1.5147e-08 0 1.5261e-08 0 1.5264e-08 0.0021 1.5267e-08 0 1.5381e-08 0 1.5384e-08 0.0021 1.5387e-08 0 1.5501e-08 0 1.5504e-08 0.0021 1.5507e-08 0 1.5621e-08 0 1.5624e-08 0.0021 1.5627e-08 0 1.5741e-08 0 1.5744e-08 0.0021 1.5747e-08 0 1.5861e-08 0 1.5864e-08 0.0021 1.5867e-08 0 1.5981e-08 0 1.5984e-08 0.0021 1.5987e-08 0 1.6101e-08 0 1.6104e-08 0.0021 1.6107e-08 0 1.6221e-08 0 1.6224e-08 0.0021 1.6227e-08 0 1.6341e-08 0 1.6344e-08 0.0021 1.6347e-08 0 1.6461e-08 0 1.6464e-08 0.0021 1.6467e-08 0 1.6581e-08 0 1.6584e-08 0.0021 1.6587e-08 0 1.6701e-08 0 1.6704e-08 0.0021 1.6707e-08 0 1.6821e-08 0 1.6824e-08 0.0021 1.6827e-08 0 1.6941e-08 0 1.6944e-08 0.0021 1.6947e-08 0 1.7061e-08 0 1.7064e-08 0.0021 1.7067e-08 0 1.7181e-08 0 1.7184e-08 0.0021 1.7187e-08 0 1.7301e-08 0 1.7304e-08 0.0021 1.7307e-08 0 1.7421e-08 0 1.7424e-08 0.0021 1.7427e-08 0 1.7541e-08 0 1.7544e-08 0.0021 1.7547e-08 0 1.7661e-08 0 1.7664e-08 0.0021 1.7667e-08 0 1.7781e-08 0 1.7784e-08 0.0021 1.7787e-08 0 1.7901e-08 0 1.7904e-08 0.0021 1.7907e-08 0 1.8021e-08 0 1.8024e-08 0.0021 1.8027e-08 0 1.8141e-08 0 1.8144e-08 0.0021 1.8147e-08 0 1.8261e-08 0 1.8264e-08 0.0021 1.8267e-08 0 1.8381e-08 0 1.8384e-08 0.0021 1.8387e-08 0 1.8501e-08 0 1.8504e-08 0.0021 1.8507e-08 0 1.8621e-08 0 1.8624e-08 0.0021 1.8627e-08 0 1.8741e-08 0 1.8744e-08 0.0021 1.8747e-08 0 1.8861e-08 0 1.8864e-08 0.0021 1.8867e-08 0 1.8981e-08 0 1.8984e-08 0.0021 1.8987e-08 0 1.9101e-08 0 1.9104e-08 0.0021 1.9107e-08 0 1.9221e-08 0 1.9224e-08 0.0021 1.9227e-08 0 1.9341e-08 0 1.9344e-08 0.0021 1.9347e-08 0 1.9461e-08 0 1.9464e-08 0.0021 1.9467e-08 0 1.9581e-08 0 1.9584e-08 0.0021 1.9587e-08 0 1.9701e-08 0 1.9704e-08 0.0021 1.9707e-08 0 1.9821e-08 0 1.9824e-08 0.0021 1.9827e-08 0 1.9941e-08 0 1.9944e-08 0.0021 1.9947e-08 0 2.0061e-08 0 2.0064e-08 0.0021 2.0067e-08 0 2.0181e-08 0 2.0184e-08 0.0021 2.0187e-08 0 2.0301e-08 0 2.0304e-08 0.0021 2.0307e-08 0 2.0421e-08 0 2.0424e-08 0.0021 2.0427e-08 0 2.0541e-08 0 2.0544e-08 0.0021 2.0547e-08 0 2.0661e-08 0 2.0664e-08 0.0021 2.0667e-08 0 2.0781e-08 0 2.0784e-08 0.0021 2.0787e-08 0 2.0901e-08 0 2.0904e-08 0.0021 2.0907e-08 0 2.1021e-08 0 2.1024e-08 0.0021 2.1027e-08 0 2.1141e-08 0 2.1144e-08 0.0021 2.1147e-08 0 2.1261e-08 0 2.1264e-08 0.0021 2.1267e-08 0 2.1381e-08 0 2.1384e-08 0.0021 2.1387e-08 0 2.1501e-08 0 2.1504e-08 0.0021 2.1507e-08 0 2.1621e-08 0 2.1624e-08 0.0021 2.1627e-08 0 2.1741e-08 0 2.1744e-08 0.0021 2.1747e-08 0 2.1861e-08 0 2.1864e-08 0.0021 2.1867e-08 0 2.1981e-08 0 2.1984e-08 0.0021 2.1987e-08 0 2.2101e-08 0 2.2104e-08 0.0021 2.2107e-08 0 2.2221e-08 0 2.2224e-08 0.0021 2.2227e-08 0 2.2341e-08 0 2.2344e-08 0.0021 2.2347e-08 0 2.2461e-08 0 2.2464e-08 0.0021 2.2467e-08 0 2.2581e-08 0 2.2584e-08 0.0021 2.2587e-08 0 2.2701e-08 0 2.2704e-08 0.0021 2.2707e-08 0 2.2821e-08 0 2.2824e-08 0.0021 2.2827e-08 0 2.2941e-08 0 2.2944e-08 0.0021 2.2947e-08 0 2.3061e-08 0 2.3064e-08 0.0021 2.3067e-08 0 2.3181e-08 0 2.3184e-08 0.0021 2.3187e-08 0 2.3301e-08 0 2.3304e-08 0.0021 2.3307e-08 0 2.3421e-08 0 2.3424e-08 0.0021 2.3427e-08 0 2.3541e-08 0 2.3544e-08 0.0021 2.3547e-08 0 2.3661e-08 0 2.3664e-08 0.0021 2.3667e-08 0 2.3781e-08 0 2.3784e-08 0.0021 2.3787e-08 0 2.3901e-08 0 2.3904e-08 0.0021 2.3907e-08 0 2.4021e-08 0 2.4024e-08 0.0021 2.4027e-08 0 2.4141e-08 0 2.4144e-08 0.0021 2.4147e-08 0 2.4261e-08 0 2.4264e-08 0.0021 2.4267e-08 0 2.4381e-08 0 2.4384e-08 0.0021 2.4387e-08 0 2.4501e-08 0 2.4504e-08 0.0021 2.4507e-08 0 2.4621e-08 0 2.4624e-08 0.0021 2.4627e-08 0 2.4741e-08 0 2.4744e-08 0.0021 2.4747e-08 0 2.4861e-08 0 2.4864e-08 0.0021 2.4867e-08 0 2.4981e-08 0 2.4984e-08 0.0021 2.4987e-08 0 2.5101e-08 0 2.5104e-08 0.0021 2.5107e-08 0 2.5221e-08 0 2.5224e-08 0.0021 2.5227e-08 0 2.5341e-08 0 2.5344e-08 0.0021 2.5347e-08 0 2.5461e-08 0 2.5464e-08 0.0021 2.5467e-08 0 2.5581e-08 0 2.5584e-08 0.0021 2.5587e-08 0 2.5701e-08 0 2.5704e-08 0.0021 2.5707e-08 0 2.5821e-08 0 2.5824e-08 0.0021 2.5827e-08 0 2.5941e-08 0 2.5944e-08 0.0021 2.5947e-08 0 2.6061e-08 0 2.6064e-08 0.0021 2.6067e-08 0 2.6181e-08 0 2.6184e-08 0.0021 2.6187e-08 0 2.6301e-08 0 2.6304e-08 0.0021 2.6307e-08 0 2.6421e-08 0 2.6424e-08 0.0021 2.6427e-08 0 2.6541e-08 0 2.6544e-08 0.0021 2.6547e-08 0 2.6661e-08 0 2.6664e-08 0.0021 2.6667e-08 0 2.6781e-08 0 2.6784e-08 0.0021 2.6787e-08 0 2.6901e-08 0 2.6904e-08 0.0021 2.6907e-08 0 2.7021e-08 0 2.7024e-08 0.0021 2.7027e-08 0 2.7141e-08 0 2.7144e-08 0.0021 2.7147e-08 0 2.7261e-08 0 2.7264e-08 0.0021 2.7267e-08 0 2.7381e-08 0 2.7384e-08 0.0021 2.7387e-08 0 2.7501e-08 0 2.7504e-08 0.0021 2.7507e-08 0 2.7621e-08 0 2.7624e-08 0.0021 2.7627e-08 0 2.7741e-08 0 2.7744e-08 0.0021 2.7747e-08 0 2.7861e-08 0 2.7864e-08 0.0021 2.7867e-08 0 2.7981e-08 0 2.7984e-08 0.0021 2.7987e-08 0 2.8101e-08 0 2.8104e-08 0.0021 2.8107e-08 0 2.8221e-08 0 2.8224e-08 0.0021 2.8227e-08 0 2.8341e-08 0 2.8344e-08 0.0021 2.8347e-08 0 2.8461e-08 0 2.8464e-08 0.0021 2.8467e-08 0 2.8581e-08 0 2.8584e-08 0.0021 2.8587e-08 0 2.8701e-08 0 2.8704e-08 0.0021 2.8707e-08 0 2.8821e-08 0 2.8824e-08 0.0021 2.8827e-08 0 2.8941e-08 0 2.8944e-08 0.0021 2.8947e-08 0 2.9061e-08 0 2.9064e-08 0.0021 2.9067e-08 0 2.9181e-08 0 2.9184e-08 0.0021 2.9187e-08 0 2.9301e-08 0 2.9304e-08 0.0021 2.9307e-08 0 2.9421e-08 0 2.9424e-08 0.0021 2.9427e-08 0 2.9541e-08 0 2.9544e-08 0.0021 2.9547e-08 0 2.9661e-08 0 2.9664e-08 0.0021 2.9667e-08 0 2.9781e-08 0 2.9784e-08 0.0021 2.9787e-08 0 2.9901e-08 0 2.9904e-08 0.0021 2.9907e-08 0 3.0021e-08 0 3.0024e-08 0.0021 3.0027e-08 0 3.0141e-08 0 3.0144e-08 0.0021 3.0147e-08 0 3.0261e-08 0 3.0264e-08 0.0021 3.0267e-08 0 3.0381e-08 0 3.0384e-08 0.0021 3.0387e-08 0 3.0501e-08 0 3.0504e-08 0.0021 3.0507e-08 0 3.0621e-08 0 3.0624e-08 0.0021 3.0627e-08 0 3.0741e-08 0 3.0744e-08 0.0021 3.0747e-08 0 3.0861e-08 0 3.0864e-08 0.0021 3.0867e-08 0 3.0981e-08 0 3.0984e-08 0.0021 3.0987e-08 0 3.1101e-08 0 3.1104e-08 0.0021 3.1107e-08 0 3.1221e-08 0 3.1224e-08 0.0021 3.1227e-08 0 3.1341e-08 0 3.1344e-08 0.0021 3.1347e-08 0 3.1461e-08 0 3.1464e-08 0.0021 3.1467e-08 0 3.1581e-08 0 3.1584e-08 0.0021 3.1587e-08 0 3.1701e-08 0 3.1704e-08 0.0021 3.1707e-08 0 3.1821e-08 0 3.1824e-08 0.0021 3.1827e-08 0 3.1941e-08 0 3.1944e-08 0.0021 3.1947e-08 0 3.2061e-08 0 3.2064e-08 0.0021 3.2067e-08 0 3.2181e-08 0 3.2184e-08 0.0021 3.2187e-08 0 3.2301e-08 0 3.2304e-08 0.0021 3.2307e-08 0 3.2421e-08 0 3.2424e-08 0.0021 3.2427e-08 0 3.2541e-08 0 3.2544e-08 0.0021 3.2547e-08 0 3.2661e-08 0 3.2664e-08 0.0021 3.2667e-08 0 3.2781e-08 0 3.2784e-08 0.0021 3.2787e-08 0 3.2901e-08 0 3.2904e-08 0.0021 3.2907e-08 0 3.3021e-08 0 3.3024e-08 0.0021 3.3027e-08 0 3.3141e-08 0 3.3144e-08 0.0021 3.3147e-08 0 3.3261e-08 0 3.3264e-08 0.0021 3.3267e-08 0 3.3381e-08 0 3.3384e-08 0.0021 3.3387e-08 0 3.3501e-08 0 3.3504e-08 0.0021 3.3507e-08 0 3.3621e-08 0 3.3624e-08 0.0021 3.3627e-08 0 3.3741e-08 0 3.3744e-08 0.0021 3.3747e-08 0 3.3861e-08 0 3.3864e-08 0.0021 3.3867e-08 0 3.3981e-08 0 3.3984e-08 0.0021 3.3987e-08 0 3.4101e-08 0 3.4104e-08 0.0021 3.4107e-08 0 3.4221e-08 0 3.4224e-08 0.0021 3.4227e-08 0 3.4341e-08 0 3.4344e-08 0.0021 3.4347e-08 0 3.4461e-08 0 3.4464e-08 0.0021 3.4467e-08 0 3.4581e-08 0 3.4584e-08 0.0021 3.4587e-08 0 3.4701e-08 0 3.4704e-08 0.0021 3.4707e-08 0 3.4821e-08 0 3.4824e-08 0.0021 3.4827e-08 0 3.4941e-08 0 3.4944e-08 0.0021 3.4947e-08 0 3.5061e-08 0 3.5064e-08 0.0021 3.5067e-08 0 3.5181e-08 0 3.5184e-08 0.0021 3.5187e-08 0 3.5301e-08 0 3.5304e-08 0.0021 3.5307e-08 0 3.5421e-08 0 3.5424e-08 0.0021 3.5427e-08 0 3.5541e-08 0 3.5544e-08 0.0021 3.5547e-08 0 3.5661e-08 0 3.5664e-08 0.0021 3.5667e-08 0 3.5781e-08 0 3.5784e-08 0.0021 3.5787e-08 0 3.5901e-08 0 3.5904e-08 0.0021 3.5907e-08 0 3.6021e-08 0 3.6024e-08 0.0021 3.6027e-08 0 3.6141e-08 0 3.6144e-08 0.0021 3.6147e-08 0 3.6261e-08 0 3.6264e-08 0.0021 3.6267e-08 0 3.6381e-08 0 3.6384e-08 0.0021 3.6387e-08 0 3.6501e-08 0 3.6504e-08 0.0021 3.6507e-08 0 3.6621e-08 0 3.6624e-08 0.0021 3.6627e-08 0 3.6741e-08 0 3.6744e-08 0.0021 3.6747e-08 0 3.6861e-08 0 3.6864e-08 0.0021 3.6867e-08 0 3.6981e-08 0 3.6984e-08 0.0021 3.6987e-08 0 3.7101e-08 0 3.7104e-08 0.0021 3.7107e-08 0 3.7221e-08 0 3.7224e-08 0.0021 3.7227e-08 0 3.7341e-08 0 3.7344e-08 0.0021 3.7347e-08 0 3.7461e-08 0 3.7464e-08 0.0021 3.7467e-08 0 3.7581e-08 0 3.7584e-08 0.0021 3.7587e-08 0 3.7701e-08 0 3.7704e-08 0.0021 3.7707e-08 0 3.7821e-08 0 3.7824e-08 0.0021 3.7827e-08 0 3.7941e-08 0 3.7944e-08 0.0021 3.7947e-08 0 3.8061e-08 0 3.8064e-08 0.0021 3.8067e-08 0 3.8181e-08 0 3.8184e-08 0.0021 3.8187e-08 0 3.8301e-08 0 3.8304e-08 0.0021 3.8307e-08 0 3.8421e-08 0 3.8424e-08 0.0021 3.8427e-08 0 3.8541e-08 0 3.8544e-08 0.0021 3.8547e-08 0 3.8661e-08 0 3.8664e-08 0.0021 3.8667e-08 0 3.8781e-08 0 3.8784e-08 0.0021 3.8787e-08 0 3.8901e-08 0 3.8904e-08 0.0021 3.8907e-08 0 3.9021e-08 0 3.9024e-08 0.0021 3.9027e-08 0 3.9141e-08 0 3.9144e-08 0.0021 3.9147e-08 0 3.9261e-08 0 3.9264e-08 0.0021 3.9267e-08 0 3.9381e-08 0 3.9384e-08 0.0021 3.9387e-08 0 3.9501e-08 0 3.9504e-08 0.0021 3.9507e-08 0 3.9621e-08 0 3.9624e-08 0.0021 3.9627e-08 0 3.9741e-08 0 3.9744e-08 0.0021 3.9747e-08 0 3.9861e-08 0 3.9864e-08 0.0021 3.9867e-08 0 3.9981e-08 0 3.9984e-08 0.0021 3.9987e-08 0 4.0101e-08 0 4.0104e-08 0.0021 4.0107e-08 0 4.0221e-08 0 4.0224e-08 0.0021 4.0227e-08 0 4.0341e-08 0 4.0344e-08 0.0021 4.0347e-08 0 4.0461e-08 0 4.0464e-08 0.0021 4.0467e-08 0 4.0581e-08 0 4.0584e-08 0.0021 4.0587e-08 0 4.0701e-08 0 4.0704e-08 0.0021 4.0707e-08 0 4.0821e-08 0 4.0824e-08 0.0021 4.0827e-08 0 4.0941e-08 0 4.0944e-08 0.0021 4.0947e-08 0 4.1061e-08 0 4.1064e-08 0.0021 4.1067e-08 0 4.1181e-08 0 4.1184e-08 0.0021 4.1187e-08 0 4.1301e-08 0 4.1304e-08 0.0021 4.1307e-08 0 4.1421e-08 0 4.1424e-08 0.0021 4.1427e-08 0 4.1541e-08 0 4.1544e-08 0.0021 4.1547e-08 0 4.1661e-08 0 4.1664e-08 0.0021 4.1667e-08 0 4.1781e-08 0 4.1784e-08 0.0021 4.1787e-08 0 4.1901e-08 0 4.1904e-08 0.0021 4.1907e-08 0 4.2021e-08 0 4.2024e-08 0.0021 4.2027e-08 0 4.2141e-08 0 4.2144e-08 0.0021 4.2147e-08 0 4.2261e-08 0 4.2264e-08 0.0021 4.2267e-08 0 4.2381e-08 0 4.2384e-08 0.0021 4.2387e-08 0 4.2501e-08 0 4.2504e-08 0.0021 4.2507e-08 0 4.2621e-08 0 4.2624e-08 0.0021 4.2627e-08 0 4.2741e-08 0 4.2744e-08 0.0021 4.2747e-08 0 4.2861e-08 0 4.2864e-08 0.0021 4.2867e-08 0 4.2981e-08 0 4.2984e-08 0.0021 4.2987e-08 0 4.3101e-08 0 4.3104e-08 0.0021 4.3107e-08 0 4.3221e-08 0 4.3224e-08 0.0021 4.3227e-08 0 4.3341e-08 0 4.3344e-08 0.0021 4.3347e-08 0 4.3461e-08 0 4.3464e-08 0.0021 4.3467e-08 0 4.3581e-08 0 4.3584e-08 0.0021 4.3587e-08 0 4.3701e-08 0 4.3704e-08 0.0021 4.3707e-08 0 4.3821e-08 0 4.3824e-08 0.0021 4.3827e-08 0 4.3941e-08 0 4.3944e-08 0.0021 4.3947e-08 0 4.4061e-08 0 4.4064e-08 0.0021 4.4067e-08 0 4.4181e-08 0 4.4184e-08 0.0021 4.4187e-08 0 4.4301e-08 0 4.4304e-08 0.0021 4.4307e-08 0 4.4421e-08 0 4.4424e-08 0.0021 4.4427e-08 0 4.4541e-08 0 4.4544e-08 0.0021 4.4547e-08 0 4.4661e-08 0 4.4664e-08 0.0021 4.4667e-08 0 4.4781e-08 0 4.4784e-08 0.0021 4.4787e-08 0 4.4901e-08 0 4.4904e-08 0.0021 4.4907e-08 0 4.5021e-08 0 4.5024e-08 0.0021 4.5027e-08 0 4.5141e-08 0 4.5144e-08 0.0021 4.5147e-08 0 4.5261e-08 0 4.5264e-08 0.0021 4.5267e-08 0 4.5381e-08 0 4.5384e-08 0.0021 4.5387e-08 0 4.5501e-08 0 4.5504e-08 0.0021 4.5507e-08 0 4.5621e-08 0 4.5624e-08 0.0021 4.5627e-08 0 4.5741e-08 0 4.5744e-08 0.0021 4.5747e-08 0 4.5861e-08 0 4.5864e-08 0.0021 4.5867e-08 0 4.5981e-08 0 4.5984e-08 0.0021 4.5987e-08 0 4.6101e-08 0 4.6104e-08 0.0021 4.6107e-08 0 4.6221e-08 0 4.6224e-08 0.0021 4.6227e-08 0 4.6341e-08 0 4.6344e-08 0.0021 4.6347e-08 0 4.6461e-08 0 4.6464e-08 0.0021 4.6467e-08 0 4.6581e-08 0 4.6584e-08 0.0021 4.6587e-08 0 4.6701e-08 0 4.6704e-08 0.0021 4.6707e-08 0 4.6821e-08 0 4.6824e-08 0.0021 4.6827e-08 0 4.6941e-08 0 4.6944e-08 0.0021 4.6947e-08 0 4.7061e-08 0 4.7064e-08 0.0021 4.7067e-08 0 4.7181e-08 0 4.7184e-08 0.0021 4.7187e-08 0 4.7301e-08 0 4.7304e-08 0.0021 4.7307e-08 0 4.7421e-08 0 4.7424e-08 0.0021 4.7427e-08 0 4.7541e-08 0 4.7544e-08 0.0021 4.7547e-08 0 4.7661e-08 0 4.7664e-08 0.0021 4.7667e-08 0 4.7781e-08 0 4.7784e-08 0.0021 4.7787e-08 0)
IT02|T 0 T02  PWL(0 0 2.1e-11 0 2.4e-11 0.0021 2.7e-11 0 1.41e-10 0 1.44e-10 0.0021 1.47e-10 0 2.61e-10 0 2.64e-10 0.0021 2.67e-10 0 3.81e-10 0 3.84e-10 0.0021 3.87e-10 0 5.01e-10 0 5.04e-10 0.0021 5.07e-10 0 6.21e-10 0 6.24e-10 0.0021 6.27e-10 0 7.41e-10 0 7.44e-10 0.0021 7.47e-10 0 8.61e-10 0 8.64e-10 0.0021 8.67e-10 0 9.81e-10 0 9.84e-10 0.0021 9.87e-10 0 1.101e-09 0 1.104e-09 0.0021 1.107e-09 0 1.221e-09 0 1.224e-09 0.0021 1.227e-09 0 1.341e-09 0 1.344e-09 0.0021 1.347e-09 0 1.461e-09 0 1.464e-09 0.0021 1.467e-09 0 1.581e-09 0 1.584e-09 0.0021 1.587e-09 0 1.701e-09 0 1.704e-09 0.0021 1.707e-09 0 1.821e-09 0 1.824e-09 0.0021 1.827e-09 0 1.941e-09 0 1.944e-09 0.0021 1.947e-09 0 2.061e-09 0 2.064e-09 0.0021 2.067e-09 0 2.181e-09 0 2.184e-09 0.0021 2.187e-09 0 2.301e-09 0 2.304e-09 0.0021 2.307e-09 0 2.421e-09 0 2.424e-09 0.0021 2.427e-09 0 2.541e-09 0 2.544e-09 0.0021 2.547e-09 0 2.661e-09 0 2.664e-09 0.0021 2.667e-09 0 2.781e-09 0 2.784e-09 0.0021 2.787e-09 0 2.901e-09 0 2.904e-09 0.0021 2.907e-09 0 3.021e-09 0 3.024e-09 0.0021 3.027e-09 0 3.141e-09 0 3.144e-09 0.0021 3.147e-09 0 3.261e-09 0 3.264e-09 0.0021 3.267e-09 0 3.381e-09 0 3.384e-09 0.0021 3.387e-09 0 3.501e-09 0 3.504e-09 0.0021 3.507e-09 0 3.621e-09 0 3.624e-09 0.0021 3.627e-09 0 3.741e-09 0 3.744e-09 0.0021 3.747e-09 0 3.861e-09 0 3.864e-09 0.0021 3.867e-09 0 3.981e-09 0 3.984e-09 0.0021 3.987e-09 0 4.101e-09 0 4.104e-09 0.0021 4.107e-09 0 4.221e-09 0 4.224e-09 0.0021 4.227e-09 0 4.341e-09 0 4.344e-09 0.0021 4.347e-09 0 4.461e-09 0 4.464e-09 0.0021 4.467e-09 0 4.581e-09 0 4.584e-09 0.0021 4.587e-09 0 4.701e-09 0 4.704e-09 0.0021 4.707e-09 0 4.821e-09 0 4.824e-09 0.0021 4.827e-09 0 4.941e-09 0 4.944e-09 0.0021 4.947e-09 0 5.061e-09 0 5.064e-09 0.0021 5.067e-09 0 5.181e-09 0 5.184e-09 0.0021 5.187e-09 0 5.301e-09 0 5.304e-09 0.0021 5.307e-09 0 5.421e-09 0 5.424e-09 0.0021 5.427e-09 0 5.541e-09 0 5.544e-09 0.0021 5.547e-09 0 5.661e-09 0 5.664e-09 0.0021 5.667e-09 0 5.781e-09 0 5.784e-09 0.0021 5.787e-09 0 5.901e-09 0 5.904e-09 0.0021 5.907e-09 0 6.021e-09 0 6.024e-09 0.0021 6.027e-09 0 6.141e-09 0 6.144e-09 0.0021 6.147e-09 0 6.261e-09 0 6.264e-09 0.0021 6.267e-09 0 6.381e-09 0 6.384e-09 0.0021 6.387e-09 0 6.501e-09 0 6.504e-09 0.0021 6.507e-09 0 6.621e-09 0 6.624e-09 0.0021 6.627e-09 0 6.741e-09 0 6.744e-09 0.0021 6.747e-09 0 6.861e-09 0 6.864e-09 0.0021 6.867e-09 0 6.981e-09 0 6.984e-09 0.0021 6.987e-09 0 7.101e-09 0 7.104e-09 0.0021 7.107e-09 0 7.221e-09 0 7.224e-09 0.0021 7.227e-09 0 7.341e-09 0 7.344e-09 0.0021 7.347e-09 0 7.461e-09 0 7.464e-09 0.0021 7.467e-09 0 7.581e-09 0 7.584e-09 0.0021 7.587e-09 0 7.701e-09 0 7.704e-09 0.0021 7.707e-09 0 7.821e-09 0 7.824e-09 0.0021 7.827e-09 0 7.941e-09 0 7.944e-09 0.0021 7.947e-09 0 8.061e-09 0 8.064e-09 0.0021 8.067e-09 0 8.181e-09 0 8.184e-09 0.0021 8.187e-09 0 8.301e-09 0 8.304e-09 0.0021 8.307e-09 0 8.421e-09 0 8.424e-09 0.0021 8.427e-09 0 8.541e-09 0 8.544e-09 0.0021 8.547e-09 0 8.661e-09 0 8.664e-09 0.0021 8.667e-09 0 8.781e-09 0 8.784e-09 0.0021 8.787e-09 0 8.901e-09 0 8.904e-09 0.0021 8.907e-09 0 9.021e-09 0 9.024e-09 0.0021 9.027e-09 0 9.141e-09 0 9.144e-09 0.0021 9.147e-09 0 9.261e-09 0 9.264e-09 0.0021 9.267e-09 0 9.381e-09 0 9.384e-09 0.0021 9.387e-09 0 9.501e-09 0 9.504e-09 0.0021 9.507e-09 0 9.621e-09 0 9.624e-09 0.0021 9.627e-09 0 9.741e-09 0 9.744e-09 0.0021 9.747e-09 0 9.861e-09 0 9.864e-09 0.0021 9.867e-09 0 9.981e-09 0 9.984e-09 0.0021 9.987e-09 0 1.0101e-08 0 1.0104e-08 0.0021 1.0107e-08 0 1.0221e-08 0 1.0224e-08 0.0021 1.0227e-08 0 1.0341e-08 0 1.0344e-08 0.0021 1.0347e-08 0 1.0461e-08 0 1.0464e-08 0.0021 1.0467e-08 0 1.0581e-08 0 1.0584e-08 0.0021 1.0587e-08 0 1.0701e-08 0 1.0704e-08 0.0021 1.0707e-08 0 1.0821e-08 0 1.0824e-08 0.0021 1.0827e-08 0 1.0941e-08 0 1.0944e-08 0.0021 1.0947e-08 0 1.1061e-08 0 1.1064e-08 0.0021 1.1067e-08 0 1.1181e-08 0 1.1184e-08 0.0021 1.1187e-08 0 1.1301e-08 0 1.1304e-08 0.0021 1.1307e-08 0 1.1421e-08 0 1.1424e-08 0.0021 1.1427e-08 0 1.1541e-08 0 1.1544e-08 0.0021 1.1547e-08 0 1.1661e-08 0 1.1664e-08 0.0021 1.1667e-08 0 1.1781e-08 0 1.1784e-08 0.0021 1.1787e-08 0 1.1901e-08 0 1.1904e-08 0.0021 1.1907e-08 0 1.2021e-08 0 1.2024e-08 0.0021 1.2027e-08 0 1.2141e-08 0 1.2144e-08 0.0021 1.2147e-08 0 1.2261e-08 0 1.2264e-08 0.0021 1.2267e-08 0 1.2381e-08 0 1.2384e-08 0.0021 1.2387e-08 0 1.2501e-08 0 1.2504e-08 0.0021 1.2507e-08 0 1.2621e-08 0 1.2624e-08 0.0021 1.2627e-08 0 1.2741e-08 0 1.2744e-08 0.0021 1.2747e-08 0 1.2861e-08 0 1.2864e-08 0.0021 1.2867e-08 0 1.2981e-08 0 1.2984e-08 0.0021 1.2987e-08 0 1.3101e-08 0 1.3104e-08 0.0021 1.3107e-08 0 1.3221e-08 0 1.3224e-08 0.0021 1.3227e-08 0 1.3341e-08 0 1.3344e-08 0.0021 1.3347e-08 0 1.3461e-08 0 1.3464e-08 0.0021 1.3467e-08 0 1.3581e-08 0 1.3584e-08 0.0021 1.3587e-08 0 1.3701e-08 0 1.3704e-08 0.0021 1.3707e-08 0 1.3821e-08 0 1.3824e-08 0.0021 1.3827e-08 0 1.3941e-08 0 1.3944e-08 0.0021 1.3947e-08 0 1.4061e-08 0 1.4064e-08 0.0021 1.4067e-08 0 1.4181e-08 0 1.4184e-08 0.0021 1.4187e-08 0 1.4301e-08 0 1.4304e-08 0.0021 1.4307e-08 0 1.4421e-08 0 1.4424e-08 0.0021 1.4427e-08 0 1.4541e-08 0 1.4544e-08 0.0021 1.4547e-08 0 1.4661e-08 0 1.4664e-08 0.0021 1.4667e-08 0 1.4781e-08 0 1.4784e-08 0.0021 1.4787e-08 0 1.4901e-08 0 1.4904e-08 0.0021 1.4907e-08 0 1.5021e-08 0 1.5024e-08 0.0021 1.5027e-08 0 1.5141e-08 0 1.5144e-08 0.0021 1.5147e-08 0 1.5261e-08 0 1.5264e-08 0.0021 1.5267e-08 0 1.5381e-08 0 1.5384e-08 0.0021 1.5387e-08 0 1.5501e-08 0 1.5504e-08 0.0021 1.5507e-08 0 1.5621e-08 0 1.5624e-08 0.0021 1.5627e-08 0 1.5741e-08 0 1.5744e-08 0.0021 1.5747e-08 0 1.5861e-08 0 1.5864e-08 0.0021 1.5867e-08 0 1.5981e-08 0 1.5984e-08 0.0021 1.5987e-08 0 1.6101e-08 0 1.6104e-08 0.0021 1.6107e-08 0 1.6221e-08 0 1.6224e-08 0.0021 1.6227e-08 0 1.6341e-08 0 1.6344e-08 0.0021 1.6347e-08 0 1.6461e-08 0 1.6464e-08 0.0021 1.6467e-08 0 1.6581e-08 0 1.6584e-08 0.0021 1.6587e-08 0 1.6701e-08 0 1.6704e-08 0.0021 1.6707e-08 0 1.6821e-08 0 1.6824e-08 0.0021 1.6827e-08 0 1.6941e-08 0 1.6944e-08 0.0021 1.6947e-08 0 1.7061e-08 0 1.7064e-08 0.0021 1.7067e-08 0 1.7181e-08 0 1.7184e-08 0.0021 1.7187e-08 0 1.7301e-08 0 1.7304e-08 0.0021 1.7307e-08 0 1.7421e-08 0 1.7424e-08 0.0021 1.7427e-08 0 1.7541e-08 0 1.7544e-08 0.0021 1.7547e-08 0 1.7661e-08 0 1.7664e-08 0.0021 1.7667e-08 0 1.7781e-08 0 1.7784e-08 0.0021 1.7787e-08 0 1.7901e-08 0 1.7904e-08 0.0021 1.7907e-08 0 1.8021e-08 0 1.8024e-08 0.0021 1.8027e-08 0 1.8141e-08 0 1.8144e-08 0.0021 1.8147e-08 0 1.8261e-08 0 1.8264e-08 0.0021 1.8267e-08 0 1.8381e-08 0 1.8384e-08 0.0021 1.8387e-08 0 1.8501e-08 0 1.8504e-08 0.0021 1.8507e-08 0 1.8621e-08 0 1.8624e-08 0.0021 1.8627e-08 0 1.8741e-08 0 1.8744e-08 0.0021 1.8747e-08 0 1.8861e-08 0 1.8864e-08 0.0021 1.8867e-08 0 1.8981e-08 0 1.8984e-08 0.0021 1.8987e-08 0 1.9101e-08 0 1.9104e-08 0.0021 1.9107e-08 0 1.9221e-08 0 1.9224e-08 0.0021 1.9227e-08 0 1.9341e-08 0 1.9344e-08 0.0021 1.9347e-08 0 1.9461e-08 0 1.9464e-08 0.0021 1.9467e-08 0 1.9581e-08 0 1.9584e-08 0.0021 1.9587e-08 0 1.9701e-08 0 1.9704e-08 0.0021 1.9707e-08 0 1.9821e-08 0 1.9824e-08 0.0021 1.9827e-08 0 1.9941e-08 0 1.9944e-08 0.0021 1.9947e-08 0 2.0061e-08 0 2.0064e-08 0.0021 2.0067e-08 0 2.0181e-08 0 2.0184e-08 0.0021 2.0187e-08 0 2.0301e-08 0 2.0304e-08 0.0021 2.0307e-08 0 2.0421e-08 0 2.0424e-08 0.0021 2.0427e-08 0 2.0541e-08 0 2.0544e-08 0.0021 2.0547e-08 0 2.0661e-08 0 2.0664e-08 0.0021 2.0667e-08 0 2.0781e-08 0 2.0784e-08 0.0021 2.0787e-08 0 2.0901e-08 0 2.0904e-08 0.0021 2.0907e-08 0 2.1021e-08 0 2.1024e-08 0.0021 2.1027e-08 0 2.1141e-08 0 2.1144e-08 0.0021 2.1147e-08 0 2.1261e-08 0 2.1264e-08 0.0021 2.1267e-08 0 2.1381e-08 0 2.1384e-08 0.0021 2.1387e-08 0 2.1501e-08 0 2.1504e-08 0.0021 2.1507e-08 0 2.1621e-08 0 2.1624e-08 0.0021 2.1627e-08 0 2.1741e-08 0 2.1744e-08 0.0021 2.1747e-08 0 2.1861e-08 0 2.1864e-08 0.0021 2.1867e-08 0 2.1981e-08 0 2.1984e-08 0.0021 2.1987e-08 0 2.2101e-08 0 2.2104e-08 0.0021 2.2107e-08 0 2.2221e-08 0 2.2224e-08 0.0021 2.2227e-08 0 2.2341e-08 0 2.2344e-08 0.0021 2.2347e-08 0 2.2461e-08 0 2.2464e-08 0.0021 2.2467e-08 0 2.2581e-08 0 2.2584e-08 0.0021 2.2587e-08 0 2.2701e-08 0 2.2704e-08 0.0021 2.2707e-08 0 2.2821e-08 0 2.2824e-08 0.0021 2.2827e-08 0 2.2941e-08 0 2.2944e-08 0.0021 2.2947e-08 0 2.3061e-08 0 2.3064e-08 0.0021 2.3067e-08 0 2.3181e-08 0 2.3184e-08 0.0021 2.3187e-08 0 2.3301e-08 0 2.3304e-08 0.0021 2.3307e-08 0 2.3421e-08 0 2.3424e-08 0.0021 2.3427e-08 0 2.3541e-08 0 2.3544e-08 0.0021 2.3547e-08 0 2.3661e-08 0 2.3664e-08 0.0021 2.3667e-08 0 2.3781e-08 0 2.3784e-08 0.0021 2.3787e-08 0 2.3901e-08 0 2.3904e-08 0.0021 2.3907e-08 0 2.4021e-08 0 2.4024e-08 0.0021 2.4027e-08 0 2.4141e-08 0 2.4144e-08 0.0021 2.4147e-08 0 2.4261e-08 0 2.4264e-08 0.0021 2.4267e-08 0 2.4381e-08 0 2.4384e-08 0.0021 2.4387e-08 0 2.4501e-08 0 2.4504e-08 0.0021 2.4507e-08 0 2.4621e-08 0 2.4624e-08 0.0021 2.4627e-08 0 2.4741e-08 0 2.4744e-08 0.0021 2.4747e-08 0 2.4861e-08 0 2.4864e-08 0.0021 2.4867e-08 0 2.4981e-08 0 2.4984e-08 0.0021 2.4987e-08 0 2.5101e-08 0 2.5104e-08 0.0021 2.5107e-08 0 2.5221e-08 0 2.5224e-08 0.0021 2.5227e-08 0 2.5341e-08 0 2.5344e-08 0.0021 2.5347e-08 0 2.5461e-08 0 2.5464e-08 0.0021 2.5467e-08 0 2.5581e-08 0 2.5584e-08 0.0021 2.5587e-08 0 2.5701e-08 0 2.5704e-08 0.0021 2.5707e-08 0 2.5821e-08 0 2.5824e-08 0.0021 2.5827e-08 0 2.5941e-08 0 2.5944e-08 0.0021 2.5947e-08 0 2.6061e-08 0 2.6064e-08 0.0021 2.6067e-08 0 2.6181e-08 0 2.6184e-08 0.0021 2.6187e-08 0 2.6301e-08 0 2.6304e-08 0.0021 2.6307e-08 0 2.6421e-08 0 2.6424e-08 0.0021 2.6427e-08 0 2.6541e-08 0 2.6544e-08 0.0021 2.6547e-08 0 2.6661e-08 0 2.6664e-08 0.0021 2.6667e-08 0 2.6781e-08 0 2.6784e-08 0.0021 2.6787e-08 0 2.6901e-08 0 2.6904e-08 0.0021 2.6907e-08 0 2.7021e-08 0 2.7024e-08 0.0021 2.7027e-08 0 2.7141e-08 0 2.7144e-08 0.0021 2.7147e-08 0 2.7261e-08 0 2.7264e-08 0.0021 2.7267e-08 0 2.7381e-08 0 2.7384e-08 0.0021 2.7387e-08 0 2.7501e-08 0 2.7504e-08 0.0021 2.7507e-08 0 2.7621e-08 0 2.7624e-08 0.0021 2.7627e-08 0 2.7741e-08 0 2.7744e-08 0.0021 2.7747e-08 0 2.7861e-08 0 2.7864e-08 0.0021 2.7867e-08 0 2.7981e-08 0 2.7984e-08 0.0021 2.7987e-08 0 2.8101e-08 0 2.8104e-08 0.0021 2.8107e-08 0 2.8221e-08 0 2.8224e-08 0.0021 2.8227e-08 0 2.8341e-08 0 2.8344e-08 0.0021 2.8347e-08 0 2.8461e-08 0 2.8464e-08 0.0021 2.8467e-08 0 2.8581e-08 0 2.8584e-08 0.0021 2.8587e-08 0 2.8701e-08 0 2.8704e-08 0.0021 2.8707e-08 0 2.8821e-08 0 2.8824e-08 0.0021 2.8827e-08 0 2.8941e-08 0 2.8944e-08 0.0021 2.8947e-08 0 2.9061e-08 0 2.9064e-08 0.0021 2.9067e-08 0 2.9181e-08 0 2.9184e-08 0.0021 2.9187e-08 0 2.9301e-08 0 2.9304e-08 0.0021 2.9307e-08 0 2.9421e-08 0 2.9424e-08 0.0021 2.9427e-08 0 2.9541e-08 0 2.9544e-08 0.0021 2.9547e-08 0 2.9661e-08 0 2.9664e-08 0.0021 2.9667e-08 0 2.9781e-08 0 2.9784e-08 0.0021 2.9787e-08 0 2.9901e-08 0 2.9904e-08 0.0021 2.9907e-08 0 3.0021e-08 0 3.0024e-08 0.0021 3.0027e-08 0 3.0141e-08 0 3.0144e-08 0.0021 3.0147e-08 0 3.0261e-08 0 3.0264e-08 0.0021 3.0267e-08 0 3.0381e-08 0 3.0384e-08 0.0021 3.0387e-08 0 3.0501e-08 0 3.0504e-08 0.0021 3.0507e-08 0 3.0621e-08 0 3.0624e-08 0.0021 3.0627e-08 0 3.0741e-08 0 3.0744e-08 0.0021 3.0747e-08 0 3.0861e-08 0 3.0864e-08 0.0021 3.0867e-08 0 3.0981e-08 0 3.0984e-08 0.0021 3.0987e-08 0 3.1101e-08 0 3.1104e-08 0.0021 3.1107e-08 0 3.1221e-08 0 3.1224e-08 0.0021 3.1227e-08 0 3.1341e-08 0 3.1344e-08 0.0021 3.1347e-08 0 3.1461e-08 0 3.1464e-08 0.0021 3.1467e-08 0 3.1581e-08 0 3.1584e-08 0.0021 3.1587e-08 0 3.1701e-08 0 3.1704e-08 0.0021 3.1707e-08 0 3.1821e-08 0 3.1824e-08 0.0021 3.1827e-08 0 3.1941e-08 0 3.1944e-08 0.0021 3.1947e-08 0 3.2061e-08 0 3.2064e-08 0.0021 3.2067e-08 0 3.2181e-08 0 3.2184e-08 0.0021 3.2187e-08 0 3.2301e-08 0 3.2304e-08 0.0021 3.2307e-08 0 3.2421e-08 0 3.2424e-08 0.0021 3.2427e-08 0 3.2541e-08 0 3.2544e-08 0.0021 3.2547e-08 0 3.2661e-08 0 3.2664e-08 0.0021 3.2667e-08 0 3.2781e-08 0 3.2784e-08 0.0021 3.2787e-08 0 3.2901e-08 0 3.2904e-08 0.0021 3.2907e-08 0 3.3021e-08 0 3.3024e-08 0.0021 3.3027e-08 0 3.3141e-08 0 3.3144e-08 0.0021 3.3147e-08 0 3.3261e-08 0 3.3264e-08 0.0021 3.3267e-08 0 3.3381e-08 0 3.3384e-08 0.0021 3.3387e-08 0 3.3501e-08 0 3.3504e-08 0.0021 3.3507e-08 0 3.3621e-08 0 3.3624e-08 0.0021 3.3627e-08 0 3.3741e-08 0 3.3744e-08 0.0021 3.3747e-08 0 3.3861e-08 0 3.3864e-08 0.0021 3.3867e-08 0 3.3981e-08 0 3.3984e-08 0.0021 3.3987e-08 0 3.4101e-08 0 3.4104e-08 0.0021 3.4107e-08 0 3.4221e-08 0 3.4224e-08 0.0021 3.4227e-08 0 3.4341e-08 0 3.4344e-08 0.0021 3.4347e-08 0 3.4461e-08 0 3.4464e-08 0.0021 3.4467e-08 0 3.4581e-08 0 3.4584e-08 0.0021 3.4587e-08 0 3.4701e-08 0 3.4704e-08 0.0021 3.4707e-08 0 3.4821e-08 0 3.4824e-08 0.0021 3.4827e-08 0 3.4941e-08 0 3.4944e-08 0.0021 3.4947e-08 0 3.5061e-08 0 3.5064e-08 0.0021 3.5067e-08 0 3.5181e-08 0 3.5184e-08 0.0021 3.5187e-08 0 3.5301e-08 0 3.5304e-08 0.0021 3.5307e-08 0 3.5421e-08 0 3.5424e-08 0.0021 3.5427e-08 0 3.5541e-08 0 3.5544e-08 0.0021 3.5547e-08 0 3.5661e-08 0 3.5664e-08 0.0021 3.5667e-08 0 3.5781e-08 0 3.5784e-08 0.0021 3.5787e-08 0 3.5901e-08 0 3.5904e-08 0.0021 3.5907e-08 0 3.6021e-08 0 3.6024e-08 0.0021 3.6027e-08 0 3.6141e-08 0 3.6144e-08 0.0021 3.6147e-08 0 3.6261e-08 0 3.6264e-08 0.0021 3.6267e-08 0 3.6381e-08 0 3.6384e-08 0.0021 3.6387e-08 0 3.6501e-08 0 3.6504e-08 0.0021 3.6507e-08 0 3.6621e-08 0 3.6624e-08 0.0021 3.6627e-08 0 3.6741e-08 0 3.6744e-08 0.0021 3.6747e-08 0 3.6861e-08 0 3.6864e-08 0.0021 3.6867e-08 0 3.6981e-08 0 3.6984e-08 0.0021 3.6987e-08 0 3.7101e-08 0 3.7104e-08 0.0021 3.7107e-08 0 3.7221e-08 0 3.7224e-08 0.0021 3.7227e-08 0 3.7341e-08 0 3.7344e-08 0.0021 3.7347e-08 0 3.7461e-08 0 3.7464e-08 0.0021 3.7467e-08 0 3.7581e-08 0 3.7584e-08 0.0021 3.7587e-08 0 3.7701e-08 0 3.7704e-08 0.0021 3.7707e-08 0 3.7821e-08 0 3.7824e-08 0.0021 3.7827e-08 0 3.7941e-08 0 3.7944e-08 0.0021 3.7947e-08 0 3.8061e-08 0 3.8064e-08 0.0021 3.8067e-08 0 3.8181e-08 0 3.8184e-08 0.0021 3.8187e-08 0 3.8301e-08 0 3.8304e-08 0.0021 3.8307e-08 0 3.8421e-08 0 3.8424e-08 0.0021 3.8427e-08 0 3.8541e-08 0 3.8544e-08 0.0021 3.8547e-08 0 3.8661e-08 0 3.8664e-08 0.0021 3.8667e-08 0 3.8781e-08 0 3.8784e-08 0.0021 3.8787e-08 0 3.8901e-08 0 3.8904e-08 0.0021 3.8907e-08 0 3.9021e-08 0 3.9024e-08 0.0021 3.9027e-08 0 3.9141e-08 0 3.9144e-08 0.0021 3.9147e-08 0 3.9261e-08 0 3.9264e-08 0.0021 3.9267e-08 0 3.9381e-08 0 3.9384e-08 0.0021 3.9387e-08 0 3.9501e-08 0 3.9504e-08 0.0021 3.9507e-08 0 3.9621e-08 0 3.9624e-08 0.0021 3.9627e-08 0 3.9741e-08 0 3.9744e-08 0.0021 3.9747e-08 0 3.9861e-08 0 3.9864e-08 0.0021 3.9867e-08 0 3.9981e-08 0 3.9984e-08 0.0021 3.9987e-08 0 4.0101e-08 0 4.0104e-08 0.0021 4.0107e-08 0 4.0221e-08 0 4.0224e-08 0.0021 4.0227e-08 0 4.0341e-08 0 4.0344e-08 0.0021 4.0347e-08 0 4.0461e-08 0 4.0464e-08 0.0021 4.0467e-08 0 4.0581e-08 0 4.0584e-08 0.0021 4.0587e-08 0 4.0701e-08 0 4.0704e-08 0.0021 4.0707e-08 0 4.0821e-08 0 4.0824e-08 0.0021 4.0827e-08 0 4.0941e-08 0 4.0944e-08 0.0021 4.0947e-08 0 4.1061e-08 0 4.1064e-08 0.0021 4.1067e-08 0 4.1181e-08 0 4.1184e-08 0.0021 4.1187e-08 0 4.1301e-08 0 4.1304e-08 0.0021 4.1307e-08 0 4.1421e-08 0 4.1424e-08 0.0021 4.1427e-08 0 4.1541e-08 0 4.1544e-08 0.0021 4.1547e-08 0 4.1661e-08 0 4.1664e-08 0.0021 4.1667e-08 0 4.1781e-08 0 4.1784e-08 0.0021 4.1787e-08 0 4.1901e-08 0 4.1904e-08 0.0021 4.1907e-08 0 4.2021e-08 0 4.2024e-08 0.0021 4.2027e-08 0 4.2141e-08 0 4.2144e-08 0.0021 4.2147e-08 0 4.2261e-08 0 4.2264e-08 0.0021 4.2267e-08 0 4.2381e-08 0 4.2384e-08 0.0021 4.2387e-08 0 4.2501e-08 0 4.2504e-08 0.0021 4.2507e-08 0 4.2621e-08 0 4.2624e-08 0.0021 4.2627e-08 0 4.2741e-08 0 4.2744e-08 0.0021 4.2747e-08 0 4.2861e-08 0 4.2864e-08 0.0021 4.2867e-08 0 4.2981e-08 0 4.2984e-08 0.0021 4.2987e-08 0 4.3101e-08 0 4.3104e-08 0.0021 4.3107e-08 0 4.3221e-08 0 4.3224e-08 0.0021 4.3227e-08 0 4.3341e-08 0 4.3344e-08 0.0021 4.3347e-08 0 4.3461e-08 0 4.3464e-08 0.0021 4.3467e-08 0 4.3581e-08 0 4.3584e-08 0.0021 4.3587e-08 0 4.3701e-08 0 4.3704e-08 0.0021 4.3707e-08 0 4.3821e-08 0 4.3824e-08 0.0021 4.3827e-08 0 4.3941e-08 0 4.3944e-08 0.0021 4.3947e-08 0 4.4061e-08 0 4.4064e-08 0.0021 4.4067e-08 0 4.4181e-08 0 4.4184e-08 0.0021 4.4187e-08 0 4.4301e-08 0 4.4304e-08 0.0021 4.4307e-08 0 4.4421e-08 0 4.4424e-08 0.0021 4.4427e-08 0 4.4541e-08 0 4.4544e-08 0.0021 4.4547e-08 0 4.4661e-08 0 4.4664e-08 0.0021 4.4667e-08 0 4.4781e-08 0 4.4784e-08 0.0021 4.4787e-08 0 4.4901e-08 0 4.4904e-08 0.0021 4.4907e-08 0 4.5021e-08 0 4.5024e-08 0.0021 4.5027e-08 0 4.5141e-08 0 4.5144e-08 0.0021 4.5147e-08 0 4.5261e-08 0 4.5264e-08 0.0021 4.5267e-08 0 4.5381e-08 0 4.5384e-08 0.0021 4.5387e-08 0 4.5501e-08 0 4.5504e-08 0.0021 4.5507e-08 0 4.5621e-08 0 4.5624e-08 0.0021 4.5627e-08 0 4.5741e-08 0 4.5744e-08 0.0021 4.5747e-08 0 4.5861e-08 0 4.5864e-08 0.0021 4.5867e-08 0 4.5981e-08 0 4.5984e-08 0.0021 4.5987e-08 0 4.6101e-08 0 4.6104e-08 0.0021 4.6107e-08 0 4.6221e-08 0 4.6224e-08 0.0021 4.6227e-08 0 4.6341e-08 0 4.6344e-08 0.0021 4.6347e-08 0 4.6461e-08 0 4.6464e-08 0.0021 4.6467e-08 0 4.6581e-08 0 4.6584e-08 0.0021 4.6587e-08 0 4.6701e-08 0 4.6704e-08 0.0021 4.6707e-08 0 4.6821e-08 0 4.6824e-08 0.0021 4.6827e-08 0 4.6941e-08 0 4.6944e-08 0.0021 4.6947e-08 0 4.7061e-08 0 4.7064e-08 0.0021 4.7067e-08 0 4.7181e-08 0 4.7184e-08 0.0021 4.7187e-08 0 4.7301e-08 0 4.7304e-08 0.0021 4.7307e-08 0 4.7421e-08 0 4.7424e-08 0.0021 4.7427e-08 0 4.7541e-08 0 4.7544e-08 0.0021 4.7547e-08 0 4.7661e-08 0 4.7664e-08 0.0021 4.7667e-08 0 4.7781e-08 0 4.7784e-08 0.0021 4.7787e-08 0)
IT03|T 0 T03  PWL(0 0 2.1e-11 0 2.4e-11 0.0021 2.7e-11 0 1.41e-10 0 1.44e-10 0.0021 1.47e-10 0 2.61e-10 0 2.64e-10 0.0021 2.67e-10 0 3.81e-10 0 3.84e-10 0.0021 3.87e-10 0 5.01e-10 0 5.04e-10 0.0021 5.07e-10 0 6.21e-10 0 6.24e-10 0.0021 6.27e-10 0 7.41e-10 0 7.44e-10 0.0021 7.47e-10 0 8.61e-10 0 8.64e-10 0.0021 8.67e-10 0 9.81e-10 0 9.84e-10 0.0021 9.87e-10 0 1.101e-09 0 1.104e-09 0.0021 1.107e-09 0 1.221e-09 0 1.224e-09 0.0021 1.227e-09 0 1.341e-09 0 1.344e-09 0.0021 1.347e-09 0 1.461e-09 0 1.464e-09 0.0021 1.467e-09 0 1.581e-09 0 1.584e-09 0.0021 1.587e-09 0 1.701e-09 0 1.704e-09 0.0021 1.707e-09 0 1.821e-09 0 1.824e-09 0.0021 1.827e-09 0 1.941e-09 0 1.944e-09 0.0021 1.947e-09 0 2.061e-09 0 2.064e-09 0.0021 2.067e-09 0 2.181e-09 0 2.184e-09 0.0021 2.187e-09 0 2.301e-09 0 2.304e-09 0.0021 2.307e-09 0 2.421e-09 0 2.424e-09 0.0021 2.427e-09 0 2.541e-09 0 2.544e-09 0.0021 2.547e-09 0 2.661e-09 0 2.664e-09 0.0021 2.667e-09 0 2.781e-09 0 2.784e-09 0.0021 2.787e-09 0 2.901e-09 0 2.904e-09 0.0021 2.907e-09 0 3.021e-09 0 3.024e-09 0.0021 3.027e-09 0 3.141e-09 0 3.144e-09 0.0021 3.147e-09 0 3.261e-09 0 3.264e-09 0.0021 3.267e-09 0 3.381e-09 0 3.384e-09 0.0021 3.387e-09 0 3.501e-09 0 3.504e-09 0.0021 3.507e-09 0 3.621e-09 0 3.624e-09 0.0021 3.627e-09 0 3.741e-09 0 3.744e-09 0.0021 3.747e-09 0 3.861e-09 0 3.864e-09 0.0021 3.867e-09 0 3.981e-09 0 3.984e-09 0.0021 3.987e-09 0 4.101e-09 0 4.104e-09 0.0021 4.107e-09 0 4.221e-09 0 4.224e-09 0.0021 4.227e-09 0 4.341e-09 0 4.344e-09 0.0021 4.347e-09 0 4.461e-09 0 4.464e-09 0.0021 4.467e-09 0 4.581e-09 0 4.584e-09 0.0021 4.587e-09 0 4.701e-09 0 4.704e-09 0.0021 4.707e-09 0 4.821e-09 0 4.824e-09 0.0021 4.827e-09 0 4.941e-09 0 4.944e-09 0.0021 4.947e-09 0 5.061e-09 0 5.064e-09 0.0021 5.067e-09 0 5.181e-09 0 5.184e-09 0.0021 5.187e-09 0 5.301e-09 0 5.304e-09 0.0021 5.307e-09 0 5.421e-09 0 5.424e-09 0.0021 5.427e-09 0 5.541e-09 0 5.544e-09 0.0021 5.547e-09 0 5.661e-09 0 5.664e-09 0.0021 5.667e-09 0 5.781e-09 0 5.784e-09 0.0021 5.787e-09 0 5.901e-09 0 5.904e-09 0.0021 5.907e-09 0 6.021e-09 0 6.024e-09 0.0021 6.027e-09 0 6.141e-09 0 6.144e-09 0.0021 6.147e-09 0 6.261e-09 0 6.264e-09 0.0021 6.267e-09 0 6.381e-09 0 6.384e-09 0.0021 6.387e-09 0 6.501e-09 0 6.504e-09 0.0021 6.507e-09 0 6.621e-09 0 6.624e-09 0.0021 6.627e-09 0 6.741e-09 0 6.744e-09 0.0021 6.747e-09 0 6.861e-09 0 6.864e-09 0.0021 6.867e-09 0 6.981e-09 0 6.984e-09 0.0021 6.987e-09 0 7.101e-09 0 7.104e-09 0.0021 7.107e-09 0 7.221e-09 0 7.224e-09 0.0021 7.227e-09 0 7.341e-09 0 7.344e-09 0.0021 7.347e-09 0 7.461e-09 0 7.464e-09 0.0021 7.467e-09 0 7.581e-09 0 7.584e-09 0.0021 7.587e-09 0 7.701e-09 0 7.704e-09 0.0021 7.707e-09 0 7.821e-09 0 7.824e-09 0.0021 7.827e-09 0 7.941e-09 0 7.944e-09 0.0021 7.947e-09 0 8.061e-09 0 8.064e-09 0.0021 8.067e-09 0 8.181e-09 0 8.184e-09 0.0021 8.187e-09 0 8.301e-09 0 8.304e-09 0.0021 8.307e-09 0 8.421e-09 0 8.424e-09 0.0021 8.427e-09 0 8.541e-09 0 8.544e-09 0.0021 8.547e-09 0 8.661e-09 0 8.664e-09 0.0021 8.667e-09 0 8.781e-09 0 8.784e-09 0.0021 8.787e-09 0 8.901e-09 0 8.904e-09 0.0021 8.907e-09 0 9.021e-09 0 9.024e-09 0.0021 9.027e-09 0 9.141e-09 0 9.144e-09 0.0021 9.147e-09 0 9.261e-09 0 9.264e-09 0.0021 9.267e-09 0 9.381e-09 0 9.384e-09 0.0021 9.387e-09 0 9.501e-09 0 9.504e-09 0.0021 9.507e-09 0 9.621e-09 0 9.624e-09 0.0021 9.627e-09 0 9.741e-09 0 9.744e-09 0.0021 9.747e-09 0 9.861e-09 0 9.864e-09 0.0021 9.867e-09 0 9.981e-09 0 9.984e-09 0.0021 9.987e-09 0 1.0101e-08 0 1.0104e-08 0.0021 1.0107e-08 0 1.0221e-08 0 1.0224e-08 0.0021 1.0227e-08 0 1.0341e-08 0 1.0344e-08 0.0021 1.0347e-08 0 1.0461e-08 0 1.0464e-08 0.0021 1.0467e-08 0 1.0581e-08 0 1.0584e-08 0.0021 1.0587e-08 0 1.0701e-08 0 1.0704e-08 0.0021 1.0707e-08 0 1.0821e-08 0 1.0824e-08 0.0021 1.0827e-08 0 1.0941e-08 0 1.0944e-08 0.0021 1.0947e-08 0 1.1061e-08 0 1.1064e-08 0.0021 1.1067e-08 0 1.1181e-08 0 1.1184e-08 0.0021 1.1187e-08 0 1.1301e-08 0 1.1304e-08 0.0021 1.1307e-08 0 1.1421e-08 0 1.1424e-08 0.0021 1.1427e-08 0 1.1541e-08 0 1.1544e-08 0.0021 1.1547e-08 0 1.1661e-08 0 1.1664e-08 0.0021 1.1667e-08 0 1.1781e-08 0 1.1784e-08 0.0021 1.1787e-08 0 1.1901e-08 0 1.1904e-08 0.0021 1.1907e-08 0 1.2021e-08 0 1.2024e-08 0.0021 1.2027e-08 0 1.2141e-08 0 1.2144e-08 0.0021 1.2147e-08 0 1.2261e-08 0 1.2264e-08 0.0021 1.2267e-08 0 1.2381e-08 0 1.2384e-08 0.0021 1.2387e-08 0 1.2501e-08 0 1.2504e-08 0.0021 1.2507e-08 0 1.2621e-08 0 1.2624e-08 0.0021 1.2627e-08 0 1.2741e-08 0 1.2744e-08 0.0021 1.2747e-08 0 1.2861e-08 0 1.2864e-08 0.0021 1.2867e-08 0 1.2981e-08 0 1.2984e-08 0.0021 1.2987e-08 0 1.3101e-08 0 1.3104e-08 0.0021 1.3107e-08 0 1.3221e-08 0 1.3224e-08 0.0021 1.3227e-08 0 1.3341e-08 0 1.3344e-08 0.0021 1.3347e-08 0 1.3461e-08 0 1.3464e-08 0.0021 1.3467e-08 0 1.3581e-08 0 1.3584e-08 0.0021 1.3587e-08 0 1.3701e-08 0 1.3704e-08 0.0021 1.3707e-08 0 1.3821e-08 0 1.3824e-08 0.0021 1.3827e-08 0 1.3941e-08 0 1.3944e-08 0.0021 1.3947e-08 0 1.4061e-08 0 1.4064e-08 0.0021 1.4067e-08 0 1.4181e-08 0 1.4184e-08 0.0021 1.4187e-08 0 1.4301e-08 0 1.4304e-08 0.0021 1.4307e-08 0 1.4421e-08 0 1.4424e-08 0.0021 1.4427e-08 0 1.4541e-08 0 1.4544e-08 0.0021 1.4547e-08 0 1.4661e-08 0 1.4664e-08 0.0021 1.4667e-08 0 1.4781e-08 0 1.4784e-08 0.0021 1.4787e-08 0 1.4901e-08 0 1.4904e-08 0.0021 1.4907e-08 0 1.5021e-08 0 1.5024e-08 0.0021 1.5027e-08 0 1.5141e-08 0 1.5144e-08 0.0021 1.5147e-08 0 1.5261e-08 0 1.5264e-08 0.0021 1.5267e-08 0 1.5381e-08 0 1.5384e-08 0.0021 1.5387e-08 0 1.5501e-08 0 1.5504e-08 0.0021 1.5507e-08 0 1.5621e-08 0 1.5624e-08 0.0021 1.5627e-08 0 1.5741e-08 0 1.5744e-08 0.0021 1.5747e-08 0 1.5861e-08 0 1.5864e-08 0.0021 1.5867e-08 0 1.5981e-08 0 1.5984e-08 0.0021 1.5987e-08 0 1.6101e-08 0 1.6104e-08 0.0021 1.6107e-08 0 1.6221e-08 0 1.6224e-08 0.0021 1.6227e-08 0 1.6341e-08 0 1.6344e-08 0.0021 1.6347e-08 0 1.6461e-08 0 1.6464e-08 0.0021 1.6467e-08 0 1.6581e-08 0 1.6584e-08 0.0021 1.6587e-08 0 1.6701e-08 0 1.6704e-08 0.0021 1.6707e-08 0 1.6821e-08 0 1.6824e-08 0.0021 1.6827e-08 0 1.6941e-08 0 1.6944e-08 0.0021 1.6947e-08 0 1.7061e-08 0 1.7064e-08 0.0021 1.7067e-08 0 1.7181e-08 0 1.7184e-08 0.0021 1.7187e-08 0 1.7301e-08 0 1.7304e-08 0.0021 1.7307e-08 0 1.7421e-08 0 1.7424e-08 0.0021 1.7427e-08 0 1.7541e-08 0 1.7544e-08 0.0021 1.7547e-08 0 1.7661e-08 0 1.7664e-08 0.0021 1.7667e-08 0 1.7781e-08 0 1.7784e-08 0.0021 1.7787e-08 0 1.7901e-08 0 1.7904e-08 0.0021 1.7907e-08 0 1.8021e-08 0 1.8024e-08 0.0021 1.8027e-08 0 1.8141e-08 0 1.8144e-08 0.0021 1.8147e-08 0 1.8261e-08 0 1.8264e-08 0.0021 1.8267e-08 0 1.8381e-08 0 1.8384e-08 0.0021 1.8387e-08 0 1.8501e-08 0 1.8504e-08 0.0021 1.8507e-08 0 1.8621e-08 0 1.8624e-08 0.0021 1.8627e-08 0 1.8741e-08 0 1.8744e-08 0.0021 1.8747e-08 0 1.8861e-08 0 1.8864e-08 0.0021 1.8867e-08 0 1.8981e-08 0 1.8984e-08 0.0021 1.8987e-08 0 1.9101e-08 0 1.9104e-08 0.0021 1.9107e-08 0 1.9221e-08 0 1.9224e-08 0.0021 1.9227e-08 0 1.9341e-08 0 1.9344e-08 0.0021 1.9347e-08 0 1.9461e-08 0 1.9464e-08 0.0021 1.9467e-08 0 1.9581e-08 0 1.9584e-08 0.0021 1.9587e-08 0 1.9701e-08 0 1.9704e-08 0.0021 1.9707e-08 0 1.9821e-08 0 1.9824e-08 0.0021 1.9827e-08 0 1.9941e-08 0 1.9944e-08 0.0021 1.9947e-08 0 2.0061e-08 0 2.0064e-08 0.0021 2.0067e-08 0 2.0181e-08 0 2.0184e-08 0.0021 2.0187e-08 0 2.0301e-08 0 2.0304e-08 0.0021 2.0307e-08 0 2.0421e-08 0 2.0424e-08 0.0021 2.0427e-08 0 2.0541e-08 0 2.0544e-08 0.0021 2.0547e-08 0 2.0661e-08 0 2.0664e-08 0.0021 2.0667e-08 0 2.0781e-08 0 2.0784e-08 0.0021 2.0787e-08 0 2.0901e-08 0 2.0904e-08 0.0021 2.0907e-08 0 2.1021e-08 0 2.1024e-08 0.0021 2.1027e-08 0 2.1141e-08 0 2.1144e-08 0.0021 2.1147e-08 0 2.1261e-08 0 2.1264e-08 0.0021 2.1267e-08 0 2.1381e-08 0 2.1384e-08 0.0021 2.1387e-08 0 2.1501e-08 0 2.1504e-08 0.0021 2.1507e-08 0 2.1621e-08 0 2.1624e-08 0.0021 2.1627e-08 0 2.1741e-08 0 2.1744e-08 0.0021 2.1747e-08 0 2.1861e-08 0 2.1864e-08 0.0021 2.1867e-08 0 2.1981e-08 0 2.1984e-08 0.0021 2.1987e-08 0 2.2101e-08 0 2.2104e-08 0.0021 2.2107e-08 0 2.2221e-08 0 2.2224e-08 0.0021 2.2227e-08 0 2.2341e-08 0 2.2344e-08 0.0021 2.2347e-08 0 2.2461e-08 0 2.2464e-08 0.0021 2.2467e-08 0 2.2581e-08 0 2.2584e-08 0.0021 2.2587e-08 0 2.2701e-08 0 2.2704e-08 0.0021 2.2707e-08 0 2.2821e-08 0 2.2824e-08 0.0021 2.2827e-08 0 2.2941e-08 0 2.2944e-08 0.0021 2.2947e-08 0 2.3061e-08 0 2.3064e-08 0.0021 2.3067e-08 0 2.3181e-08 0 2.3184e-08 0.0021 2.3187e-08 0 2.3301e-08 0 2.3304e-08 0.0021 2.3307e-08 0 2.3421e-08 0 2.3424e-08 0.0021 2.3427e-08 0 2.3541e-08 0 2.3544e-08 0.0021 2.3547e-08 0 2.3661e-08 0 2.3664e-08 0.0021 2.3667e-08 0 2.3781e-08 0 2.3784e-08 0.0021 2.3787e-08 0 2.3901e-08 0 2.3904e-08 0.0021 2.3907e-08 0 2.4021e-08 0 2.4024e-08 0.0021 2.4027e-08 0 2.4141e-08 0 2.4144e-08 0.0021 2.4147e-08 0 2.4261e-08 0 2.4264e-08 0.0021 2.4267e-08 0 2.4381e-08 0 2.4384e-08 0.0021 2.4387e-08 0 2.4501e-08 0 2.4504e-08 0.0021 2.4507e-08 0 2.4621e-08 0 2.4624e-08 0.0021 2.4627e-08 0 2.4741e-08 0 2.4744e-08 0.0021 2.4747e-08 0 2.4861e-08 0 2.4864e-08 0.0021 2.4867e-08 0 2.4981e-08 0 2.4984e-08 0.0021 2.4987e-08 0 2.5101e-08 0 2.5104e-08 0.0021 2.5107e-08 0 2.5221e-08 0 2.5224e-08 0.0021 2.5227e-08 0 2.5341e-08 0 2.5344e-08 0.0021 2.5347e-08 0 2.5461e-08 0 2.5464e-08 0.0021 2.5467e-08 0 2.5581e-08 0 2.5584e-08 0.0021 2.5587e-08 0 2.5701e-08 0 2.5704e-08 0.0021 2.5707e-08 0 2.5821e-08 0 2.5824e-08 0.0021 2.5827e-08 0 2.5941e-08 0 2.5944e-08 0.0021 2.5947e-08 0 2.6061e-08 0 2.6064e-08 0.0021 2.6067e-08 0 2.6181e-08 0 2.6184e-08 0.0021 2.6187e-08 0 2.6301e-08 0 2.6304e-08 0.0021 2.6307e-08 0 2.6421e-08 0 2.6424e-08 0.0021 2.6427e-08 0 2.6541e-08 0 2.6544e-08 0.0021 2.6547e-08 0 2.6661e-08 0 2.6664e-08 0.0021 2.6667e-08 0 2.6781e-08 0 2.6784e-08 0.0021 2.6787e-08 0 2.6901e-08 0 2.6904e-08 0.0021 2.6907e-08 0 2.7021e-08 0 2.7024e-08 0.0021 2.7027e-08 0 2.7141e-08 0 2.7144e-08 0.0021 2.7147e-08 0 2.7261e-08 0 2.7264e-08 0.0021 2.7267e-08 0 2.7381e-08 0 2.7384e-08 0.0021 2.7387e-08 0 2.7501e-08 0 2.7504e-08 0.0021 2.7507e-08 0 2.7621e-08 0 2.7624e-08 0.0021 2.7627e-08 0 2.7741e-08 0 2.7744e-08 0.0021 2.7747e-08 0 2.7861e-08 0 2.7864e-08 0.0021 2.7867e-08 0 2.7981e-08 0 2.7984e-08 0.0021 2.7987e-08 0 2.8101e-08 0 2.8104e-08 0.0021 2.8107e-08 0 2.8221e-08 0 2.8224e-08 0.0021 2.8227e-08 0 2.8341e-08 0 2.8344e-08 0.0021 2.8347e-08 0 2.8461e-08 0 2.8464e-08 0.0021 2.8467e-08 0 2.8581e-08 0 2.8584e-08 0.0021 2.8587e-08 0 2.8701e-08 0 2.8704e-08 0.0021 2.8707e-08 0 2.8821e-08 0 2.8824e-08 0.0021 2.8827e-08 0 2.8941e-08 0 2.8944e-08 0.0021 2.8947e-08 0 2.9061e-08 0 2.9064e-08 0.0021 2.9067e-08 0 2.9181e-08 0 2.9184e-08 0.0021 2.9187e-08 0 2.9301e-08 0 2.9304e-08 0.0021 2.9307e-08 0 2.9421e-08 0 2.9424e-08 0.0021 2.9427e-08 0 2.9541e-08 0 2.9544e-08 0.0021 2.9547e-08 0 2.9661e-08 0 2.9664e-08 0.0021 2.9667e-08 0 2.9781e-08 0 2.9784e-08 0.0021 2.9787e-08 0 2.9901e-08 0 2.9904e-08 0.0021 2.9907e-08 0 3.0021e-08 0 3.0024e-08 0.0021 3.0027e-08 0 3.0141e-08 0 3.0144e-08 0.0021 3.0147e-08 0 3.0261e-08 0 3.0264e-08 0.0021 3.0267e-08 0 3.0381e-08 0 3.0384e-08 0.0021 3.0387e-08 0 3.0501e-08 0 3.0504e-08 0.0021 3.0507e-08 0 3.0621e-08 0 3.0624e-08 0.0021 3.0627e-08 0 3.0741e-08 0 3.0744e-08 0.0021 3.0747e-08 0 3.0861e-08 0 3.0864e-08 0.0021 3.0867e-08 0 3.0981e-08 0 3.0984e-08 0.0021 3.0987e-08 0 3.1101e-08 0 3.1104e-08 0.0021 3.1107e-08 0 3.1221e-08 0 3.1224e-08 0.0021 3.1227e-08 0 3.1341e-08 0 3.1344e-08 0.0021 3.1347e-08 0 3.1461e-08 0 3.1464e-08 0.0021 3.1467e-08 0 3.1581e-08 0 3.1584e-08 0.0021 3.1587e-08 0 3.1701e-08 0 3.1704e-08 0.0021 3.1707e-08 0 3.1821e-08 0 3.1824e-08 0.0021 3.1827e-08 0 3.1941e-08 0 3.1944e-08 0.0021 3.1947e-08 0 3.2061e-08 0 3.2064e-08 0.0021 3.2067e-08 0 3.2181e-08 0 3.2184e-08 0.0021 3.2187e-08 0 3.2301e-08 0 3.2304e-08 0.0021 3.2307e-08 0 3.2421e-08 0 3.2424e-08 0.0021 3.2427e-08 0 3.2541e-08 0 3.2544e-08 0.0021 3.2547e-08 0 3.2661e-08 0 3.2664e-08 0.0021 3.2667e-08 0 3.2781e-08 0 3.2784e-08 0.0021 3.2787e-08 0 3.2901e-08 0 3.2904e-08 0.0021 3.2907e-08 0 3.3021e-08 0 3.3024e-08 0.0021 3.3027e-08 0 3.3141e-08 0 3.3144e-08 0.0021 3.3147e-08 0 3.3261e-08 0 3.3264e-08 0.0021 3.3267e-08 0 3.3381e-08 0 3.3384e-08 0.0021 3.3387e-08 0 3.3501e-08 0 3.3504e-08 0.0021 3.3507e-08 0 3.3621e-08 0 3.3624e-08 0.0021 3.3627e-08 0 3.3741e-08 0 3.3744e-08 0.0021 3.3747e-08 0 3.3861e-08 0 3.3864e-08 0.0021 3.3867e-08 0 3.3981e-08 0 3.3984e-08 0.0021 3.3987e-08 0 3.4101e-08 0 3.4104e-08 0.0021 3.4107e-08 0 3.4221e-08 0 3.4224e-08 0.0021 3.4227e-08 0 3.4341e-08 0 3.4344e-08 0.0021 3.4347e-08 0 3.4461e-08 0 3.4464e-08 0.0021 3.4467e-08 0 3.4581e-08 0 3.4584e-08 0.0021 3.4587e-08 0 3.4701e-08 0 3.4704e-08 0.0021 3.4707e-08 0 3.4821e-08 0 3.4824e-08 0.0021 3.4827e-08 0 3.4941e-08 0 3.4944e-08 0.0021 3.4947e-08 0 3.5061e-08 0 3.5064e-08 0.0021 3.5067e-08 0 3.5181e-08 0 3.5184e-08 0.0021 3.5187e-08 0 3.5301e-08 0 3.5304e-08 0.0021 3.5307e-08 0 3.5421e-08 0 3.5424e-08 0.0021 3.5427e-08 0 3.5541e-08 0 3.5544e-08 0.0021 3.5547e-08 0 3.5661e-08 0 3.5664e-08 0.0021 3.5667e-08 0 3.5781e-08 0 3.5784e-08 0.0021 3.5787e-08 0 3.5901e-08 0 3.5904e-08 0.0021 3.5907e-08 0 3.6021e-08 0 3.6024e-08 0.0021 3.6027e-08 0 3.6141e-08 0 3.6144e-08 0.0021 3.6147e-08 0 3.6261e-08 0 3.6264e-08 0.0021 3.6267e-08 0 3.6381e-08 0 3.6384e-08 0.0021 3.6387e-08 0 3.6501e-08 0 3.6504e-08 0.0021 3.6507e-08 0 3.6621e-08 0 3.6624e-08 0.0021 3.6627e-08 0 3.6741e-08 0 3.6744e-08 0.0021 3.6747e-08 0 3.6861e-08 0 3.6864e-08 0.0021 3.6867e-08 0 3.6981e-08 0 3.6984e-08 0.0021 3.6987e-08 0 3.7101e-08 0 3.7104e-08 0.0021 3.7107e-08 0 3.7221e-08 0 3.7224e-08 0.0021 3.7227e-08 0 3.7341e-08 0 3.7344e-08 0.0021 3.7347e-08 0 3.7461e-08 0 3.7464e-08 0.0021 3.7467e-08 0 3.7581e-08 0 3.7584e-08 0.0021 3.7587e-08 0 3.7701e-08 0 3.7704e-08 0.0021 3.7707e-08 0 3.7821e-08 0 3.7824e-08 0.0021 3.7827e-08 0 3.7941e-08 0 3.7944e-08 0.0021 3.7947e-08 0 3.8061e-08 0 3.8064e-08 0.0021 3.8067e-08 0 3.8181e-08 0 3.8184e-08 0.0021 3.8187e-08 0 3.8301e-08 0 3.8304e-08 0.0021 3.8307e-08 0 3.8421e-08 0 3.8424e-08 0.0021 3.8427e-08 0 3.8541e-08 0 3.8544e-08 0.0021 3.8547e-08 0 3.8661e-08 0 3.8664e-08 0.0021 3.8667e-08 0 3.8781e-08 0 3.8784e-08 0.0021 3.8787e-08 0 3.8901e-08 0 3.8904e-08 0.0021 3.8907e-08 0 3.9021e-08 0 3.9024e-08 0.0021 3.9027e-08 0 3.9141e-08 0 3.9144e-08 0.0021 3.9147e-08 0 3.9261e-08 0 3.9264e-08 0.0021 3.9267e-08 0 3.9381e-08 0 3.9384e-08 0.0021 3.9387e-08 0 3.9501e-08 0 3.9504e-08 0.0021 3.9507e-08 0 3.9621e-08 0 3.9624e-08 0.0021 3.9627e-08 0 3.9741e-08 0 3.9744e-08 0.0021 3.9747e-08 0 3.9861e-08 0 3.9864e-08 0.0021 3.9867e-08 0 3.9981e-08 0 3.9984e-08 0.0021 3.9987e-08 0 4.0101e-08 0 4.0104e-08 0.0021 4.0107e-08 0 4.0221e-08 0 4.0224e-08 0.0021 4.0227e-08 0 4.0341e-08 0 4.0344e-08 0.0021 4.0347e-08 0 4.0461e-08 0 4.0464e-08 0.0021 4.0467e-08 0 4.0581e-08 0 4.0584e-08 0.0021 4.0587e-08 0 4.0701e-08 0 4.0704e-08 0.0021 4.0707e-08 0 4.0821e-08 0 4.0824e-08 0.0021 4.0827e-08 0 4.0941e-08 0 4.0944e-08 0.0021 4.0947e-08 0 4.1061e-08 0 4.1064e-08 0.0021 4.1067e-08 0 4.1181e-08 0 4.1184e-08 0.0021 4.1187e-08 0 4.1301e-08 0 4.1304e-08 0.0021 4.1307e-08 0 4.1421e-08 0 4.1424e-08 0.0021 4.1427e-08 0 4.1541e-08 0 4.1544e-08 0.0021 4.1547e-08 0 4.1661e-08 0 4.1664e-08 0.0021 4.1667e-08 0 4.1781e-08 0 4.1784e-08 0.0021 4.1787e-08 0 4.1901e-08 0 4.1904e-08 0.0021 4.1907e-08 0 4.2021e-08 0 4.2024e-08 0.0021 4.2027e-08 0 4.2141e-08 0 4.2144e-08 0.0021 4.2147e-08 0 4.2261e-08 0 4.2264e-08 0.0021 4.2267e-08 0 4.2381e-08 0 4.2384e-08 0.0021 4.2387e-08 0 4.2501e-08 0 4.2504e-08 0.0021 4.2507e-08 0 4.2621e-08 0 4.2624e-08 0.0021 4.2627e-08 0 4.2741e-08 0 4.2744e-08 0.0021 4.2747e-08 0 4.2861e-08 0 4.2864e-08 0.0021 4.2867e-08 0 4.2981e-08 0 4.2984e-08 0.0021 4.2987e-08 0 4.3101e-08 0 4.3104e-08 0.0021 4.3107e-08 0 4.3221e-08 0 4.3224e-08 0.0021 4.3227e-08 0 4.3341e-08 0 4.3344e-08 0.0021 4.3347e-08 0 4.3461e-08 0 4.3464e-08 0.0021 4.3467e-08 0 4.3581e-08 0 4.3584e-08 0.0021 4.3587e-08 0 4.3701e-08 0 4.3704e-08 0.0021 4.3707e-08 0 4.3821e-08 0 4.3824e-08 0.0021 4.3827e-08 0 4.3941e-08 0 4.3944e-08 0.0021 4.3947e-08 0 4.4061e-08 0 4.4064e-08 0.0021 4.4067e-08 0 4.4181e-08 0 4.4184e-08 0.0021 4.4187e-08 0 4.4301e-08 0 4.4304e-08 0.0021 4.4307e-08 0 4.4421e-08 0 4.4424e-08 0.0021 4.4427e-08 0 4.4541e-08 0 4.4544e-08 0.0021 4.4547e-08 0 4.4661e-08 0 4.4664e-08 0.0021 4.4667e-08 0 4.4781e-08 0 4.4784e-08 0.0021 4.4787e-08 0 4.4901e-08 0 4.4904e-08 0.0021 4.4907e-08 0 4.5021e-08 0 4.5024e-08 0.0021 4.5027e-08 0 4.5141e-08 0 4.5144e-08 0.0021 4.5147e-08 0 4.5261e-08 0 4.5264e-08 0.0021 4.5267e-08 0 4.5381e-08 0 4.5384e-08 0.0021 4.5387e-08 0 4.5501e-08 0 4.5504e-08 0.0021 4.5507e-08 0 4.5621e-08 0 4.5624e-08 0.0021 4.5627e-08 0 4.5741e-08 0 4.5744e-08 0.0021 4.5747e-08 0 4.5861e-08 0 4.5864e-08 0.0021 4.5867e-08 0 4.5981e-08 0 4.5984e-08 0.0021 4.5987e-08 0 4.6101e-08 0 4.6104e-08 0.0021 4.6107e-08 0 4.6221e-08 0 4.6224e-08 0.0021 4.6227e-08 0 4.6341e-08 0 4.6344e-08 0.0021 4.6347e-08 0 4.6461e-08 0 4.6464e-08 0.0021 4.6467e-08 0 4.6581e-08 0 4.6584e-08 0.0021 4.6587e-08 0 4.6701e-08 0 4.6704e-08 0.0021 4.6707e-08 0 4.6821e-08 0 4.6824e-08 0.0021 4.6827e-08 0 4.6941e-08 0 4.6944e-08 0.0021 4.6947e-08 0 4.7061e-08 0 4.7064e-08 0.0021 4.7067e-08 0 4.7181e-08 0 4.7184e-08 0.0021 4.7187e-08 0 4.7301e-08 0 4.7304e-08 0.0021 4.7307e-08 0 4.7421e-08 0 4.7424e-08 0.0021 4.7427e-08 0 4.7541e-08 0 4.7544e-08 0.0021 4.7547e-08 0 4.7661e-08 0 4.7664e-08 0.0021 4.7667e-08 0 4.7781e-08 0 4.7784e-08 0.0021 4.7787e-08 0)
LSPL_IG0_0|1 IG0_0_RX SPL_IG0_0|D1  2e-12
LSPL_IG0_0|2 SPL_IG0_0|D1 SPL_IG0_0|D2  4.135667696e-12
LSPL_IG0_0|3 SPL_IG0_0|D2 SPL_IG0_0|JCT  9.84682784761905e-13
LSPL_IG0_0|4 SPL_IG0_0|JCT SPL_IG0_0|QA1  9.84682784761905e-13
LSPL_IG0_0|5 SPL_IG0_0|QA1 IG0_0_TO0  2e-12
LSPL_IG0_0|6 SPL_IG0_0|JCT SPL_IG0_0|QB1  9.84682784761905e-13
LSPL_IG0_0|7 SPL_IG0_0|QB1 IG0_0_TO1  2e-12
LSPL_IP1_0|1 IP1_0_RX SPL_IP1_0|D1  2e-12
LSPL_IP1_0|2 SPL_IP1_0|D1 SPL_IP1_0|D2  4.135667696e-12
LSPL_IP1_0|3 SPL_IP1_0|D2 SPL_IP1_0|JCT  9.84682784761905e-13
LSPL_IP1_0|4 SPL_IP1_0|JCT SPL_IP1_0|QA1  9.84682784761905e-13
LSPL_IP1_0|5 SPL_IP1_0|QA1 IP1_0_TO1  2e-12
LSPL_IP1_0|6 SPL_IP1_0|JCT SPL_IP1_0|QB1  9.84682784761905e-13
LSPL_IP1_0|7 SPL_IP1_0|QB1 IP1_0_OUT  2e-12
LSPL_IG2_0|1 IG2_0_RX SPL_IG2_0|D1  2e-12
LSPL_IG2_0|2 SPL_IG2_0|D1 SPL_IG2_0|D2  4.135667696e-12
LSPL_IG2_0|3 SPL_IG2_0|D2 SPL_IG2_0|JCT  9.84682784761905e-13
LSPL_IG2_0|4 SPL_IG2_0|JCT SPL_IG2_0|QA1  9.84682784761905e-13
LSPL_IG2_0|5 SPL_IG2_0|QA1 IG2_0_TO2  2e-12
LSPL_IG2_0|6 SPL_IG2_0|JCT SPL_IG2_0|QB1  9.84682784761905e-13
LSPL_IG2_0|7 SPL_IG2_0|QB1 IG2_0_TO3  2e-12
LSPL_IP3_0|1 IP3_0_RX SPL_IP3_0|D1  2e-12
LSPL_IP3_0|2 SPL_IP3_0|D1 SPL_IP3_0|D2  4.135667696e-12
LSPL_IP3_0|3 SPL_IP3_0|D2 SPL_IP3_0|JCT  9.84682784761905e-13
LSPL_IP3_0|4 SPL_IP3_0|JCT SPL_IP3_0|QA1  9.84682784761905e-13
LSPL_IP3_0|5 SPL_IP3_0|QA1 IP3_0_TO1  2e-12
LSPL_IP3_0|6 SPL_IP3_0|JCT SPL_IP3_0|QB1  9.84682784761905e-13
LSPL_IP3_0|7 SPL_IP3_0|QB1 IP3_0_OUT  2e-12
IT04|T 0 T04  PWL(0 0 1.5e-11 0 1.8e-11 0.0014 2.1e-11 0 1.35e-10 0 1.38e-10 0.0014 1.41e-10 0 2.55e-10 0 2.58e-10 0.0014 2.61e-10 0 3.75e-10 0 3.78e-10 0.0014 3.81e-10 0 4.95e-10 0 4.98e-10 0.0014 5.01e-10 0 6.15e-10 0 6.18e-10 0.0014 6.21e-10 0 7.35e-10 0 7.38e-10 0.0014 7.41e-10 0 8.55e-10 0 8.58e-10 0.0014 8.61e-10 0 9.75e-10 0 9.78e-10 0.0014 9.81e-10 0 1.095e-09 0 1.098e-09 0.0014 1.101e-09 0 1.215e-09 0 1.218e-09 0.0014 1.221e-09 0 1.335e-09 0 1.338e-09 0.0014 1.341e-09 0 1.455e-09 0 1.458e-09 0.0014 1.461e-09 0 1.575e-09 0 1.578e-09 0.0014 1.581e-09 0 1.695e-09 0 1.698e-09 0.0014 1.701e-09 0 1.815e-09 0 1.818e-09 0.0014 1.821e-09 0 1.935e-09 0 1.938e-09 0.0014 1.941e-09 0 2.055e-09 0 2.058e-09 0.0014 2.061e-09 0 2.175e-09 0 2.178e-09 0.0014 2.181e-09 0 2.295e-09 0 2.298e-09 0.0014 2.301e-09 0 2.415e-09 0 2.418e-09 0.0014 2.421e-09 0 2.535e-09 0 2.538e-09 0.0014 2.541e-09 0 2.655e-09 0 2.658e-09 0.0014 2.661e-09 0 2.775e-09 0 2.778e-09 0.0014 2.781e-09 0 2.895e-09 0 2.898e-09 0.0014 2.901e-09 0 3.015e-09 0 3.018e-09 0.0014 3.021e-09 0 3.135e-09 0 3.138e-09 0.0014 3.141e-09 0 3.255e-09 0 3.258e-09 0.0014 3.261e-09 0 3.375e-09 0 3.378e-09 0.0014 3.381e-09 0 3.495e-09 0 3.498e-09 0.0014 3.501e-09 0 3.615e-09 0 3.618e-09 0.0014 3.621e-09 0 3.735e-09 0 3.738e-09 0.0014 3.741e-09 0 3.855e-09 0 3.858e-09 0.0014 3.861e-09 0 3.975e-09 0 3.978e-09 0.0014 3.981e-09 0 4.095e-09 0 4.098e-09 0.0014 4.101e-09 0 4.215e-09 0 4.218e-09 0.0014 4.221e-09 0 4.335e-09 0 4.338e-09 0.0014 4.341e-09 0 4.455e-09 0 4.458e-09 0.0014 4.461e-09 0 4.575e-09 0 4.578e-09 0.0014 4.581e-09 0 4.695e-09 0 4.698e-09 0.0014 4.701e-09 0 4.815e-09 0 4.818e-09 0.0014 4.821e-09 0 4.935e-09 0 4.938e-09 0.0014 4.941e-09 0 5.055e-09 0 5.058e-09 0.0014 5.061e-09 0 5.175e-09 0 5.178e-09 0.0014 5.181e-09 0 5.295e-09 0 5.298e-09 0.0014 5.301e-09 0 5.415e-09 0 5.418e-09 0.0014 5.421e-09 0 5.535e-09 0 5.538e-09 0.0014 5.541e-09 0 5.655e-09 0 5.658e-09 0.0014 5.661e-09 0 5.775e-09 0 5.778e-09 0.0014 5.781e-09 0 5.895e-09 0 5.898e-09 0.0014 5.901e-09 0 6.015e-09 0 6.018e-09 0.0014 6.021e-09 0 6.135e-09 0 6.138e-09 0.0014 6.141e-09 0 6.255e-09 0 6.258e-09 0.0014 6.261e-09 0 6.375e-09 0 6.378e-09 0.0014 6.381e-09 0 6.495e-09 0 6.498e-09 0.0014 6.501e-09 0 6.615e-09 0 6.618e-09 0.0014 6.621e-09 0 6.735e-09 0 6.738e-09 0.0014 6.741e-09 0 6.855e-09 0 6.858e-09 0.0014 6.861e-09 0 6.975e-09 0 6.978e-09 0.0014 6.981e-09 0 7.095e-09 0 7.098e-09 0.0014 7.101e-09 0 7.215e-09 0 7.218e-09 0.0014 7.221e-09 0 7.335e-09 0 7.338e-09 0.0014 7.341e-09 0 7.455e-09 0 7.458e-09 0.0014 7.461e-09 0 7.575e-09 0 7.578e-09 0.0014 7.581e-09 0 7.695e-09 0 7.698e-09 0.0014 7.701e-09 0 7.815e-09 0 7.818e-09 0.0014 7.821e-09 0 7.935e-09 0 7.938e-09 0.0014 7.941e-09 0 8.055e-09 0 8.058e-09 0.0014 8.061e-09 0 8.175e-09 0 8.178e-09 0.0014 8.181e-09 0 8.295e-09 0 8.298e-09 0.0014 8.301e-09 0 8.415e-09 0 8.418e-09 0.0014 8.421e-09 0 8.535e-09 0 8.538e-09 0.0014 8.541e-09 0 8.655e-09 0 8.658e-09 0.0014 8.661e-09 0 8.775e-09 0 8.778e-09 0.0014 8.781e-09 0 8.895e-09 0 8.898e-09 0.0014 8.901e-09 0 9.015e-09 0 9.018e-09 0.0014 9.021e-09 0 9.135e-09 0 9.138e-09 0.0014 9.141e-09 0 9.255e-09 0 9.258e-09 0.0014 9.261e-09 0 9.375e-09 0 9.378e-09 0.0014 9.381e-09 0 9.495e-09 0 9.498e-09 0.0014 9.501e-09 0 9.615e-09 0 9.618e-09 0.0014 9.621e-09 0 9.735e-09 0 9.738e-09 0.0014 9.741e-09 0 9.855e-09 0 9.858e-09 0.0014 9.861e-09 0 9.975e-09 0 9.978e-09 0.0014 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0014 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0014 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0014 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0014 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0014 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0014 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0014 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0014 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0014 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0014 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0014 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0014 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0014 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0014 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0014 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0014 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0014 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0014 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0014 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0014 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0014 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0014 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0014 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0014 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0014 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0014 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0014 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0014 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0014 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0014 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0014 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0014 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0014 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0014 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0014 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0014 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0014 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0014 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0014 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0014 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0014 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0014 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0014 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0014 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0014 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0014 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0014 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0014 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0014 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0014 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0014 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0014 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0014 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0014 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0014 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0014 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0014 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0014 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0014 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0014 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0014 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0014 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0014 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0014 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0014 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0014 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0014 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0014 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0014 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0014 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0014 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0014 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0014 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0014 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0014 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0014 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0014 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0014 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0014 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0014 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0014 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0014 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0014 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0014 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0014 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0014 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0014 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0014 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0014 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0014 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0014 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0014 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0014 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0014 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0014 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0014 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0014 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0014 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0014 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0014 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0014 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0014 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0014 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0014 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0014 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0014 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0014 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0014 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0014 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0014 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0014 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0014 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0014 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0014 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0014 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0014 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0014 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0014 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0014 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0014 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0014 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0014 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0014 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0014 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0014 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0014 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0014 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0014 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0014 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0014 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0014 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0014 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0014 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0014 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0014 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0014 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0014 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0014 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0014 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0014 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0014 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0014 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0014 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0014 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0014 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0014 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0014 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0014 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0014 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0014 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0014 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0014 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0014 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0014 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0014 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0014 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0014 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0014 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0014 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0014 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0014 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0014 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0014 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0014 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0014 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0014 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0014 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0014 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0014 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0014 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0014 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0014 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0014 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0014 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0014 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0014 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0014 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0014 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0014 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0014 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0014 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0014 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0014 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0014 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0014 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0014 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0014 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0014 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0014 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0014 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0014 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0014 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0014 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0014 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0014 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0014 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0014 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0014 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0014 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0014 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0014 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0014 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0014 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0014 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0014 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0014 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0014 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0014 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0014 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0014 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0014 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0014 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0014 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0014 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0014 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0014 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0014 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0014 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0014 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0014 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0014 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0014 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0014 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0014 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0014 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0014 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0014 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0014 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0014 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0014 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0014 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0014 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0014 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0014 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0014 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0014 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0014 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0014 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0014 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0014 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0014 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0014 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0014 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0014 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0014 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0014 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0014 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0014 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0014 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0014 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0014 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0014 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0014 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0014 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0014 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0014 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0014 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0014 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0014 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0014 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0014 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0014 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0014 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0014 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0014 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0014 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0014 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0014 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0014 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0014 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0014 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0014 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0014 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0014 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0014 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0014 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0014 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0014 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0014 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0014 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0014 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0014 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0014 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0014 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0014 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0014 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0014 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0014 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0014 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0014 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0014 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0014 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0014 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0014 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0014 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0014 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0014 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0014 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0014 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0014 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0014 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0014 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0014 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0014 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0014 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0014 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0014 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0014 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0014 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0014 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0014 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0014 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0014 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0014 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0014 4.7781e-08 0)
IT05|T 0 T05  PWL(0 0 1.5e-11 0 1.8e-11 0.0014 2.1e-11 0 1.35e-10 0 1.38e-10 0.0014 1.41e-10 0 2.55e-10 0 2.58e-10 0.0014 2.61e-10 0 3.75e-10 0 3.78e-10 0.0014 3.81e-10 0 4.95e-10 0 4.98e-10 0.0014 5.01e-10 0 6.15e-10 0 6.18e-10 0.0014 6.21e-10 0 7.35e-10 0 7.38e-10 0.0014 7.41e-10 0 8.55e-10 0 8.58e-10 0.0014 8.61e-10 0 9.75e-10 0 9.78e-10 0.0014 9.81e-10 0 1.095e-09 0 1.098e-09 0.0014 1.101e-09 0 1.215e-09 0 1.218e-09 0.0014 1.221e-09 0 1.335e-09 0 1.338e-09 0.0014 1.341e-09 0 1.455e-09 0 1.458e-09 0.0014 1.461e-09 0 1.575e-09 0 1.578e-09 0.0014 1.581e-09 0 1.695e-09 0 1.698e-09 0.0014 1.701e-09 0 1.815e-09 0 1.818e-09 0.0014 1.821e-09 0 1.935e-09 0 1.938e-09 0.0014 1.941e-09 0 2.055e-09 0 2.058e-09 0.0014 2.061e-09 0 2.175e-09 0 2.178e-09 0.0014 2.181e-09 0 2.295e-09 0 2.298e-09 0.0014 2.301e-09 0 2.415e-09 0 2.418e-09 0.0014 2.421e-09 0 2.535e-09 0 2.538e-09 0.0014 2.541e-09 0 2.655e-09 0 2.658e-09 0.0014 2.661e-09 0 2.775e-09 0 2.778e-09 0.0014 2.781e-09 0 2.895e-09 0 2.898e-09 0.0014 2.901e-09 0 3.015e-09 0 3.018e-09 0.0014 3.021e-09 0 3.135e-09 0 3.138e-09 0.0014 3.141e-09 0 3.255e-09 0 3.258e-09 0.0014 3.261e-09 0 3.375e-09 0 3.378e-09 0.0014 3.381e-09 0 3.495e-09 0 3.498e-09 0.0014 3.501e-09 0 3.615e-09 0 3.618e-09 0.0014 3.621e-09 0 3.735e-09 0 3.738e-09 0.0014 3.741e-09 0 3.855e-09 0 3.858e-09 0.0014 3.861e-09 0 3.975e-09 0 3.978e-09 0.0014 3.981e-09 0 4.095e-09 0 4.098e-09 0.0014 4.101e-09 0 4.215e-09 0 4.218e-09 0.0014 4.221e-09 0 4.335e-09 0 4.338e-09 0.0014 4.341e-09 0 4.455e-09 0 4.458e-09 0.0014 4.461e-09 0 4.575e-09 0 4.578e-09 0.0014 4.581e-09 0 4.695e-09 0 4.698e-09 0.0014 4.701e-09 0 4.815e-09 0 4.818e-09 0.0014 4.821e-09 0 4.935e-09 0 4.938e-09 0.0014 4.941e-09 0 5.055e-09 0 5.058e-09 0.0014 5.061e-09 0 5.175e-09 0 5.178e-09 0.0014 5.181e-09 0 5.295e-09 0 5.298e-09 0.0014 5.301e-09 0 5.415e-09 0 5.418e-09 0.0014 5.421e-09 0 5.535e-09 0 5.538e-09 0.0014 5.541e-09 0 5.655e-09 0 5.658e-09 0.0014 5.661e-09 0 5.775e-09 0 5.778e-09 0.0014 5.781e-09 0 5.895e-09 0 5.898e-09 0.0014 5.901e-09 0 6.015e-09 0 6.018e-09 0.0014 6.021e-09 0 6.135e-09 0 6.138e-09 0.0014 6.141e-09 0 6.255e-09 0 6.258e-09 0.0014 6.261e-09 0 6.375e-09 0 6.378e-09 0.0014 6.381e-09 0 6.495e-09 0 6.498e-09 0.0014 6.501e-09 0 6.615e-09 0 6.618e-09 0.0014 6.621e-09 0 6.735e-09 0 6.738e-09 0.0014 6.741e-09 0 6.855e-09 0 6.858e-09 0.0014 6.861e-09 0 6.975e-09 0 6.978e-09 0.0014 6.981e-09 0 7.095e-09 0 7.098e-09 0.0014 7.101e-09 0 7.215e-09 0 7.218e-09 0.0014 7.221e-09 0 7.335e-09 0 7.338e-09 0.0014 7.341e-09 0 7.455e-09 0 7.458e-09 0.0014 7.461e-09 0 7.575e-09 0 7.578e-09 0.0014 7.581e-09 0 7.695e-09 0 7.698e-09 0.0014 7.701e-09 0 7.815e-09 0 7.818e-09 0.0014 7.821e-09 0 7.935e-09 0 7.938e-09 0.0014 7.941e-09 0 8.055e-09 0 8.058e-09 0.0014 8.061e-09 0 8.175e-09 0 8.178e-09 0.0014 8.181e-09 0 8.295e-09 0 8.298e-09 0.0014 8.301e-09 0 8.415e-09 0 8.418e-09 0.0014 8.421e-09 0 8.535e-09 0 8.538e-09 0.0014 8.541e-09 0 8.655e-09 0 8.658e-09 0.0014 8.661e-09 0 8.775e-09 0 8.778e-09 0.0014 8.781e-09 0 8.895e-09 0 8.898e-09 0.0014 8.901e-09 0 9.015e-09 0 9.018e-09 0.0014 9.021e-09 0 9.135e-09 0 9.138e-09 0.0014 9.141e-09 0 9.255e-09 0 9.258e-09 0.0014 9.261e-09 0 9.375e-09 0 9.378e-09 0.0014 9.381e-09 0 9.495e-09 0 9.498e-09 0.0014 9.501e-09 0 9.615e-09 0 9.618e-09 0.0014 9.621e-09 0 9.735e-09 0 9.738e-09 0.0014 9.741e-09 0 9.855e-09 0 9.858e-09 0.0014 9.861e-09 0 9.975e-09 0 9.978e-09 0.0014 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0014 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0014 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0014 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0014 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0014 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0014 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0014 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0014 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0014 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0014 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0014 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0014 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0014 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0014 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0014 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0014 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0014 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0014 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0014 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0014 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0014 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0014 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0014 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0014 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0014 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0014 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0014 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0014 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0014 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0014 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0014 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0014 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0014 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0014 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0014 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0014 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0014 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0014 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0014 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0014 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0014 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0014 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0014 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0014 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0014 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0014 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0014 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0014 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0014 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0014 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0014 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0014 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0014 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0014 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0014 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0014 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0014 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0014 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0014 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0014 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0014 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0014 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0014 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0014 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0014 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0014 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0014 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0014 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0014 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0014 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0014 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0014 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0014 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0014 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0014 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0014 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0014 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0014 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0014 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0014 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0014 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0014 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0014 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0014 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0014 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0014 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0014 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0014 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0014 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0014 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0014 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0014 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0014 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0014 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0014 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0014 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0014 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0014 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0014 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0014 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0014 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0014 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0014 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0014 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0014 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0014 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0014 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0014 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0014 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0014 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0014 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0014 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0014 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0014 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0014 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0014 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0014 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0014 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0014 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0014 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0014 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0014 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0014 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0014 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0014 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0014 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0014 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0014 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0014 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0014 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0014 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0014 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0014 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0014 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0014 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0014 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0014 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0014 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0014 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0014 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0014 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0014 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0014 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0014 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0014 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0014 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0014 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0014 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0014 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0014 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0014 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0014 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0014 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0014 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0014 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0014 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0014 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0014 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0014 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0014 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0014 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0014 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0014 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0014 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0014 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0014 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0014 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0014 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0014 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0014 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0014 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0014 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0014 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0014 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0014 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0014 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0014 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0014 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0014 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0014 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0014 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0014 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0014 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0014 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0014 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0014 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0014 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0014 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0014 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0014 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0014 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0014 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0014 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0014 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0014 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0014 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0014 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0014 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0014 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0014 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0014 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0014 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0014 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0014 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0014 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0014 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0014 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0014 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0014 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0014 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0014 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0014 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0014 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0014 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0014 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0014 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0014 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0014 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0014 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0014 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0014 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0014 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0014 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0014 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0014 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0014 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0014 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0014 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0014 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0014 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0014 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0014 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0014 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0014 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0014 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0014 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0014 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0014 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0014 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0014 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0014 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0014 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0014 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0014 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0014 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0014 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0014 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0014 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0014 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0014 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0014 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0014 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0014 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0014 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0014 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0014 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0014 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0014 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0014 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0014 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0014 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0014 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0014 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0014 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0014 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0014 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0014 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0014 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0014 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0014 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0014 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0014 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0014 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0014 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0014 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0014 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0014 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0014 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0014 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0014 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0014 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0014 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0014 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0014 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0014 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0014 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0014 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0014 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0014 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0014 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0014 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0014 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0014 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0014 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0014 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0014 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0014 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0014 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0014 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0014 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0014 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0014 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0014 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0014 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0014 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0014 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0014 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0014 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0014 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0014 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0014 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0014 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0014 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0014 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0014 4.7781e-08 0)
IT06|T 0 T06  PWL(0 0 1.5e-11 0 1.8e-11 0.0014 2.1e-11 0 1.35e-10 0 1.38e-10 0.0014 1.41e-10 0 2.55e-10 0 2.58e-10 0.0014 2.61e-10 0 3.75e-10 0 3.78e-10 0.0014 3.81e-10 0 4.95e-10 0 4.98e-10 0.0014 5.01e-10 0 6.15e-10 0 6.18e-10 0.0014 6.21e-10 0 7.35e-10 0 7.38e-10 0.0014 7.41e-10 0 8.55e-10 0 8.58e-10 0.0014 8.61e-10 0 9.75e-10 0 9.78e-10 0.0014 9.81e-10 0 1.095e-09 0 1.098e-09 0.0014 1.101e-09 0 1.215e-09 0 1.218e-09 0.0014 1.221e-09 0 1.335e-09 0 1.338e-09 0.0014 1.341e-09 0 1.455e-09 0 1.458e-09 0.0014 1.461e-09 0 1.575e-09 0 1.578e-09 0.0014 1.581e-09 0 1.695e-09 0 1.698e-09 0.0014 1.701e-09 0 1.815e-09 0 1.818e-09 0.0014 1.821e-09 0 1.935e-09 0 1.938e-09 0.0014 1.941e-09 0 2.055e-09 0 2.058e-09 0.0014 2.061e-09 0 2.175e-09 0 2.178e-09 0.0014 2.181e-09 0 2.295e-09 0 2.298e-09 0.0014 2.301e-09 0 2.415e-09 0 2.418e-09 0.0014 2.421e-09 0 2.535e-09 0 2.538e-09 0.0014 2.541e-09 0 2.655e-09 0 2.658e-09 0.0014 2.661e-09 0 2.775e-09 0 2.778e-09 0.0014 2.781e-09 0 2.895e-09 0 2.898e-09 0.0014 2.901e-09 0 3.015e-09 0 3.018e-09 0.0014 3.021e-09 0 3.135e-09 0 3.138e-09 0.0014 3.141e-09 0 3.255e-09 0 3.258e-09 0.0014 3.261e-09 0 3.375e-09 0 3.378e-09 0.0014 3.381e-09 0 3.495e-09 0 3.498e-09 0.0014 3.501e-09 0 3.615e-09 0 3.618e-09 0.0014 3.621e-09 0 3.735e-09 0 3.738e-09 0.0014 3.741e-09 0 3.855e-09 0 3.858e-09 0.0014 3.861e-09 0 3.975e-09 0 3.978e-09 0.0014 3.981e-09 0 4.095e-09 0 4.098e-09 0.0014 4.101e-09 0 4.215e-09 0 4.218e-09 0.0014 4.221e-09 0 4.335e-09 0 4.338e-09 0.0014 4.341e-09 0 4.455e-09 0 4.458e-09 0.0014 4.461e-09 0 4.575e-09 0 4.578e-09 0.0014 4.581e-09 0 4.695e-09 0 4.698e-09 0.0014 4.701e-09 0 4.815e-09 0 4.818e-09 0.0014 4.821e-09 0 4.935e-09 0 4.938e-09 0.0014 4.941e-09 0 5.055e-09 0 5.058e-09 0.0014 5.061e-09 0 5.175e-09 0 5.178e-09 0.0014 5.181e-09 0 5.295e-09 0 5.298e-09 0.0014 5.301e-09 0 5.415e-09 0 5.418e-09 0.0014 5.421e-09 0 5.535e-09 0 5.538e-09 0.0014 5.541e-09 0 5.655e-09 0 5.658e-09 0.0014 5.661e-09 0 5.775e-09 0 5.778e-09 0.0014 5.781e-09 0 5.895e-09 0 5.898e-09 0.0014 5.901e-09 0 6.015e-09 0 6.018e-09 0.0014 6.021e-09 0 6.135e-09 0 6.138e-09 0.0014 6.141e-09 0 6.255e-09 0 6.258e-09 0.0014 6.261e-09 0 6.375e-09 0 6.378e-09 0.0014 6.381e-09 0 6.495e-09 0 6.498e-09 0.0014 6.501e-09 0 6.615e-09 0 6.618e-09 0.0014 6.621e-09 0 6.735e-09 0 6.738e-09 0.0014 6.741e-09 0 6.855e-09 0 6.858e-09 0.0014 6.861e-09 0 6.975e-09 0 6.978e-09 0.0014 6.981e-09 0 7.095e-09 0 7.098e-09 0.0014 7.101e-09 0 7.215e-09 0 7.218e-09 0.0014 7.221e-09 0 7.335e-09 0 7.338e-09 0.0014 7.341e-09 0 7.455e-09 0 7.458e-09 0.0014 7.461e-09 0 7.575e-09 0 7.578e-09 0.0014 7.581e-09 0 7.695e-09 0 7.698e-09 0.0014 7.701e-09 0 7.815e-09 0 7.818e-09 0.0014 7.821e-09 0 7.935e-09 0 7.938e-09 0.0014 7.941e-09 0 8.055e-09 0 8.058e-09 0.0014 8.061e-09 0 8.175e-09 0 8.178e-09 0.0014 8.181e-09 0 8.295e-09 0 8.298e-09 0.0014 8.301e-09 0 8.415e-09 0 8.418e-09 0.0014 8.421e-09 0 8.535e-09 0 8.538e-09 0.0014 8.541e-09 0 8.655e-09 0 8.658e-09 0.0014 8.661e-09 0 8.775e-09 0 8.778e-09 0.0014 8.781e-09 0 8.895e-09 0 8.898e-09 0.0014 8.901e-09 0 9.015e-09 0 9.018e-09 0.0014 9.021e-09 0 9.135e-09 0 9.138e-09 0.0014 9.141e-09 0 9.255e-09 0 9.258e-09 0.0014 9.261e-09 0 9.375e-09 0 9.378e-09 0.0014 9.381e-09 0 9.495e-09 0 9.498e-09 0.0014 9.501e-09 0 9.615e-09 0 9.618e-09 0.0014 9.621e-09 0 9.735e-09 0 9.738e-09 0.0014 9.741e-09 0 9.855e-09 0 9.858e-09 0.0014 9.861e-09 0 9.975e-09 0 9.978e-09 0.0014 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0014 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0014 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0014 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0014 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0014 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0014 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0014 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0014 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0014 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0014 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0014 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0014 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0014 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0014 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0014 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0014 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0014 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0014 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0014 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0014 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0014 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0014 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0014 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0014 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0014 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0014 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0014 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0014 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0014 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0014 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0014 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0014 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0014 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0014 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0014 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0014 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0014 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0014 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0014 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0014 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0014 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0014 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0014 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0014 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0014 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0014 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0014 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0014 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0014 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0014 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0014 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0014 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0014 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0014 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0014 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0014 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0014 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0014 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0014 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0014 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0014 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0014 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0014 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0014 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0014 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0014 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0014 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0014 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0014 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0014 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0014 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0014 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0014 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0014 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0014 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0014 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0014 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0014 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0014 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0014 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0014 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0014 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0014 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0014 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0014 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0014 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0014 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0014 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0014 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0014 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0014 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0014 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0014 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0014 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0014 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0014 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0014 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0014 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0014 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0014 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0014 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0014 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0014 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0014 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0014 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0014 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0014 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0014 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0014 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0014 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0014 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0014 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0014 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0014 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0014 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0014 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0014 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0014 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0014 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0014 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0014 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0014 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0014 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0014 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0014 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0014 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0014 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0014 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0014 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0014 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0014 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0014 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0014 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0014 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0014 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0014 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0014 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0014 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0014 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0014 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0014 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0014 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0014 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0014 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0014 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0014 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0014 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0014 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0014 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0014 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0014 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0014 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0014 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0014 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0014 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0014 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0014 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0014 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0014 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0014 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0014 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0014 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0014 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0014 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0014 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0014 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0014 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0014 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0014 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0014 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0014 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0014 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0014 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0014 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0014 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0014 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0014 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0014 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0014 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0014 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0014 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0014 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0014 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0014 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0014 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0014 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0014 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0014 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0014 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0014 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0014 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0014 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0014 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0014 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0014 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0014 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0014 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0014 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0014 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0014 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0014 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0014 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0014 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0014 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0014 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0014 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0014 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0014 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0014 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0014 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0014 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0014 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0014 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0014 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0014 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0014 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0014 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0014 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0014 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0014 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0014 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0014 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0014 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0014 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0014 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0014 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0014 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0014 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0014 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0014 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0014 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0014 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0014 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0014 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0014 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0014 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0014 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0014 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0014 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0014 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0014 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0014 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0014 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0014 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0014 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0014 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0014 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0014 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0014 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0014 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0014 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0014 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0014 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0014 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0014 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0014 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0014 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0014 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0014 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0014 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0014 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0014 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0014 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0014 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0014 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0014 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0014 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0014 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0014 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0014 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0014 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0014 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0014 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0014 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0014 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0014 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0014 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0014 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0014 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0014 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0014 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0014 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0014 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0014 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0014 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0014 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0014 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0014 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0014 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0014 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0014 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0014 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0014 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0014 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0014 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0014 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0014 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0014 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0014 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0014 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0014 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0014 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0014 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0014 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0014 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0014 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0014 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0014 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0014 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0014 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0014 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0014 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0014 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0014 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0014 4.7781e-08 0)
IT07|T 0 T07  PWL(0 0 1.5e-11 0 1.8e-11 0.0028 2.1e-11 0 1.35e-10 0 1.38e-10 0.0028 1.41e-10 0 2.55e-10 0 2.58e-10 0.0028 2.61e-10 0 3.75e-10 0 3.78e-10 0.0028 3.81e-10 0 4.95e-10 0 4.98e-10 0.0028 5.01e-10 0 6.15e-10 0 6.18e-10 0.0028 6.21e-10 0 7.35e-10 0 7.38e-10 0.0028 7.41e-10 0 8.55e-10 0 8.58e-10 0.0028 8.61e-10 0 9.75e-10 0 9.78e-10 0.0028 9.81e-10 0 1.095e-09 0 1.098e-09 0.0028 1.101e-09 0 1.215e-09 0 1.218e-09 0.0028 1.221e-09 0 1.335e-09 0 1.338e-09 0.0028 1.341e-09 0 1.455e-09 0 1.458e-09 0.0028 1.461e-09 0 1.575e-09 0 1.578e-09 0.0028 1.581e-09 0 1.695e-09 0 1.698e-09 0.0028 1.701e-09 0 1.815e-09 0 1.818e-09 0.0028 1.821e-09 0 1.935e-09 0 1.938e-09 0.0028 1.941e-09 0 2.055e-09 0 2.058e-09 0.0028 2.061e-09 0 2.175e-09 0 2.178e-09 0.0028 2.181e-09 0 2.295e-09 0 2.298e-09 0.0028 2.301e-09 0 2.415e-09 0 2.418e-09 0.0028 2.421e-09 0 2.535e-09 0 2.538e-09 0.0028 2.541e-09 0 2.655e-09 0 2.658e-09 0.0028 2.661e-09 0 2.775e-09 0 2.778e-09 0.0028 2.781e-09 0 2.895e-09 0 2.898e-09 0.0028 2.901e-09 0 3.015e-09 0 3.018e-09 0.0028 3.021e-09 0 3.135e-09 0 3.138e-09 0.0028 3.141e-09 0 3.255e-09 0 3.258e-09 0.0028 3.261e-09 0 3.375e-09 0 3.378e-09 0.0028 3.381e-09 0 3.495e-09 0 3.498e-09 0.0028 3.501e-09 0 3.615e-09 0 3.618e-09 0.0028 3.621e-09 0 3.735e-09 0 3.738e-09 0.0028 3.741e-09 0 3.855e-09 0 3.858e-09 0.0028 3.861e-09 0 3.975e-09 0 3.978e-09 0.0028 3.981e-09 0 4.095e-09 0 4.098e-09 0.0028 4.101e-09 0 4.215e-09 0 4.218e-09 0.0028 4.221e-09 0 4.335e-09 0 4.338e-09 0.0028 4.341e-09 0 4.455e-09 0 4.458e-09 0.0028 4.461e-09 0 4.575e-09 0 4.578e-09 0.0028 4.581e-09 0 4.695e-09 0 4.698e-09 0.0028 4.701e-09 0 4.815e-09 0 4.818e-09 0.0028 4.821e-09 0 4.935e-09 0 4.938e-09 0.0028 4.941e-09 0 5.055e-09 0 5.058e-09 0.0028 5.061e-09 0 5.175e-09 0 5.178e-09 0.0028 5.181e-09 0 5.295e-09 0 5.298e-09 0.0028 5.301e-09 0 5.415e-09 0 5.418e-09 0.0028 5.421e-09 0 5.535e-09 0 5.538e-09 0.0028 5.541e-09 0 5.655e-09 0 5.658e-09 0.0028 5.661e-09 0 5.775e-09 0 5.778e-09 0.0028 5.781e-09 0 5.895e-09 0 5.898e-09 0.0028 5.901e-09 0 6.015e-09 0 6.018e-09 0.0028 6.021e-09 0 6.135e-09 0 6.138e-09 0.0028 6.141e-09 0 6.255e-09 0 6.258e-09 0.0028 6.261e-09 0 6.375e-09 0 6.378e-09 0.0028 6.381e-09 0 6.495e-09 0 6.498e-09 0.0028 6.501e-09 0 6.615e-09 0 6.618e-09 0.0028 6.621e-09 0 6.735e-09 0 6.738e-09 0.0028 6.741e-09 0 6.855e-09 0 6.858e-09 0.0028 6.861e-09 0 6.975e-09 0 6.978e-09 0.0028 6.981e-09 0 7.095e-09 0 7.098e-09 0.0028 7.101e-09 0 7.215e-09 0 7.218e-09 0.0028 7.221e-09 0 7.335e-09 0 7.338e-09 0.0028 7.341e-09 0 7.455e-09 0 7.458e-09 0.0028 7.461e-09 0 7.575e-09 0 7.578e-09 0.0028 7.581e-09 0 7.695e-09 0 7.698e-09 0.0028 7.701e-09 0 7.815e-09 0 7.818e-09 0.0028 7.821e-09 0 7.935e-09 0 7.938e-09 0.0028 7.941e-09 0 8.055e-09 0 8.058e-09 0.0028 8.061e-09 0 8.175e-09 0 8.178e-09 0.0028 8.181e-09 0 8.295e-09 0 8.298e-09 0.0028 8.301e-09 0 8.415e-09 0 8.418e-09 0.0028 8.421e-09 0 8.535e-09 0 8.538e-09 0.0028 8.541e-09 0 8.655e-09 0 8.658e-09 0.0028 8.661e-09 0 8.775e-09 0 8.778e-09 0.0028 8.781e-09 0 8.895e-09 0 8.898e-09 0.0028 8.901e-09 0 9.015e-09 0 9.018e-09 0.0028 9.021e-09 0 9.135e-09 0 9.138e-09 0.0028 9.141e-09 0 9.255e-09 0 9.258e-09 0.0028 9.261e-09 0 9.375e-09 0 9.378e-09 0.0028 9.381e-09 0 9.495e-09 0 9.498e-09 0.0028 9.501e-09 0 9.615e-09 0 9.618e-09 0.0028 9.621e-09 0 9.735e-09 0 9.738e-09 0.0028 9.741e-09 0 9.855e-09 0 9.858e-09 0.0028 9.861e-09 0 9.975e-09 0 9.978e-09 0.0028 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0028 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0028 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0028 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0028 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0028 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0028 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0028 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0028 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0028 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0028 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0028 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0028 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0028 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0028 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0028 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0028 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0028 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0028 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0028 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0028 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0028 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0028 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0028 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0028 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0028 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0028 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0028 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0028 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0028 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0028 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0028 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0028 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0028 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0028 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0028 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0028 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0028 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0028 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0028 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0028 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0028 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0028 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0028 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0028 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0028 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0028 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0028 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0028 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0028 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0028 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0028 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0028 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0028 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0028 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0028 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0028 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0028 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0028 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0028 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0028 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0028 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0028 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0028 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0028 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0028 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0028 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0028 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0028 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0028 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0028 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0028 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0028 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0028 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0028 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0028 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0028 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0028 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0028 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0028 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0028 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0028 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0028 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0028 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0028 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0028 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0028 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0028 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0028 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0028 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0028 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0028 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0028 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0028 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0028 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0028 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0028 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0028 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0028 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0028 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0028 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0028 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0028 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0028 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0028 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0028 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0028 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0028 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0028 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0028 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0028 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0028 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0028 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0028 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0028 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0028 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0028 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0028 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0028 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0028 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0028 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0028 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0028 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0028 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0028 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0028 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0028 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0028 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0028 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0028 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0028 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0028 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0028 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0028 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0028 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0028 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0028 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0028 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0028 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0028 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0028 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0028 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0028 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0028 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0028 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0028 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0028 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0028 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0028 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0028 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0028 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0028 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0028 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0028 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0028 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0028 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0028 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0028 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0028 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0028 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0028 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0028 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0028 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0028 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0028 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0028 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0028 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0028 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0028 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0028 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0028 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0028 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0028 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0028 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0028 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0028 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0028 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0028 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0028 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0028 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0028 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0028 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0028 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0028 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0028 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0028 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0028 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0028 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0028 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0028 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0028 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0028 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0028 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0028 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0028 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0028 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0028 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0028 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0028 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0028 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0028 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0028 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0028 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0028 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0028 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0028 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0028 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0028 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0028 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0028 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0028 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0028 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0028 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0028 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0028 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0028 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0028 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0028 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0028 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0028 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0028 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0028 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0028 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0028 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0028 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0028 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0028 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0028 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0028 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0028 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0028 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0028 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0028 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0028 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0028 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0028 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0028 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0028 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0028 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0028 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0028 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0028 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0028 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0028 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0028 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0028 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0028 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0028 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0028 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0028 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0028 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0028 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0028 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0028 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0028 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0028 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0028 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0028 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0028 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0028 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0028 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0028 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0028 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0028 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0028 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0028 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0028 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0028 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0028 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0028 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0028 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0028 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0028 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0028 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0028 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0028 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0028 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0028 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0028 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0028 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0028 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0028 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0028 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0028 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0028 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0028 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0028 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0028 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0028 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0028 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0028 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0028 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0028 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0028 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0028 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0028 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0028 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0028 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0028 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0028 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0028 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0028 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0028 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0028 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0028 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0028 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0028 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0028 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0028 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0028 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0028 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0028 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0028 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0028 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0028 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0028 4.7781e-08 0)
ID01|T 0 D01  PWL(0 0 1.5e-11 0 1.8e-11 0.0007 2.1e-11 0 1.35e-10 0 1.38e-10 0.0007 1.41e-10 0 2.55e-10 0 2.58e-10 0.0007 2.61e-10 0 3.75e-10 0 3.78e-10 0.0007 3.81e-10 0 4.95e-10 0 4.98e-10 0.0007 5.01e-10 0 6.15e-10 0 6.18e-10 0.0007 6.21e-10 0 7.35e-10 0 7.38e-10 0.0007 7.41e-10 0 8.55e-10 0 8.58e-10 0.0007 8.61e-10 0 9.75e-10 0 9.78e-10 0.0007 9.81e-10 0 1.095e-09 0 1.098e-09 0.0007 1.101e-09 0 1.215e-09 0 1.218e-09 0.0007 1.221e-09 0 1.335e-09 0 1.338e-09 0.0007 1.341e-09 0 1.455e-09 0 1.458e-09 0.0007 1.461e-09 0 1.575e-09 0 1.578e-09 0.0007 1.581e-09 0 1.695e-09 0 1.698e-09 0.0007 1.701e-09 0 1.815e-09 0 1.818e-09 0.0007 1.821e-09 0 1.935e-09 0 1.938e-09 0.0007 1.941e-09 0 2.055e-09 0 2.058e-09 0.0007 2.061e-09 0 2.175e-09 0 2.178e-09 0.0007 2.181e-09 0 2.295e-09 0 2.298e-09 0.0007 2.301e-09 0 2.415e-09 0 2.418e-09 0.0007 2.421e-09 0 2.535e-09 0 2.538e-09 0.0007 2.541e-09 0 2.655e-09 0 2.658e-09 0.0007 2.661e-09 0 2.775e-09 0 2.778e-09 0.0007 2.781e-09 0 2.895e-09 0 2.898e-09 0.0007 2.901e-09 0 3.015e-09 0 3.018e-09 0.0007 3.021e-09 0 3.135e-09 0 3.138e-09 0.0007 3.141e-09 0 3.255e-09 0 3.258e-09 0.0007 3.261e-09 0 3.375e-09 0 3.378e-09 0.0007 3.381e-09 0 3.495e-09 0 3.498e-09 0.0007 3.501e-09 0 3.615e-09 0 3.618e-09 0.0007 3.621e-09 0 3.735e-09 0 3.738e-09 0.0007 3.741e-09 0 3.855e-09 0 3.858e-09 0.0007 3.861e-09 0 3.975e-09 0 3.978e-09 0.0007 3.981e-09 0 4.095e-09 0 4.098e-09 0.0007 4.101e-09 0 4.215e-09 0 4.218e-09 0.0007 4.221e-09 0 4.335e-09 0 4.338e-09 0.0007 4.341e-09 0 4.455e-09 0 4.458e-09 0.0007 4.461e-09 0 4.575e-09 0 4.578e-09 0.0007 4.581e-09 0 4.695e-09 0 4.698e-09 0.0007 4.701e-09 0 4.815e-09 0 4.818e-09 0.0007 4.821e-09 0 4.935e-09 0 4.938e-09 0.0007 4.941e-09 0 5.055e-09 0 5.058e-09 0.0007 5.061e-09 0 5.175e-09 0 5.178e-09 0.0007 5.181e-09 0 5.295e-09 0 5.298e-09 0.0007 5.301e-09 0 5.415e-09 0 5.418e-09 0.0007 5.421e-09 0 5.535e-09 0 5.538e-09 0.0007 5.541e-09 0 5.655e-09 0 5.658e-09 0.0007 5.661e-09 0 5.775e-09 0 5.778e-09 0.0007 5.781e-09 0 5.895e-09 0 5.898e-09 0.0007 5.901e-09 0 6.015e-09 0 6.018e-09 0.0007 6.021e-09 0 6.135e-09 0 6.138e-09 0.0007 6.141e-09 0 6.255e-09 0 6.258e-09 0.0007 6.261e-09 0 6.375e-09 0 6.378e-09 0.0007 6.381e-09 0 6.495e-09 0 6.498e-09 0.0007 6.501e-09 0 6.615e-09 0 6.618e-09 0.0007 6.621e-09 0 6.735e-09 0 6.738e-09 0.0007 6.741e-09 0 6.855e-09 0 6.858e-09 0.0007 6.861e-09 0 6.975e-09 0 6.978e-09 0.0007 6.981e-09 0 7.095e-09 0 7.098e-09 0.0007 7.101e-09 0 7.215e-09 0 7.218e-09 0.0007 7.221e-09 0 7.335e-09 0 7.338e-09 0.0007 7.341e-09 0 7.455e-09 0 7.458e-09 0.0007 7.461e-09 0 7.575e-09 0 7.578e-09 0.0007 7.581e-09 0 7.695e-09 0 7.698e-09 0.0007 7.701e-09 0 7.815e-09 0 7.818e-09 0.0007 7.821e-09 0 7.935e-09 0 7.938e-09 0.0007 7.941e-09 0 8.055e-09 0 8.058e-09 0.0007 8.061e-09 0 8.175e-09 0 8.178e-09 0.0007 8.181e-09 0 8.295e-09 0 8.298e-09 0.0007 8.301e-09 0 8.415e-09 0 8.418e-09 0.0007 8.421e-09 0 8.535e-09 0 8.538e-09 0.0007 8.541e-09 0 8.655e-09 0 8.658e-09 0.0007 8.661e-09 0 8.775e-09 0 8.778e-09 0.0007 8.781e-09 0 8.895e-09 0 8.898e-09 0.0007 8.901e-09 0 9.015e-09 0 9.018e-09 0.0007 9.021e-09 0 9.135e-09 0 9.138e-09 0.0007 9.141e-09 0 9.255e-09 0 9.258e-09 0.0007 9.261e-09 0 9.375e-09 0 9.378e-09 0.0007 9.381e-09 0 9.495e-09 0 9.498e-09 0.0007 9.501e-09 0 9.615e-09 0 9.618e-09 0.0007 9.621e-09 0 9.735e-09 0 9.738e-09 0.0007 9.741e-09 0 9.855e-09 0 9.858e-09 0.0007 9.861e-09 0 9.975e-09 0 9.978e-09 0.0007 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0007 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0007 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0007 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0007 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0007 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0007 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0007 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0007 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0007 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0007 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0007 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0007 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0007 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0007 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0007 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0007 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0007 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0007 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0007 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0007 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0007 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0007 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0007 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0007 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0007 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0007 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0007 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0007 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0007 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0007 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0007 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0007 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0007 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0007 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0007 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0007 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0007 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0007 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0007 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0007 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0007 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0007 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0007 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0007 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0007 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0007 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0007 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0007 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0007 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0007 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0007 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0007 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0007 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0007 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0007 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0007 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0007 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0007 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0007 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0007 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0007 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0007 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0007 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0007 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0007 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0007 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0007 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0007 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0007 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0007 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0007 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0007 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0007 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0007 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0007 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0007 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0007 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0007 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0007 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0007 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0007 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0007 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0007 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0007 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0007 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0007 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0007 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0007 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0007 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0007 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0007 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0007 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0007 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0007 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0007 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0007 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0007 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0007 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0007 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0007 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0007 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0007 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0007 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0007 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0007 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0007 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0007 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0007 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0007 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0007 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0007 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0007 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0007 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0007 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0007 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0007 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0007 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0007 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0007 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0007 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0007 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0007 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0007 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0007 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0007 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0007 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0007 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0007 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0007 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0007 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0007 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0007 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0007 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0007 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0007 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0007 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0007 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0007 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0007 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0007 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0007 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0007 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0007 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0007 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0007 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0007 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0007 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0007 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0007 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0007 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0007 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0007 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0007 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0007 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0007 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0007 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0007 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0007 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0007 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0007 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0007 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0007 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0007 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0007 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0007 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0007 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0007 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0007 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0007 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0007 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0007 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0007 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0007 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0007 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0007 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0007 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0007 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0007 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0007 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0007 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0007 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0007 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0007 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0007 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0007 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0007 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0007 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0007 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0007 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0007 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0007 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0007 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0007 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0007 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0007 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0007 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0007 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0007 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0007 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0007 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0007 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0007 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0007 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0007 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0007 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0007 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0007 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0007 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0007 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0007 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0007 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0007 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0007 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0007 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0007 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0007 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0007 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0007 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0007 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0007 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0007 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0007 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0007 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0007 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0007 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0007 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0007 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0007 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0007 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0007 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0007 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0007 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0007 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0007 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0007 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0007 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0007 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0007 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0007 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0007 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0007 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0007 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0007 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0007 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0007 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0007 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0007 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0007 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0007 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0007 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0007 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0007 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0007 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0007 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0007 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0007 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0007 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0007 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0007 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0007 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0007 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0007 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0007 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0007 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0007 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0007 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0007 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0007 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0007 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0007 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0007 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0007 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0007 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0007 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0007 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0007 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0007 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0007 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0007 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0007 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0007 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0007 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0007 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0007 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0007 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0007 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0007 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0007 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0007 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0007 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0007 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0007 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0007 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0007 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0007 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0007 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0007 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0007 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0007 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0007 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0007 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0007 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0007 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0007 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0007 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0007 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0007 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0007 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0007 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0007 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0007 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0007 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0007 4.7781e-08 0)
L_DFF_IP1_01|1 IP1_0_OUT _DFF_IP1_01|A1  2.067833848e-12
L_DFF_IP1_01|2 _DFF_IP1_01|A1 _DFF_IP1_01|A2  4.135667696e-12
L_DFF_IP1_01|3 _DFF_IP1_01|A3 _DFF_IP1_01|A4  8.271335392e-12
L_DFF_IP1_01|T D01 _DFF_IP1_01|T1  2.067833848e-12
L_DFF_IP1_01|4 _DFF_IP1_01|T1 _DFF_IP1_01|T2  4.135667696e-12
L_DFF_IP1_01|5 _DFF_IP1_01|A4 _DFF_IP1_01|Q1  4.135667696e-12
L_DFF_IP1_01|6 _DFF_IP1_01|Q1 IP1_1_OUT  2.067833848e-12
ID02|T 0 D02  PWL(0 0 1.5e-11 0 1.8e-11 0.0007 2.1e-11 0 1.35e-10 0 1.38e-10 0.0007 1.41e-10 0 2.55e-10 0 2.58e-10 0.0007 2.61e-10 0 3.75e-10 0 3.78e-10 0.0007 3.81e-10 0 4.95e-10 0 4.98e-10 0.0007 5.01e-10 0 6.15e-10 0 6.18e-10 0.0007 6.21e-10 0 7.35e-10 0 7.38e-10 0.0007 7.41e-10 0 8.55e-10 0 8.58e-10 0.0007 8.61e-10 0 9.75e-10 0 9.78e-10 0.0007 9.81e-10 0 1.095e-09 0 1.098e-09 0.0007 1.101e-09 0 1.215e-09 0 1.218e-09 0.0007 1.221e-09 0 1.335e-09 0 1.338e-09 0.0007 1.341e-09 0 1.455e-09 0 1.458e-09 0.0007 1.461e-09 0 1.575e-09 0 1.578e-09 0.0007 1.581e-09 0 1.695e-09 0 1.698e-09 0.0007 1.701e-09 0 1.815e-09 0 1.818e-09 0.0007 1.821e-09 0 1.935e-09 0 1.938e-09 0.0007 1.941e-09 0 2.055e-09 0 2.058e-09 0.0007 2.061e-09 0 2.175e-09 0 2.178e-09 0.0007 2.181e-09 0 2.295e-09 0 2.298e-09 0.0007 2.301e-09 0 2.415e-09 0 2.418e-09 0.0007 2.421e-09 0 2.535e-09 0 2.538e-09 0.0007 2.541e-09 0 2.655e-09 0 2.658e-09 0.0007 2.661e-09 0 2.775e-09 0 2.778e-09 0.0007 2.781e-09 0 2.895e-09 0 2.898e-09 0.0007 2.901e-09 0 3.015e-09 0 3.018e-09 0.0007 3.021e-09 0 3.135e-09 0 3.138e-09 0.0007 3.141e-09 0 3.255e-09 0 3.258e-09 0.0007 3.261e-09 0 3.375e-09 0 3.378e-09 0.0007 3.381e-09 0 3.495e-09 0 3.498e-09 0.0007 3.501e-09 0 3.615e-09 0 3.618e-09 0.0007 3.621e-09 0 3.735e-09 0 3.738e-09 0.0007 3.741e-09 0 3.855e-09 0 3.858e-09 0.0007 3.861e-09 0 3.975e-09 0 3.978e-09 0.0007 3.981e-09 0 4.095e-09 0 4.098e-09 0.0007 4.101e-09 0 4.215e-09 0 4.218e-09 0.0007 4.221e-09 0 4.335e-09 0 4.338e-09 0.0007 4.341e-09 0 4.455e-09 0 4.458e-09 0.0007 4.461e-09 0 4.575e-09 0 4.578e-09 0.0007 4.581e-09 0 4.695e-09 0 4.698e-09 0.0007 4.701e-09 0 4.815e-09 0 4.818e-09 0.0007 4.821e-09 0 4.935e-09 0 4.938e-09 0.0007 4.941e-09 0 5.055e-09 0 5.058e-09 0.0007 5.061e-09 0 5.175e-09 0 5.178e-09 0.0007 5.181e-09 0 5.295e-09 0 5.298e-09 0.0007 5.301e-09 0 5.415e-09 0 5.418e-09 0.0007 5.421e-09 0 5.535e-09 0 5.538e-09 0.0007 5.541e-09 0 5.655e-09 0 5.658e-09 0.0007 5.661e-09 0 5.775e-09 0 5.778e-09 0.0007 5.781e-09 0 5.895e-09 0 5.898e-09 0.0007 5.901e-09 0 6.015e-09 0 6.018e-09 0.0007 6.021e-09 0 6.135e-09 0 6.138e-09 0.0007 6.141e-09 0 6.255e-09 0 6.258e-09 0.0007 6.261e-09 0 6.375e-09 0 6.378e-09 0.0007 6.381e-09 0 6.495e-09 0 6.498e-09 0.0007 6.501e-09 0 6.615e-09 0 6.618e-09 0.0007 6.621e-09 0 6.735e-09 0 6.738e-09 0.0007 6.741e-09 0 6.855e-09 0 6.858e-09 0.0007 6.861e-09 0 6.975e-09 0 6.978e-09 0.0007 6.981e-09 0 7.095e-09 0 7.098e-09 0.0007 7.101e-09 0 7.215e-09 0 7.218e-09 0.0007 7.221e-09 0 7.335e-09 0 7.338e-09 0.0007 7.341e-09 0 7.455e-09 0 7.458e-09 0.0007 7.461e-09 0 7.575e-09 0 7.578e-09 0.0007 7.581e-09 0 7.695e-09 0 7.698e-09 0.0007 7.701e-09 0 7.815e-09 0 7.818e-09 0.0007 7.821e-09 0 7.935e-09 0 7.938e-09 0.0007 7.941e-09 0 8.055e-09 0 8.058e-09 0.0007 8.061e-09 0 8.175e-09 0 8.178e-09 0.0007 8.181e-09 0 8.295e-09 0 8.298e-09 0.0007 8.301e-09 0 8.415e-09 0 8.418e-09 0.0007 8.421e-09 0 8.535e-09 0 8.538e-09 0.0007 8.541e-09 0 8.655e-09 0 8.658e-09 0.0007 8.661e-09 0 8.775e-09 0 8.778e-09 0.0007 8.781e-09 0 8.895e-09 0 8.898e-09 0.0007 8.901e-09 0 9.015e-09 0 9.018e-09 0.0007 9.021e-09 0 9.135e-09 0 9.138e-09 0.0007 9.141e-09 0 9.255e-09 0 9.258e-09 0.0007 9.261e-09 0 9.375e-09 0 9.378e-09 0.0007 9.381e-09 0 9.495e-09 0 9.498e-09 0.0007 9.501e-09 0 9.615e-09 0 9.618e-09 0.0007 9.621e-09 0 9.735e-09 0 9.738e-09 0.0007 9.741e-09 0 9.855e-09 0 9.858e-09 0.0007 9.861e-09 0 9.975e-09 0 9.978e-09 0.0007 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0007 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0007 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0007 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0007 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0007 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0007 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0007 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0007 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0007 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0007 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0007 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0007 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0007 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0007 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0007 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0007 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0007 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0007 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0007 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0007 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0007 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0007 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0007 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0007 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0007 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0007 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0007 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0007 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0007 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0007 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0007 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0007 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0007 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0007 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0007 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0007 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0007 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0007 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0007 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0007 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0007 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0007 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0007 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0007 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0007 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0007 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0007 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0007 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0007 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0007 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0007 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0007 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0007 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0007 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0007 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0007 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0007 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0007 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0007 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0007 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0007 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0007 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0007 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0007 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0007 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0007 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0007 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0007 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0007 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0007 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0007 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0007 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0007 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0007 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0007 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0007 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0007 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0007 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0007 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0007 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0007 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0007 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0007 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0007 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0007 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0007 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0007 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0007 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0007 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0007 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0007 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0007 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0007 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0007 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0007 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0007 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0007 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0007 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0007 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0007 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0007 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0007 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0007 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0007 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0007 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0007 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0007 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0007 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0007 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0007 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0007 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0007 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0007 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0007 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0007 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0007 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0007 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0007 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0007 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0007 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0007 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0007 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0007 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0007 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0007 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0007 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0007 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0007 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0007 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0007 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0007 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0007 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0007 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0007 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0007 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0007 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0007 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0007 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0007 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0007 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0007 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0007 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0007 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0007 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0007 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0007 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0007 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0007 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0007 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0007 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0007 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0007 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0007 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0007 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0007 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0007 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0007 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0007 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0007 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0007 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0007 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0007 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0007 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0007 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0007 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0007 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0007 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0007 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0007 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0007 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0007 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0007 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0007 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0007 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0007 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0007 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0007 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0007 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0007 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0007 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0007 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0007 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0007 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0007 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0007 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0007 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0007 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0007 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0007 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0007 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0007 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0007 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0007 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0007 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0007 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0007 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0007 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0007 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0007 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0007 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0007 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0007 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0007 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0007 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0007 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0007 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0007 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0007 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0007 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0007 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0007 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0007 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0007 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0007 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0007 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0007 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0007 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0007 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0007 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0007 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0007 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0007 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0007 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0007 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0007 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0007 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0007 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0007 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0007 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0007 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0007 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0007 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0007 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0007 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0007 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0007 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0007 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0007 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0007 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0007 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0007 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0007 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0007 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0007 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0007 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0007 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0007 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0007 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0007 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0007 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0007 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0007 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0007 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0007 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0007 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0007 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0007 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0007 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0007 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0007 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0007 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0007 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0007 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0007 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0007 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0007 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0007 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0007 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0007 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0007 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0007 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0007 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0007 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0007 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0007 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0007 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0007 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0007 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0007 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0007 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0007 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0007 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0007 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0007 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0007 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0007 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0007 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0007 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0007 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0007 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0007 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0007 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0007 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0007 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0007 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0007 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0007 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0007 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0007 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0007 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0007 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0007 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0007 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0007 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0007 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0007 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0007 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0007 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0007 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0007 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0007 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0007 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0007 4.7781e-08 0)
L_DFF_IP2_01|1 IP2_0_OUT _DFF_IP2_01|A1  2.067833848e-12
L_DFF_IP2_01|2 _DFF_IP2_01|A1 _DFF_IP2_01|A2  4.135667696e-12
L_DFF_IP2_01|3 _DFF_IP2_01|A3 _DFF_IP2_01|A4  8.271335392e-12
L_DFF_IP2_01|T D02 _DFF_IP2_01|T1  2.067833848e-12
L_DFF_IP2_01|4 _DFF_IP2_01|T1 _DFF_IP2_01|T2  4.135667696e-12
L_DFF_IP2_01|5 _DFF_IP2_01|A4 _DFF_IP2_01|Q1  4.135667696e-12
L_DFF_IP2_01|6 _DFF_IP2_01|Q1 IP2_1_OUT  2.067833848e-12
ID03|T 0 D03  PWL(0 0 1.5e-11 0 1.8e-11 0.0007 2.1e-11 0 1.35e-10 0 1.38e-10 0.0007 1.41e-10 0 2.55e-10 0 2.58e-10 0.0007 2.61e-10 0 3.75e-10 0 3.78e-10 0.0007 3.81e-10 0 4.95e-10 0 4.98e-10 0.0007 5.01e-10 0 6.15e-10 0 6.18e-10 0.0007 6.21e-10 0 7.35e-10 0 7.38e-10 0.0007 7.41e-10 0 8.55e-10 0 8.58e-10 0.0007 8.61e-10 0 9.75e-10 0 9.78e-10 0.0007 9.81e-10 0 1.095e-09 0 1.098e-09 0.0007 1.101e-09 0 1.215e-09 0 1.218e-09 0.0007 1.221e-09 0 1.335e-09 0 1.338e-09 0.0007 1.341e-09 0 1.455e-09 0 1.458e-09 0.0007 1.461e-09 0 1.575e-09 0 1.578e-09 0.0007 1.581e-09 0 1.695e-09 0 1.698e-09 0.0007 1.701e-09 0 1.815e-09 0 1.818e-09 0.0007 1.821e-09 0 1.935e-09 0 1.938e-09 0.0007 1.941e-09 0 2.055e-09 0 2.058e-09 0.0007 2.061e-09 0 2.175e-09 0 2.178e-09 0.0007 2.181e-09 0 2.295e-09 0 2.298e-09 0.0007 2.301e-09 0 2.415e-09 0 2.418e-09 0.0007 2.421e-09 0 2.535e-09 0 2.538e-09 0.0007 2.541e-09 0 2.655e-09 0 2.658e-09 0.0007 2.661e-09 0 2.775e-09 0 2.778e-09 0.0007 2.781e-09 0 2.895e-09 0 2.898e-09 0.0007 2.901e-09 0 3.015e-09 0 3.018e-09 0.0007 3.021e-09 0 3.135e-09 0 3.138e-09 0.0007 3.141e-09 0 3.255e-09 0 3.258e-09 0.0007 3.261e-09 0 3.375e-09 0 3.378e-09 0.0007 3.381e-09 0 3.495e-09 0 3.498e-09 0.0007 3.501e-09 0 3.615e-09 0 3.618e-09 0.0007 3.621e-09 0 3.735e-09 0 3.738e-09 0.0007 3.741e-09 0 3.855e-09 0 3.858e-09 0.0007 3.861e-09 0 3.975e-09 0 3.978e-09 0.0007 3.981e-09 0 4.095e-09 0 4.098e-09 0.0007 4.101e-09 0 4.215e-09 0 4.218e-09 0.0007 4.221e-09 0 4.335e-09 0 4.338e-09 0.0007 4.341e-09 0 4.455e-09 0 4.458e-09 0.0007 4.461e-09 0 4.575e-09 0 4.578e-09 0.0007 4.581e-09 0 4.695e-09 0 4.698e-09 0.0007 4.701e-09 0 4.815e-09 0 4.818e-09 0.0007 4.821e-09 0 4.935e-09 0 4.938e-09 0.0007 4.941e-09 0 5.055e-09 0 5.058e-09 0.0007 5.061e-09 0 5.175e-09 0 5.178e-09 0.0007 5.181e-09 0 5.295e-09 0 5.298e-09 0.0007 5.301e-09 0 5.415e-09 0 5.418e-09 0.0007 5.421e-09 0 5.535e-09 0 5.538e-09 0.0007 5.541e-09 0 5.655e-09 0 5.658e-09 0.0007 5.661e-09 0 5.775e-09 0 5.778e-09 0.0007 5.781e-09 0 5.895e-09 0 5.898e-09 0.0007 5.901e-09 0 6.015e-09 0 6.018e-09 0.0007 6.021e-09 0 6.135e-09 0 6.138e-09 0.0007 6.141e-09 0 6.255e-09 0 6.258e-09 0.0007 6.261e-09 0 6.375e-09 0 6.378e-09 0.0007 6.381e-09 0 6.495e-09 0 6.498e-09 0.0007 6.501e-09 0 6.615e-09 0 6.618e-09 0.0007 6.621e-09 0 6.735e-09 0 6.738e-09 0.0007 6.741e-09 0 6.855e-09 0 6.858e-09 0.0007 6.861e-09 0 6.975e-09 0 6.978e-09 0.0007 6.981e-09 0 7.095e-09 0 7.098e-09 0.0007 7.101e-09 0 7.215e-09 0 7.218e-09 0.0007 7.221e-09 0 7.335e-09 0 7.338e-09 0.0007 7.341e-09 0 7.455e-09 0 7.458e-09 0.0007 7.461e-09 0 7.575e-09 0 7.578e-09 0.0007 7.581e-09 0 7.695e-09 0 7.698e-09 0.0007 7.701e-09 0 7.815e-09 0 7.818e-09 0.0007 7.821e-09 0 7.935e-09 0 7.938e-09 0.0007 7.941e-09 0 8.055e-09 0 8.058e-09 0.0007 8.061e-09 0 8.175e-09 0 8.178e-09 0.0007 8.181e-09 0 8.295e-09 0 8.298e-09 0.0007 8.301e-09 0 8.415e-09 0 8.418e-09 0.0007 8.421e-09 0 8.535e-09 0 8.538e-09 0.0007 8.541e-09 0 8.655e-09 0 8.658e-09 0.0007 8.661e-09 0 8.775e-09 0 8.778e-09 0.0007 8.781e-09 0 8.895e-09 0 8.898e-09 0.0007 8.901e-09 0 9.015e-09 0 9.018e-09 0.0007 9.021e-09 0 9.135e-09 0 9.138e-09 0.0007 9.141e-09 0 9.255e-09 0 9.258e-09 0.0007 9.261e-09 0 9.375e-09 0 9.378e-09 0.0007 9.381e-09 0 9.495e-09 0 9.498e-09 0.0007 9.501e-09 0 9.615e-09 0 9.618e-09 0.0007 9.621e-09 0 9.735e-09 0 9.738e-09 0.0007 9.741e-09 0 9.855e-09 0 9.858e-09 0.0007 9.861e-09 0 9.975e-09 0 9.978e-09 0.0007 9.981e-09 0 1.0095e-08 0 1.0098e-08 0.0007 1.0101e-08 0 1.0215e-08 0 1.0218e-08 0.0007 1.0221e-08 0 1.0335e-08 0 1.0338e-08 0.0007 1.0341e-08 0 1.0455e-08 0 1.0458e-08 0.0007 1.0461e-08 0 1.0575e-08 0 1.0578e-08 0.0007 1.0581e-08 0 1.0695e-08 0 1.0698e-08 0.0007 1.0701e-08 0 1.0815e-08 0 1.0818e-08 0.0007 1.0821e-08 0 1.0935e-08 0 1.0938e-08 0.0007 1.0941e-08 0 1.1055e-08 0 1.1058e-08 0.0007 1.1061e-08 0 1.1175e-08 0 1.1178e-08 0.0007 1.1181e-08 0 1.1295e-08 0 1.1298e-08 0.0007 1.1301e-08 0 1.1415e-08 0 1.1418e-08 0.0007 1.1421e-08 0 1.1535e-08 0 1.1538e-08 0.0007 1.1541e-08 0 1.1655e-08 0 1.1658e-08 0.0007 1.1661e-08 0 1.1775e-08 0 1.1778e-08 0.0007 1.1781e-08 0 1.1895e-08 0 1.1898e-08 0.0007 1.1901e-08 0 1.2015e-08 0 1.2018e-08 0.0007 1.2021e-08 0 1.2135e-08 0 1.2138e-08 0.0007 1.2141e-08 0 1.2255e-08 0 1.2258e-08 0.0007 1.2261e-08 0 1.2375e-08 0 1.2378e-08 0.0007 1.2381e-08 0 1.2495e-08 0 1.2498e-08 0.0007 1.2501e-08 0 1.2615e-08 0 1.2618e-08 0.0007 1.2621e-08 0 1.2735e-08 0 1.2738e-08 0.0007 1.2741e-08 0 1.2855e-08 0 1.2858e-08 0.0007 1.2861e-08 0 1.2975e-08 0 1.2978e-08 0.0007 1.2981e-08 0 1.3095e-08 0 1.3098e-08 0.0007 1.3101e-08 0 1.3215e-08 0 1.3218e-08 0.0007 1.3221e-08 0 1.3335e-08 0 1.3338e-08 0.0007 1.3341e-08 0 1.3455e-08 0 1.3458e-08 0.0007 1.3461e-08 0 1.3575e-08 0 1.3578e-08 0.0007 1.3581e-08 0 1.3695e-08 0 1.3698e-08 0.0007 1.3701e-08 0 1.3815e-08 0 1.3818e-08 0.0007 1.3821e-08 0 1.3935e-08 0 1.3938e-08 0.0007 1.3941e-08 0 1.4055e-08 0 1.4058e-08 0.0007 1.4061e-08 0 1.4175e-08 0 1.4178e-08 0.0007 1.4181e-08 0 1.4295e-08 0 1.4298e-08 0.0007 1.4301e-08 0 1.4415e-08 0 1.4418e-08 0.0007 1.4421e-08 0 1.4535e-08 0 1.4538e-08 0.0007 1.4541e-08 0 1.4655e-08 0 1.4658e-08 0.0007 1.4661e-08 0 1.4775e-08 0 1.4778e-08 0.0007 1.4781e-08 0 1.4895e-08 0 1.4898e-08 0.0007 1.4901e-08 0 1.5015e-08 0 1.5018e-08 0.0007 1.5021e-08 0 1.5135e-08 0 1.5138e-08 0.0007 1.5141e-08 0 1.5255e-08 0 1.5258e-08 0.0007 1.5261e-08 0 1.5375e-08 0 1.5378e-08 0.0007 1.5381e-08 0 1.5495e-08 0 1.5498e-08 0.0007 1.5501e-08 0 1.5615e-08 0 1.5618e-08 0.0007 1.5621e-08 0 1.5735e-08 0 1.5738e-08 0.0007 1.5741e-08 0 1.5855e-08 0 1.5858e-08 0.0007 1.5861e-08 0 1.5975e-08 0 1.5978e-08 0.0007 1.5981e-08 0 1.6095e-08 0 1.6098e-08 0.0007 1.6101e-08 0 1.6215e-08 0 1.6218e-08 0.0007 1.6221e-08 0 1.6335e-08 0 1.6338e-08 0.0007 1.6341e-08 0 1.6455e-08 0 1.6458e-08 0.0007 1.6461e-08 0 1.6575e-08 0 1.6578e-08 0.0007 1.6581e-08 0 1.6695e-08 0 1.6698e-08 0.0007 1.6701e-08 0 1.6815e-08 0 1.6818e-08 0.0007 1.6821e-08 0 1.6935e-08 0 1.6938e-08 0.0007 1.6941e-08 0 1.7055e-08 0 1.7058e-08 0.0007 1.7061e-08 0 1.7175e-08 0 1.7178e-08 0.0007 1.7181e-08 0 1.7295e-08 0 1.7298e-08 0.0007 1.7301e-08 0 1.7415e-08 0 1.7418e-08 0.0007 1.7421e-08 0 1.7535e-08 0 1.7538e-08 0.0007 1.7541e-08 0 1.7655e-08 0 1.7658e-08 0.0007 1.7661e-08 0 1.7775e-08 0 1.7778e-08 0.0007 1.7781e-08 0 1.7895e-08 0 1.7898e-08 0.0007 1.7901e-08 0 1.8015e-08 0 1.8018e-08 0.0007 1.8021e-08 0 1.8135e-08 0 1.8138e-08 0.0007 1.8141e-08 0 1.8255e-08 0 1.8258e-08 0.0007 1.8261e-08 0 1.8375e-08 0 1.8378e-08 0.0007 1.8381e-08 0 1.8495e-08 0 1.8498e-08 0.0007 1.8501e-08 0 1.8615e-08 0 1.8618e-08 0.0007 1.8621e-08 0 1.8735e-08 0 1.8738e-08 0.0007 1.8741e-08 0 1.8855e-08 0 1.8858e-08 0.0007 1.8861e-08 0 1.8975e-08 0 1.8978e-08 0.0007 1.8981e-08 0 1.9095e-08 0 1.9098e-08 0.0007 1.9101e-08 0 1.9215e-08 0 1.9218e-08 0.0007 1.9221e-08 0 1.9335e-08 0 1.9338e-08 0.0007 1.9341e-08 0 1.9455e-08 0 1.9458e-08 0.0007 1.9461e-08 0 1.9575e-08 0 1.9578e-08 0.0007 1.9581e-08 0 1.9695e-08 0 1.9698e-08 0.0007 1.9701e-08 0 1.9815e-08 0 1.9818e-08 0.0007 1.9821e-08 0 1.9935e-08 0 1.9938e-08 0.0007 1.9941e-08 0 2.0055e-08 0 2.0058e-08 0.0007 2.0061e-08 0 2.0175e-08 0 2.0178e-08 0.0007 2.0181e-08 0 2.0295e-08 0 2.0298e-08 0.0007 2.0301e-08 0 2.0415e-08 0 2.0418e-08 0.0007 2.0421e-08 0 2.0535e-08 0 2.0538e-08 0.0007 2.0541e-08 0 2.0655e-08 0 2.0658e-08 0.0007 2.0661e-08 0 2.0775e-08 0 2.0778e-08 0.0007 2.0781e-08 0 2.0895e-08 0 2.0898e-08 0.0007 2.0901e-08 0 2.1015e-08 0 2.1018e-08 0.0007 2.1021e-08 0 2.1135e-08 0 2.1138e-08 0.0007 2.1141e-08 0 2.1255e-08 0 2.1258e-08 0.0007 2.1261e-08 0 2.1375e-08 0 2.1378e-08 0.0007 2.1381e-08 0 2.1495e-08 0 2.1498e-08 0.0007 2.1501e-08 0 2.1615e-08 0 2.1618e-08 0.0007 2.1621e-08 0 2.1735e-08 0 2.1738e-08 0.0007 2.1741e-08 0 2.1855e-08 0 2.1858e-08 0.0007 2.1861e-08 0 2.1975e-08 0 2.1978e-08 0.0007 2.1981e-08 0 2.2095e-08 0 2.2098e-08 0.0007 2.2101e-08 0 2.2215e-08 0 2.2218e-08 0.0007 2.2221e-08 0 2.2335e-08 0 2.2338e-08 0.0007 2.2341e-08 0 2.2455e-08 0 2.2458e-08 0.0007 2.2461e-08 0 2.2575e-08 0 2.2578e-08 0.0007 2.2581e-08 0 2.2695e-08 0 2.2698e-08 0.0007 2.2701e-08 0 2.2815e-08 0 2.2818e-08 0.0007 2.2821e-08 0 2.2935e-08 0 2.2938e-08 0.0007 2.2941e-08 0 2.3055e-08 0 2.3058e-08 0.0007 2.3061e-08 0 2.3175e-08 0 2.3178e-08 0.0007 2.3181e-08 0 2.3295e-08 0 2.3298e-08 0.0007 2.3301e-08 0 2.3415e-08 0 2.3418e-08 0.0007 2.3421e-08 0 2.3535e-08 0 2.3538e-08 0.0007 2.3541e-08 0 2.3655e-08 0 2.3658e-08 0.0007 2.3661e-08 0 2.3775e-08 0 2.3778e-08 0.0007 2.3781e-08 0 2.3895e-08 0 2.3898e-08 0.0007 2.3901e-08 0 2.4015e-08 0 2.4018e-08 0.0007 2.4021e-08 0 2.4135e-08 0 2.4138e-08 0.0007 2.4141e-08 0 2.4255e-08 0 2.4258e-08 0.0007 2.4261e-08 0 2.4375e-08 0 2.4378e-08 0.0007 2.4381e-08 0 2.4495e-08 0 2.4498e-08 0.0007 2.4501e-08 0 2.4615e-08 0 2.4618e-08 0.0007 2.4621e-08 0 2.4735e-08 0 2.4738e-08 0.0007 2.4741e-08 0 2.4855e-08 0 2.4858e-08 0.0007 2.4861e-08 0 2.4975e-08 0 2.4978e-08 0.0007 2.4981e-08 0 2.5095e-08 0 2.5098e-08 0.0007 2.5101e-08 0 2.5215e-08 0 2.5218e-08 0.0007 2.5221e-08 0 2.5335e-08 0 2.5338e-08 0.0007 2.5341e-08 0 2.5455e-08 0 2.5458e-08 0.0007 2.5461e-08 0 2.5575e-08 0 2.5578e-08 0.0007 2.5581e-08 0 2.5695e-08 0 2.5698e-08 0.0007 2.5701e-08 0 2.5815e-08 0 2.5818e-08 0.0007 2.5821e-08 0 2.5935e-08 0 2.5938e-08 0.0007 2.5941e-08 0 2.6055e-08 0 2.6058e-08 0.0007 2.6061e-08 0 2.6175e-08 0 2.6178e-08 0.0007 2.6181e-08 0 2.6295e-08 0 2.6298e-08 0.0007 2.6301e-08 0 2.6415e-08 0 2.6418e-08 0.0007 2.6421e-08 0 2.6535e-08 0 2.6538e-08 0.0007 2.6541e-08 0 2.6655e-08 0 2.6658e-08 0.0007 2.6661e-08 0 2.6775e-08 0 2.6778e-08 0.0007 2.6781e-08 0 2.6895e-08 0 2.6898e-08 0.0007 2.6901e-08 0 2.7015e-08 0 2.7018e-08 0.0007 2.7021e-08 0 2.7135e-08 0 2.7138e-08 0.0007 2.7141e-08 0 2.7255e-08 0 2.7258e-08 0.0007 2.7261e-08 0 2.7375e-08 0 2.7378e-08 0.0007 2.7381e-08 0 2.7495e-08 0 2.7498e-08 0.0007 2.7501e-08 0 2.7615e-08 0 2.7618e-08 0.0007 2.7621e-08 0 2.7735e-08 0 2.7738e-08 0.0007 2.7741e-08 0 2.7855e-08 0 2.7858e-08 0.0007 2.7861e-08 0 2.7975e-08 0 2.7978e-08 0.0007 2.7981e-08 0 2.8095e-08 0 2.8098e-08 0.0007 2.8101e-08 0 2.8215e-08 0 2.8218e-08 0.0007 2.8221e-08 0 2.8335e-08 0 2.8338e-08 0.0007 2.8341e-08 0 2.8455e-08 0 2.8458e-08 0.0007 2.8461e-08 0 2.8575e-08 0 2.8578e-08 0.0007 2.8581e-08 0 2.8695e-08 0 2.8698e-08 0.0007 2.8701e-08 0 2.8815e-08 0 2.8818e-08 0.0007 2.8821e-08 0 2.8935e-08 0 2.8938e-08 0.0007 2.8941e-08 0 2.9055e-08 0 2.9058e-08 0.0007 2.9061e-08 0 2.9175e-08 0 2.9178e-08 0.0007 2.9181e-08 0 2.9295e-08 0 2.9298e-08 0.0007 2.9301e-08 0 2.9415e-08 0 2.9418e-08 0.0007 2.9421e-08 0 2.9535e-08 0 2.9538e-08 0.0007 2.9541e-08 0 2.9655e-08 0 2.9658e-08 0.0007 2.9661e-08 0 2.9775e-08 0 2.9778e-08 0.0007 2.9781e-08 0 2.9895e-08 0 2.9898e-08 0.0007 2.9901e-08 0 3.0015e-08 0 3.0018e-08 0.0007 3.0021e-08 0 3.0135e-08 0 3.0138e-08 0.0007 3.0141e-08 0 3.0255e-08 0 3.0258e-08 0.0007 3.0261e-08 0 3.0375e-08 0 3.0378e-08 0.0007 3.0381e-08 0 3.0495e-08 0 3.0498e-08 0.0007 3.0501e-08 0 3.0615e-08 0 3.0618e-08 0.0007 3.0621e-08 0 3.0735e-08 0 3.0738e-08 0.0007 3.0741e-08 0 3.0855e-08 0 3.0858e-08 0.0007 3.0861e-08 0 3.0975e-08 0 3.0978e-08 0.0007 3.0981e-08 0 3.1095e-08 0 3.1098e-08 0.0007 3.1101e-08 0 3.1215e-08 0 3.1218e-08 0.0007 3.1221e-08 0 3.1335e-08 0 3.1338e-08 0.0007 3.1341e-08 0 3.1455e-08 0 3.1458e-08 0.0007 3.1461e-08 0 3.1575e-08 0 3.1578e-08 0.0007 3.1581e-08 0 3.1695e-08 0 3.1698e-08 0.0007 3.1701e-08 0 3.1815e-08 0 3.1818e-08 0.0007 3.1821e-08 0 3.1935e-08 0 3.1938e-08 0.0007 3.1941e-08 0 3.2055e-08 0 3.2058e-08 0.0007 3.2061e-08 0 3.2175e-08 0 3.2178e-08 0.0007 3.2181e-08 0 3.2295e-08 0 3.2298e-08 0.0007 3.2301e-08 0 3.2415e-08 0 3.2418e-08 0.0007 3.2421e-08 0 3.2535e-08 0 3.2538e-08 0.0007 3.2541e-08 0 3.2655e-08 0 3.2658e-08 0.0007 3.2661e-08 0 3.2775e-08 0 3.2778e-08 0.0007 3.2781e-08 0 3.2895e-08 0 3.2898e-08 0.0007 3.2901e-08 0 3.3015e-08 0 3.3018e-08 0.0007 3.3021e-08 0 3.3135e-08 0 3.3138e-08 0.0007 3.3141e-08 0 3.3255e-08 0 3.3258e-08 0.0007 3.3261e-08 0 3.3375e-08 0 3.3378e-08 0.0007 3.3381e-08 0 3.3495e-08 0 3.3498e-08 0.0007 3.3501e-08 0 3.3615e-08 0 3.3618e-08 0.0007 3.3621e-08 0 3.3735e-08 0 3.3738e-08 0.0007 3.3741e-08 0 3.3855e-08 0 3.3858e-08 0.0007 3.3861e-08 0 3.3975e-08 0 3.3978e-08 0.0007 3.3981e-08 0 3.4095e-08 0 3.4098e-08 0.0007 3.4101e-08 0 3.4215e-08 0 3.4218e-08 0.0007 3.4221e-08 0 3.4335e-08 0 3.4338e-08 0.0007 3.4341e-08 0 3.4455e-08 0 3.4458e-08 0.0007 3.4461e-08 0 3.4575e-08 0 3.4578e-08 0.0007 3.4581e-08 0 3.4695e-08 0 3.4698e-08 0.0007 3.4701e-08 0 3.4815e-08 0 3.4818e-08 0.0007 3.4821e-08 0 3.4935e-08 0 3.4938e-08 0.0007 3.4941e-08 0 3.5055e-08 0 3.5058e-08 0.0007 3.5061e-08 0 3.5175e-08 0 3.5178e-08 0.0007 3.5181e-08 0 3.5295e-08 0 3.5298e-08 0.0007 3.5301e-08 0 3.5415e-08 0 3.5418e-08 0.0007 3.5421e-08 0 3.5535e-08 0 3.5538e-08 0.0007 3.5541e-08 0 3.5655e-08 0 3.5658e-08 0.0007 3.5661e-08 0 3.5775e-08 0 3.5778e-08 0.0007 3.5781e-08 0 3.5895e-08 0 3.5898e-08 0.0007 3.5901e-08 0 3.6015e-08 0 3.6018e-08 0.0007 3.6021e-08 0 3.6135e-08 0 3.6138e-08 0.0007 3.6141e-08 0 3.6255e-08 0 3.6258e-08 0.0007 3.6261e-08 0 3.6375e-08 0 3.6378e-08 0.0007 3.6381e-08 0 3.6495e-08 0 3.6498e-08 0.0007 3.6501e-08 0 3.6615e-08 0 3.6618e-08 0.0007 3.6621e-08 0 3.6735e-08 0 3.6738e-08 0.0007 3.6741e-08 0 3.6855e-08 0 3.6858e-08 0.0007 3.6861e-08 0 3.6975e-08 0 3.6978e-08 0.0007 3.6981e-08 0 3.7095e-08 0 3.7098e-08 0.0007 3.7101e-08 0 3.7215e-08 0 3.7218e-08 0.0007 3.7221e-08 0 3.7335e-08 0 3.7338e-08 0.0007 3.7341e-08 0 3.7455e-08 0 3.7458e-08 0.0007 3.7461e-08 0 3.7575e-08 0 3.7578e-08 0.0007 3.7581e-08 0 3.7695e-08 0 3.7698e-08 0.0007 3.7701e-08 0 3.7815e-08 0 3.7818e-08 0.0007 3.7821e-08 0 3.7935e-08 0 3.7938e-08 0.0007 3.7941e-08 0 3.8055e-08 0 3.8058e-08 0.0007 3.8061e-08 0 3.8175e-08 0 3.8178e-08 0.0007 3.8181e-08 0 3.8295e-08 0 3.8298e-08 0.0007 3.8301e-08 0 3.8415e-08 0 3.8418e-08 0.0007 3.8421e-08 0 3.8535e-08 0 3.8538e-08 0.0007 3.8541e-08 0 3.8655e-08 0 3.8658e-08 0.0007 3.8661e-08 0 3.8775e-08 0 3.8778e-08 0.0007 3.8781e-08 0 3.8895e-08 0 3.8898e-08 0.0007 3.8901e-08 0 3.9015e-08 0 3.9018e-08 0.0007 3.9021e-08 0 3.9135e-08 0 3.9138e-08 0.0007 3.9141e-08 0 3.9255e-08 0 3.9258e-08 0.0007 3.9261e-08 0 3.9375e-08 0 3.9378e-08 0.0007 3.9381e-08 0 3.9495e-08 0 3.9498e-08 0.0007 3.9501e-08 0 3.9615e-08 0 3.9618e-08 0.0007 3.9621e-08 0 3.9735e-08 0 3.9738e-08 0.0007 3.9741e-08 0 3.9855e-08 0 3.9858e-08 0.0007 3.9861e-08 0 3.9975e-08 0 3.9978e-08 0.0007 3.9981e-08 0 4.0095e-08 0 4.0098e-08 0.0007 4.0101e-08 0 4.0215e-08 0 4.0218e-08 0.0007 4.0221e-08 0 4.0335e-08 0 4.0338e-08 0.0007 4.0341e-08 0 4.0455e-08 0 4.0458e-08 0.0007 4.0461e-08 0 4.0575e-08 0 4.0578e-08 0.0007 4.0581e-08 0 4.0695e-08 0 4.0698e-08 0.0007 4.0701e-08 0 4.0815e-08 0 4.0818e-08 0.0007 4.0821e-08 0 4.0935e-08 0 4.0938e-08 0.0007 4.0941e-08 0 4.1055e-08 0 4.1058e-08 0.0007 4.1061e-08 0 4.1175e-08 0 4.1178e-08 0.0007 4.1181e-08 0 4.1295e-08 0 4.1298e-08 0.0007 4.1301e-08 0 4.1415e-08 0 4.1418e-08 0.0007 4.1421e-08 0 4.1535e-08 0 4.1538e-08 0.0007 4.1541e-08 0 4.1655e-08 0 4.1658e-08 0.0007 4.1661e-08 0 4.1775e-08 0 4.1778e-08 0.0007 4.1781e-08 0 4.1895e-08 0 4.1898e-08 0.0007 4.1901e-08 0 4.2015e-08 0 4.2018e-08 0.0007 4.2021e-08 0 4.2135e-08 0 4.2138e-08 0.0007 4.2141e-08 0 4.2255e-08 0 4.2258e-08 0.0007 4.2261e-08 0 4.2375e-08 0 4.2378e-08 0.0007 4.2381e-08 0 4.2495e-08 0 4.2498e-08 0.0007 4.2501e-08 0 4.2615e-08 0 4.2618e-08 0.0007 4.2621e-08 0 4.2735e-08 0 4.2738e-08 0.0007 4.2741e-08 0 4.2855e-08 0 4.2858e-08 0.0007 4.2861e-08 0 4.2975e-08 0 4.2978e-08 0.0007 4.2981e-08 0 4.3095e-08 0 4.3098e-08 0.0007 4.3101e-08 0 4.3215e-08 0 4.3218e-08 0.0007 4.3221e-08 0 4.3335e-08 0 4.3338e-08 0.0007 4.3341e-08 0 4.3455e-08 0 4.3458e-08 0.0007 4.3461e-08 0 4.3575e-08 0 4.3578e-08 0.0007 4.3581e-08 0 4.3695e-08 0 4.3698e-08 0.0007 4.3701e-08 0 4.3815e-08 0 4.3818e-08 0.0007 4.3821e-08 0 4.3935e-08 0 4.3938e-08 0.0007 4.3941e-08 0 4.4055e-08 0 4.4058e-08 0.0007 4.4061e-08 0 4.4175e-08 0 4.4178e-08 0.0007 4.4181e-08 0 4.4295e-08 0 4.4298e-08 0.0007 4.4301e-08 0 4.4415e-08 0 4.4418e-08 0.0007 4.4421e-08 0 4.4535e-08 0 4.4538e-08 0.0007 4.4541e-08 0 4.4655e-08 0 4.4658e-08 0.0007 4.4661e-08 0 4.4775e-08 0 4.4778e-08 0.0007 4.4781e-08 0 4.4895e-08 0 4.4898e-08 0.0007 4.4901e-08 0 4.5015e-08 0 4.5018e-08 0.0007 4.5021e-08 0 4.5135e-08 0 4.5138e-08 0.0007 4.5141e-08 0 4.5255e-08 0 4.5258e-08 0.0007 4.5261e-08 0 4.5375e-08 0 4.5378e-08 0.0007 4.5381e-08 0 4.5495e-08 0 4.5498e-08 0.0007 4.5501e-08 0 4.5615e-08 0 4.5618e-08 0.0007 4.5621e-08 0 4.5735e-08 0 4.5738e-08 0.0007 4.5741e-08 0 4.5855e-08 0 4.5858e-08 0.0007 4.5861e-08 0 4.5975e-08 0 4.5978e-08 0.0007 4.5981e-08 0 4.6095e-08 0 4.6098e-08 0.0007 4.6101e-08 0 4.6215e-08 0 4.6218e-08 0.0007 4.6221e-08 0 4.6335e-08 0 4.6338e-08 0.0007 4.6341e-08 0 4.6455e-08 0 4.6458e-08 0.0007 4.6461e-08 0 4.6575e-08 0 4.6578e-08 0.0007 4.6581e-08 0 4.6695e-08 0 4.6698e-08 0.0007 4.6701e-08 0 4.6815e-08 0 4.6818e-08 0.0007 4.6821e-08 0 4.6935e-08 0 4.6938e-08 0.0007 4.6941e-08 0 4.7055e-08 0 4.7058e-08 0.0007 4.7061e-08 0 4.7175e-08 0 4.7178e-08 0.0007 4.7181e-08 0 4.7295e-08 0 4.7298e-08 0.0007 4.7301e-08 0 4.7415e-08 0 4.7418e-08 0.0007 4.7421e-08 0 4.7535e-08 0 4.7538e-08 0.0007 4.7541e-08 0 4.7655e-08 0 4.7658e-08 0.0007 4.7661e-08 0 4.7775e-08 0 4.7778e-08 0.0007 4.7781e-08 0)
L_DFF_IP3_01|1 IP3_0_OUT _DFF_IP3_01|A1  2.067833848e-12
L_DFF_IP3_01|2 _DFF_IP3_01|A1 _DFF_IP3_01|A2  4.135667696e-12
L_DFF_IP3_01|3 _DFF_IP3_01|A3 _DFF_IP3_01|A4  8.271335392e-12
L_DFF_IP3_01|T D03 _DFF_IP3_01|T1  2.067833848e-12
L_DFF_IP3_01|4 _DFF_IP3_01|T1 _DFF_IP3_01|T2  4.135667696e-12
L_DFF_IP3_01|5 _DFF_IP3_01|A4 _DFF_IP3_01|Q1  4.135667696e-12
L_DFF_IP3_01|6 _DFF_IP3_01|Q1 IP3_1_OUT  2.067833848e-12
IT08|T 0 T08  PWL(0 0 9e-12 0 1.2e-11 0.0014 1.5e-11 0 1.29e-10 0 1.32e-10 0.0014 1.35e-10 0 2.49e-10 0 2.52e-10 0.0014 2.55e-10 0 3.69e-10 0 3.72e-10 0.0014 3.75e-10 0 4.89e-10 0 4.92e-10 0.0014 4.95e-10 0 6.09e-10 0 6.12e-10 0.0014 6.15e-10 0 7.29e-10 0 7.32e-10 0.0014 7.35e-10 0 8.49e-10 0 8.52e-10 0.0014 8.55e-10 0 9.69e-10 0 9.72e-10 0.0014 9.75e-10 0 1.089e-09 0 1.092e-09 0.0014 1.095e-09 0 1.209e-09 0 1.212e-09 0.0014 1.215e-09 0 1.329e-09 0 1.332e-09 0.0014 1.335e-09 0 1.449e-09 0 1.452e-09 0.0014 1.455e-09 0 1.569e-09 0 1.572e-09 0.0014 1.575e-09 0 1.689e-09 0 1.692e-09 0.0014 1.695e-09 0 1.809e-09 0 1.812e-09 0.0014 1.815e-09 0 1.929e-09 0 1.932e-09 0.0014 1.935e-09 0 2.049e-09 0 2.052e-09 0.0014 2.055e-09 0 2.169e-09 0 2.172e-09 0.0014 2.175e-09 0 2.289e-09 0 2.292e-09 0.0014 2.295e-09 0 2.409e-09 0 2.412e-09 0.0014 2.415e-09 0 2.529e-09 0 2.532e-09 0.0014 2.535e-09 0 2.649e-09 0 2.652e-09 0.0014 2.655e-09 0 2.769e-09 0 2.772e-09 0.0014 2.775e-09 0 2.889e-09 0 2.892e-09 0.0014 2.895e-09 0 3.009e-09 0 3.012e-09 0.0014 3.015e-09 0 3.129e-09 0 3.132e-09 0.0014 3.135e-09 0 3.249e-09 0 3.252e-09 0.0014 3.255e-09 0 3.369e-09 0 3.372e-09 0.0014 3.375e-09 0 3.489e-09 0 3.492e-09 0.0014 3.495e-09 0 3.609e-09 0 3.612e-09 0.0014 3.615e-09 0 3.729e-09 0 3.732e-09 0.0014 3.735e-09 0 3.849e-09 0 3.852e-09 0.0014 3.855e-09 0 3.969e-09 0 3.972e-09 0.0014 3.975e-09 0 4.089e-09 0 4.092e-09 0.0014 4.095e-09 0 4.209e-09 0 4.212e-09 0.0014 4.215e-09 0 4.329e-09 0 4.332e-09 0.0014 4.335e-09 0 4.449e-09 0 4.452e-09 0.0014 4.455e-09 0 4.569e-09 0 4.572e-09 0.0014 4.575e-09 0 4.689e-09 0 4.692e-09 0.0014 4.695e-09 0 4.809e-09 0 4.812e-09 0.0014 4.815e-09 0 4.929e-09 0 4.932e-09 0.0014 4.935e-09 0 5.049e-09 0 5.052e-09 0.0014 5.055e-09 0 5.169e-09 0 5.172e-09 0.0014 5.175e-09 0 5.289e-09 0 5.292e-09 0.0014 5.295e-09 0 5.409e-09 0 5.412e-09 0.0014 5.415e-09 0 5.529e-09 0 5.532e-09 0.0014 5.535e-09 0 5.649e-09 0 5.652e-09 0.0014 5.655e-09 0 5.769e-09 0 5.772e-09 0.0014 5.775e-09 0 5.889e-09 0 5.892e-09 0.0014 5.895e-09 0 6.009e-09 0 6.012e-09 0.0014 6.015e-09 0 6.129e-09 0 6.132e-09 0.0014 6.135e-09 0 6.249e-09 0 6.252e-09 0.0014 6.255e-09 0 6.369e-09 0 6.372e-09 0.0014 6.375e-09 0 6.489e-09 0 6.492e-09 0.0014 6.495e-09 0 6.609e-09 0 6.612e-09 0.0014 6.615e-09 0 6.729e-09 0 6.732e-09 0.0014 6.735e-09 0 6.849e-09 0 6.852e-09 0.0014 6.855e-09 0 6.969e-09 0 6.972e-09 0.0014 6.975e-09 0 7.089e-09 0 7.092e-09 0.0014 7.095e-09 0 7.209e-09 0 7.212e-09 0.0014 7.215e-09 0 7.329e-09 0 7.332e-09 0.0014 7.335e-09 0 7.449e-09 0 7.452e-09 0.0014 7.455e-09 0 7.569e-09 0 7.572e-09 0.0014 7.575e-09 0 7.689e-09 0 7.692e-09 0.0014 7.695e-09 0 7.809e-09 0 7.812e-09 0.0014 7.815e-09 0 7.929e-09 0 7.932e-09 0.0014 7.935e-09 0 8.049e-09 0 8.052e-09 0.0014 8.055e-09 0 8.169e-09 0 8.172e-09 0.0014 8.175e-09 0 8.289e-09 0 8.292e-09 0.0014 8.295e-09 0 8.409e-09 0 8.412e-09 0.0014 8.415e-09 0 8.529e-09 0 8.532e-09 0.0014 8.535e-09 0 8.649e-09 0 8.652e-09 0.0014 8.655e-09 0 8.769e-09 0 8.772e-09 0.0014 8.775e-09 0 8.889e-09 0 8.892e-09 0.0014 8.895e-09 0 9.009e-09 0 9.012e-09 0.0014 9.015e-09 0 9.129e-09 0 9.132e-09 0.0014 9.135e-09 0 9.249e-09 0 9.252e-09 0.0014 9.255e-09 0 9.369e-09 0 9.372e-09 0.0014 9.375e-09 0 9.489e-09 0 9.492e-09 0.0014 9.495e-09 0 9.609e-09 0 9.612e-09 0.0014 9.615e-09 0 9.729e-09 0 9.732e-09 0.0014 9.735e-09 0 9.849e-09 0 9.852e-09 0.0014 9.855e-09 0 9.969e-09 0 9.972e-09 0.0014 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0014 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0014 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0014 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0014 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0014 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0014 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0014 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0014 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0014 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0014 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0014 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0014 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0014 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0014 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0014 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0014 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0014 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0014 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0014 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0014 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0014 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0014 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0014 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0014 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0014 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0014 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0014 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0014 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0014 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0014 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0014 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0014 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0014 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0014 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0014 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0014 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0014 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0014 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0014 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0014 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0014 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0014 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0014 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0014 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0014 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0014 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0014 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0014 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0014 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0014 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0014 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0014 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0014 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0014 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0014 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0014 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0014 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0014 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0014 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0014 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0014 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0014 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0014 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0014 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0014 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0014 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0014 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0014 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0014 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0014 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0014 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0014 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0014 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0014 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0014 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0014 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0014 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0014 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0014 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0014 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0014 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0014 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0014 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0014 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0014 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0014 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0014 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0014 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0014 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0014 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0014 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0014 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0014 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0014 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0014 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0014 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0014 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0014 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0014 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0014 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0014 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0014 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0014 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0014 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0014 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0014 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0014 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0014 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0014 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0014 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0014 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0014 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0014 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0014 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0014 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0014 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0014 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0014 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0014 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0014 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0014 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0014 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0014 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0014 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0014 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0014 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0014 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0014 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0014 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0014 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0014 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0014 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0014 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0014 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0014 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0014 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0014 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0014 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0014 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0014 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0014 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0014 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0014 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0014 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0014 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0014 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0014 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0014 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0014 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0014 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0014 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0014 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0014 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0014 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0014 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0014 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0014 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0014 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0014 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0014 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0014 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0014 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0014 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0014 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0014 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0014 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0014 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0014 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0014 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0014 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0014 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0014 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0014 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0014 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0014 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0014 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0014 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0014 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0014 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0014 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0014 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0014 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0014 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0014 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0014 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0014 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0014 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0014 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0014 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0014 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0014 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0014 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0014 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0014 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0014 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0014 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0014 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0014 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0014 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0014 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0014 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0014 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0014 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0014 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0014 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0014 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0014 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0014 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0014 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0014 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0014 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0014 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0014 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0014 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0014 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0014 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0014 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0014 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0014 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0014 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0014 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0014 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0014 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0014 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0014 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0014 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0014 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0014 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0014 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0014 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0014 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0014 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0014 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0014 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0014 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0014 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0014 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0014 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0014 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0014 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0014 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0014 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0014 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0014 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0014 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0014 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0014 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0014 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0014 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0014 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0014 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0014 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0014 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0014 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0014 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0014 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0014 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0014 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0014 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0014 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0014 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0014 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0014 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0014 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0014 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0014 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0014 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0014 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0014 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0014 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0014 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0014 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0014 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0014 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0014 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0014 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0014 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0014 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0014 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0014 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0014 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0014 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0014 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0014 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0014 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0014 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0014 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0014 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0014 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0014 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0014 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0014 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0014 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0014 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0014 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0014 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0014 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0014 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0014 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0014 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0014 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0014 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0014 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0014 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0014 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0014 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0014 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0014 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0014 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0014 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0014 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0014 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0014 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0014 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0014 4.7775e-08 0)
IT09|T 0 T09  PWL(0 0 9e-12 0 1.2e-11 0.0007 1.5e-11 0 1.29e-10 0 1.32e-10 0.0007 1.35e-10 0 2.49e-10 0 2.52e-10 0.0007 2.55e-10 0 3.69e-10 0 3.72e-10 0.0007 3.75e-10 0 4.89e-10 0 4.92e-10 0.0007 4.95e-10 0 6.09e-10 0 6.12e-10 0.0007 6.15e-10 0 7.29e-10 0 7.32e-10 0.0007 7.35e-10 0 8.49e-10 0 8.52e-10 0.0007 8.55e-10 0 9.69e-10 0 9.72e-10 0.0007 9.75e-10 0 1.089e-09 0 1.092e-09 0.0007 1.095e-09 0 1.209e-09 0 1.212e-09 0.0007 1.215e-09 0 1.329e-09 0 1.332e-09 0.0007 1.335e-09 0 1.449e-09 0 1.452e-09 0.0007 1.455e-09 0 1.569e-09 0 1.572e-09 0.0007 1.575e-09 0 1.689e-09 0 1.692e-09 0.0007 1.695e-09 0 1.809e-09 0 1.812e-09 0.0007 1.815e-09 0 1.929e-09 0 1.932e-09 0.0007 1.935e-09 0 2.049e-09 0 2.052e-09 0.0007 2.055e-09 0 2.169e-09 0 2.172e-09 0.0007 2.175e-09 0 2.289e-09 0 2.292e-09 0.0007 2.295e-09 0 2.409e-09 0 2.412e-09 0.0007 2.415e-09 0 2.529e-09 0 2.532e-09 0.0007 2.535e-09 0 2.649e-09 0 2.652e-09 0.0007 2.655e-09 0 2.769e-09 0 2.772e-09 0.0007 2.775e-09 0 2.889e-09 0 2.892e-09 0.0007 2.895e-09 0 3.009e-09 0 3.012e-09 0.0007 3.015e-09 0 3.129e-09 0 3.132e-09 0.0007 3.135e-09 0 3.249e-09 0 3.252e-09 0.0007 3.255e-09 0 3.369e-09 0 3.372e-09 0.0007 3.375e-09 0 3.489e-09 0 3.492e-09 0.0007 3.495e-09 0 3.609e-09 0 3.612e-09 0.0007 3.615e-09 0 3.729e-09 0 3.732e-09 0.0007 3.735e-09 0 3.849e-09 0 3.852e-09 0.0007 3.855e-09 0 3.969e-09 0 3.972e-09 0.0007 3.975e-09 0 4.089e-09 0 4.092e-09 0.0007 4.095e-09 0 4.209e-09 0 4.212e-09 0.0007 4.215e-09 0 4.329e-09 0 4.332e-09 0.0007 4.335e-09 0 4.449e-09 0 4.452e-09 0.0007 4.455e-09 0 4.569e-09 0 4.572e-09 0.0007 4.575e-09 0 4.689e-09 0 4.692e-09 0.0007 4.695e-09 0 4.809e-09 0 4.812e-09 0.0007 4.815e-09 0 4.929e-09 0 4.932e-09 0.0007 4.935e-09 0 5.049e-09 0 5.052e-09 0.0007 5.055e-09 0 5.169e-09 0 5.172e-09 0.0007 5.175e-09 0 5.289e-09 0 5.292e-09 0.0007 5.295e-09 0 5.409e-09 0 5.412e-09 0.0007 5.415e-09 0 5.529e-09 0 5.532e-09 0.0007 5.535e-09 0 5.649e-09 0 5.652e-09 0.0007 5.655e-09 0 5.769e-09 0 5.772e-09 0.0007 5.775e-09 0 5.889e-09 0 5.892e-09 0.0007 5.895e-09 0 6.009e-09 0 6.012e-09 0.0007 6.015e-09 0 6.129e-09 0 6.132e-09 0.0007 6.135e-09 0 6.249e-09 0 6.252e-09 0.0007 6.255e-09 0 6.369e-09 0 6.372e-09 0.0007 6.375e-09 0 6.489e-09 0 6.492e-09 0.0007 6.495e-09 0 6.609e-09 0 6.612e-09 0.0007 6.615e-09 0 6.729e-09 0 6.732e-09 0.0007 6.735e-09 0 6.849e-09 0 6.852e-09 0.0007 6.855e-09 0 6.969e-09 0 6.972e-09 0.0007 6.975e-09 0 7.089e-09 0 7.092e-09 0.0007 7.095e-09 0 7.209e-09 0 7.212e-09 0.0007 7.215e-09 0 7.329e-09 0 7.332e-09 0.0007 7.335e-09 0 7.449e-09 0 7.452e-09 0.0007 7.455e-09 0 7.569e-09 0 7.572e-09 0.0007 7.575e-09 0 7.689e-09 0 7.692e-09 0.0007 7.695e-09 0 7.809e-09 0 7.812e-09 0.0007 7.815e-09 0 7.929e-09 0 7.932e-09 0.0007 7.935e-09 0 8.049e-09 0 8.052e-09 0.0007 8.055e-09 0 8.169e-09 0 8.172e-09 0.0007 8.175e-09 0 8.289e-09 0 8.292e-09 0.0007 8.295e-09 0 8.409e-09 0 8.412e-09 0.0007 8.415e-09 0 8.529e-09 0 8.532e-09 0.0007 8.535e-09 0 8.649e-09 0 8.652e-09 0.0007 8.655e-09 0 8.769e-09 0 8.772e-09 0.0007 8.775e-09 0 8.889e-09 0 8.892e-09 0.0007 8.895e-09 0 9.009e-09 0 9.012e-09 0.0007 9.015e-09 0 9.129e-09 0 9.132e-09 0.0007 9.135e-09 0 9.249e-09 0 9.252e-09 0.0007 9.255e-09 0 9.369e-09 0 9.372e-09 0.0007 9.375e-09 0 9.489e-09 0 9.492e-09 0.0007 9.495e-09 0 9.609e-09 0 9.612e-09 0.0007 9.615e-09 0 9.729e-09 0 9.732e-09 0.0007 9.735e-09 0 9.849e-09 0 9.852e-09 0.0007 9.855e-09 0 9.969e-09 0 9.972e-09 0.0007 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0007 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0007 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0007 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0007 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0007 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0007 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0007 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0007 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0007 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0007 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0007 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0007 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0007 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0007 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0007 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0007 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0007 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0007 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0007 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0007 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0007 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0007 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0007 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0007 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0007 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0007 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0007 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0007 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0007 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0007 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0007 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0007 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0007 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0007 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0007 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0007 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0007 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0007 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0007 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0007 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0007 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0007 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0007 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0007 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0007 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0007 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0007 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0007 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0007 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0007 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0007 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0007 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0007 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0007 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0007 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0007 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0007 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0007 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0007 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0007 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0007 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0007 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0007 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0007 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0007 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0007 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0007 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0007 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0007 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0007 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0007 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0007 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0007 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0007 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0007 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0007 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0007 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0007 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0007 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0007 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0007 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0007 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0007 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0007 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0007 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0007 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0007 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0007 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0007 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0007 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0007 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0007 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0007 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0007 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0007 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0007 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0007 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0007 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0007 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0007 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0007 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0007 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0007 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0007 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0007 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0007 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0007 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0007 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0007 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0007 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0007 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0007 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0007 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0007 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0007 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0007 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0007 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0007 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0007 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0007 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0007 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0007 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0007 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0007 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0007 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0007 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0007 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0007 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0007 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0007 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0007 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0007 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0007 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0007 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0007 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0007 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0007 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0007 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0007 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0007 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0007 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0007 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0007 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0007 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0007 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0007 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0007 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0007 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0007 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0007 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0007 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0007 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0007 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0007 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0007 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0007 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0007 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0007 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0007 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0007 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0007 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0007 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0007 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0007 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0007 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0007 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0007 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0007 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0007 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0007 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0007 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0007 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0007 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0007 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0007 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0007 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0007 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0007 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0007 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0007 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0007 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0007 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0007 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0007 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0007 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0007 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0007 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0007 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0007 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0007 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0007 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0007 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0007 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0007 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0007 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0007 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0007 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0007 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0007 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0007 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0007 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0007 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0007 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0007 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0007 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0007 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0007 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0007 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0007 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0007 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0007 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0007 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0007 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0007 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0007 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0007 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0007 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0007 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0007 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0007 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0007 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0007 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0007 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0007 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0007 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0007 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0007 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0007 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0007 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0007 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0007 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0007 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0007 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0007 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0007 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0007 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0007 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0007 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0007 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0007 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0007 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0007 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0007 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0007 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0007 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0007 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0007 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0007 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0007 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0007 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0007 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0007 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0007 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0007 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0007 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0007 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0007 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0007 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0007 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0007 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0007 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0007 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0007 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0007 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0007 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0007 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0007 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0007 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0007 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0007 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0007 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0007 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0007 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0007 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0007 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0007 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0007 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0007 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0007 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0007 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0007 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0007 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0007 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0007 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0007 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0007 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0007 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0007 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0007 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0007 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0007 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0007 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0007 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0007 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0007 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0007 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0007 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0007 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0007 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0007 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0007 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0007 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0007 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0007 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0007 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0007 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0007 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0007 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0007 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0007 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0007 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0007 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0007 4.7775e-08 0)
L_PG1_12|1 G1_1_TO1 _PG1_12|A1  2.067833848e-12
L_PG1_12|2 _PG1_12|A1 _PG1_12|A2  4.135667696e-12
L_PG1_12|3 _PG1_12|A3 _PG1_12|A4  8.271335392e-12
L_PG1_12|T T09 _PG1_12|T1  2.067833848e-12
L_PG1_12|4 _PG1_12|T1 _PG1_12|T2  4.135667696e-12
L_PG1_12|5 _PG1_12|A4 _PG1_12|Q1  4.135667696e-12
L_PG1_12|6 _PG1_12|Q1 G1_2  2.067833848e-12
IT10|T 0 T10  PWL(0 0 9e-12 0 1.2e-11 0.0014 1.5e-11 0 1.29e-10 0 1.32e-10 0.0014 1.35e-10 0 2.49e-10 0 2.52e-10 0.0014 2.55e-10 0 3.69e-10 0 3.72e-10 0.0014 3.75e-10 0 4.89e-10 0 4.92e-10 0.0014 4.95e-10 0 6.09e-10 0 6.12e-10 0.0014 6.15e-10 0 7.29e-10 0 7.32e-10 0.0014 7.35e-10 0 8.49e-10 0 8.52e-10 0.0014 8.55e-10 0 9.69e-10 0 9.72e-10 0.0014 9.75e-10 0 1.089e-09 0 1.092e-09 0.0014 1.095e-09 0 1.209e-09 0 1.212e-09 0.0014 1.215e-09 0 1.329e-09 0 1.332e-09 0.0014 1.335e-09 0 1.449e-09 0 1.452e-09 0.0014 1.455e-09 0 1.569e-09 0 1.572e-09 0.0014 1.575e-09 0 1.689e-09 0 1.692e-09 0.0014 1.695e-09 0 1.809e-09 0 1.812e-09 0.0014 1.815e-09 0 1.929e-09 0 1.932e-09 0.0014 1.935e-09 0 2.049e-09 0 2.052e-09 0.0014 2.055e-09 0 2.169e-09 0 2.172e-09 0.0014 2.175e-09 0 2.289e-09 0 2.292e-09 0.0014 2.295e-09 0 2.409e-09 0 2.412e-09 0.0014 2.415e-09 0 2.529e-09 0 2.532e-09 0.0014 2.535e-09 0 2.649e-09 0 2.652e-09 0.0014 2.655e-09 0 2.769e-09 0 2.772e-09 0.0014 2.775e-09 0 2.889e-09 0 2.892e-09 0.0014 2.895e-09 0 3.009e-09 0 3.012e-09 0.0014 3.015e-09 0 3.129e-09 0 3.132e-09 0.0014 3.135e-09 0 3.249e-09 0 3.252e-09 0.0014 3.255e-09 0 3.369e-09 0 3.372e-09 0.0014 3.375e-09 0 3.489e-09 0 3.492e-09 0.0014 3.495e-09 0 3.609e-09 0 3.612e-09 0.0014 3.615e-09 0 3.729e-09 0 3.732e-09 0.0014 3.735e-09 0 3.849e-09 0 3.852e-09 0.0014 3.855e-09 0 3.969e-09 0 3.972e-09 0.0014 3.975e-09 0 4.089e-09 0 4.092e-09 0.0014 4.095e-09 0 4.209e-09 0 4.212e-09 0.0014 4.215e-09 0 4.329e-09 0 4.332e-09 0.0014 4.335e-09 0 4.449e-09 0 4.452e-09 0.0014 4.455e-09 0 4.569e-09 0 4.572e-09 0.0014 4.575e-09 0 4.689e-09 0 4.692e-09 0.0014 4.695e-09 0 4.809e-09 0 4.812e-09 0.0014 4.815e-09 0 4.929e-09 0 4.932e-09 0.0014 4.935e-09 0 5.049e-09 0 5.052e-09 0.0014 5.055e-09 0 5.169e-09 0 5.172e-09 0.0014 5.175e-09 0 5.289e-09 0 5.292e-09 0.0014 5.295e-09 0 5.409e-09 0 5.412e-09 0.0014 5.415e-09 0 5.529e-09 0 5.532e-09 0.0014 5.535e-09 0 5.649e-09 0 5.652e-09 0.0014 5.655e-09 0 5.769e-09 0 5.772e-09 0.0014 5.775e-09 0 5.889e-09 0 5.892e-09 0.0014 5.895e-09 0 6.009e-09 0 6.012e-09 0.0014 6.015e-09 0 6.129e-09 0 6.132e-09 0.0014 6.135e-09 0 6.249e-09 0 6.252e-09 0.0014 6.255e-09 0 6.369e-09 0 6.372e-09 0.0014 6.375e-09 0 6.489e-09 0 6.492e-09 0.0014 6.495e-09 0 6.609e-09 0 6.612e-09 0.0014 6.615e-09 0 6.729e-09 0 6.732e-09 0.0014 6.735e-09 0 6.849e-09 0 6.852e-09 0.0014 6.855e-09 0 6.969e-09 0 6.972e-09 0.0014 6.975e-09 0 7.089e-09 0 7.092e-09 0.0014 7.095e-09 0 7.209e-09 0 7.212e-09 0.0014 7.215e-09 0 7.329e-09 0 7.332e-09 0.0014 7.335e-09 0 7.449e-09 0 7.452e-09 0.0014 7.455e-09 0 7.569e-09 0 7.572e-09 0.0014 7.575e-09 0 7.689e-09 0 7.692e-09 0.0014 7.695e-09 0 7.809e-09 0 7.812e-09 0.0014 7.815e-09 0 7.929e-09 0 7.932e-09 0.0014 7.935e-09 0 8.049e-09 0 8.052e-09 0.0014 8.055e-09 0 8.169e-09 0 8.172e-09 0.0014 8.175e-09 0 8.289e-09 0 8.292e-09 0.0014 8.295e-09 0 8.409e-09 0 8.412e-09 0.0014 8.415e-09 0 8.529e-09 0 8.532e-09 0.0014 8.535e-09 0 8.649e-09 0 8.652e-09 0.0014 8.655e-09 0 8.769e-09 0 8.772e-09 0.0014 8.775e-09 0 8.889e-09 0 8.892e-09 0.0014 8.895e-09 0 9.009e-09 0 9.012e-09 0.0014 9.015e-09 0 9.129e-09 0 9.132e-09 0.0014 9.135e-09 0 9.249e-09 0 9.252e-09 0.0014 9.255e-09 0 9.369e-09 0 9.372e-09 0.0014 9.375e-09 0 9.489e-09 0 9.492e-09 0.0014 9.495e-09 0 9.609e-09 0 9.612e-09 0.0014 9.615e-09 0 9.729e-09 0 9.732e-09 0.0014 9.735e-09 0 9.849e-09 0 9.852e-09 0.0014 9.855e-09 0 9.969e-09 0 9.972e-09 0.0014 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0014 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0014 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0014 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0014 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0014 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0014 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0014 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0014 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0014 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0014 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0014 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0014 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0014 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0014 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0014 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0014 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0014 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0014 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0014 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0014 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0014 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0014 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0014 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0014 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0014 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0014 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0014 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0014 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0014 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0014 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0014 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0014 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0014 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0014 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0014 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0014 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0014 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0014 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0014 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0014 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0014 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0014 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0014 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0014 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0014 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0014 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0014 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0014 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0014 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0014 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0014 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0014 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0014 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0014 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0014 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0014 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0014 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0014 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0014 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0014 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0014 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0014 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0014 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0014 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0014 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0014 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0014 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0014 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0014 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0014 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0014 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0014 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0014 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0014 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0014 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0014 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0014 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0014 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0014 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0014 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0014 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0014 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0014 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0014 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0014 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0014 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0014 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0014 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0014 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0014 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0014 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0014 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0014 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0014 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0014 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0014 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0014 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0014 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0014 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0014 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0014 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0014 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0014 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0014 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0014 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0014 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0014 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0014 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0014 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0014 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0014 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0014 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0014 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0014 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0014 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0014 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0014 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0014 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0014 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0014 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0014 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0014 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0014 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0014 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0014 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0014 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0014 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0014 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0014 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0014 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0014 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0014 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0014 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0014 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0014 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0014 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0014 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0014 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0014 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0014 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0014 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0014 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0014 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0014 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0014 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0014 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0014 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0014 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0014 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0014 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0014 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0014 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0014 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0014 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0014 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0014 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0014 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0014 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0014 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0014 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0014 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0014 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0014 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0014 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0014 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0014 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0014 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0014 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0014 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0014 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0014 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0014 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0014 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0014 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0014 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0014 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0014 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0014 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0014 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0014 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0014 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0014 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0014 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0014 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0014 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0014 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0014 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0014 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0014 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0014 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0014 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0014 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0014 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0014 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0014 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0014 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0014 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0014 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0014 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0014 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0014 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0014 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0014 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0014 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0014 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0014 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0014 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0014 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0014 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0014 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0014 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0014 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0014 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0014 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0014 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0014 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0014 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0014 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0014 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0014 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0014 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0014 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0014 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0014 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0014 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0014 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0014 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0014 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0014 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0014 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0014 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0014 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0014 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0014 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0014 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0014 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0014 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0014 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0014 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0014 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0014 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0014 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0014 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0014 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0014 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0014 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0014 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0014 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0014 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0014 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0014 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0014 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0014 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0014 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0014 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0014 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0014 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0014 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0014 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0014 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0014 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0014 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0014 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0014 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0014 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0014 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0014 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0014 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0014 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0014 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0014 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0014 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0014 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0014 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0014 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0014 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0014 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0014 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0014 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0014 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0014 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0014 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0014 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0014 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0014 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0014 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0014 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0014 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0014 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0014 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0014 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0014 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0014 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0014 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0014 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0014 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0014 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0014 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0014 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0014 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0014 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0014 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0014 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0014 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0014 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0014 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0014 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0014 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0014 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0014 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0014 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0014 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0014 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0014 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0014 4.7775e-08 0)
IT11|T 0 T11  PWL(0 0 9e-12 0 1.2e-11 0.0014 1.5e-11 0 1.29e-10 0 1.32e-10 0.0014 1.35e-10 0 2.49e-10 0 2.52e-10 0.0014 2.55e-10 0 3.69e-10 0 3.72e-10 0.0014 3.75e-10 0 4.89e-10 0 4.92e-10 0.0014 4.95e-10 0 6.09e-10 0 6.12e-10 0.0014 6.15e-10 0 7.29e-10 0 7.32e-10 0.0014 7.35e-10 0 8.49e-10 0 8.52e-10 0.0014 8.55e-10 0 9.69e-10 0 9.72e-10 0.0014 9.75e-10 0 1.089e-09 0 1.092e-09 0.0014 1.095e-09 0 1.209e-09 0 1.212e-09 0.0014 1.215e-09 0 1.329e-09 0 1.332e-09 0.0014 1.335e-09 0 1.449e-09 0 1.452e-09 0.0014 1.455e-09 0 1.569e-09 0 1.572e-09 0.0014 1.575e-09 0 1.689e-09 0 1.692e-09 0.0014 1.695e-09 0 1.809e-09 0 1.812e-09 0.0014 1.815e-09 0 1.929e-09 0 1.932e-09 0.0014 1.935e-09 0 2.049e-09 0 2.052e-09 0.0014 2.055e-09 0 2.169e-09 0 2.172e-09 0.0014 2.175e-09 0 2.289e-09 0 2.292e-09 0.0014 2.295e-09 0 2.409e-09 0 2.412e-09 0.0014 2.415e-09 0 2.529e-09 0 2.532e-09 0.0014 2.535e-09 0 2.649e-09 0 2.652e-09 0.0014 2.655e-09 0 2.769e-09 0 2.772e-09 0.0014 2.775e-09 0 2.889e-09 0 2.892e-09 0.0014 2.895e-09 0 3.009e-09 0 3.012e-09 0.0014 3.015e-09 0 3.129e-09 0 3.132e-09 0.0014 3.135e-09 0 3.249e-09 0 3.252e-09 0.0014 3.255e-09 0 3.369e-09 0 3.372e-09 0.0014 3.375e-09 0 3.489e-09 0 3.492e-09 0.0014 3.495e-09 0 3.609e-09 0 3.612e-09 0.0014 3.615e-09 0 3.729e-09 0 3.732e-09 0.0014 3.735e-09 0 3.849e-09 0 3.852e-09 0.0014 3.855e-09 0 3.969e-09 0 3.972e-09 0.0014 3.975e-09 0 4.089e-09 0 4.092e-09 0.0014 4.095e-09 0 4.209e-09 0 4.212e-09 0.0014 4.215e-09 0 4.329e-09 0 4.332e-09 0.0014 4.335e-09 0 4.449e-09 0 4.452e-09 0.0014 4.455e-09 0 4.569e-09 0 4.572e-09 0.0014 4.575e-09 0 4.689e-09 0 4.692e-09 0.0014 4.695e-09 0 4.809e-09 0 4.812e-09 0.0014 4.815e-09 0 4.929e-09 0 4.932e-09 0.0014 4.935e-09 0 5.049e-09 0 5.052e-09 0.0014 5.055e-09 0 5.169e-09 0 5.172e-09 0.0014 5.175e-09 0 5.289e-09 0 5.292e-09 0.0014 5.295e-09 0 5.409e-09 0 5.412e-09 0.0014 5.415e-09 0 5.529e-09 0 5.532e-09 0.0014 5.535e-09 0 5.649e-09 0 5.652e-09 0.0014 5.655e-09 0 5.769e-09 0 5.772e-09 0.0014 5.775e-09 0 5.889e-09 0 5.892e-09 0.0014 5.895e-09 0 6.009e-09 0 6.012e-09 0.0014 6.015e-09 0 6.129e-09 0 6.132e-09 0.0014 6.135e-09 0 6.249e-09 0 6.252e-09 0.0014 6.255e-09 0 6.369e-09 0 6.372e-09 0.0014 6.375e-09 0 6.489e-09 0 6.492e-09 0.0014 6.495e-09 0 6.609e-09 0 6.612e-09 0.0014 6.615e-09 0 6.729e-09 0 6.732e-09 0.0014 6.735e-09 0 6.849e-09 0 6.852e-09 0.0014 6.855e-09 0 6.969e-09 0 6.972e-09 0.0014 6.975e-09 0 7.089e-09 0 7.092e-09 0.0014 7.095e-09 0 7.209e-09 0 7.212e-09 0.0014 7.215e-09 0 7.329e-09 0 7.332e-09 0.0014 7.335e-09 0 7.449e-09 0 7.452e-09 0.0014 7.455e-09 0 7.569e-09 0 7.572e-09 0.0014 7.575e-09 0 7.689e-09 0 7.692e-09 0.0014 7.695e-09 0 7.809e-09 0 7.812e-09 0.0014 7.815e-09 0 7.929e-09 0 7.932e-09 0.0014 7.935e-09 0 8.049e-09 0 8.052e-09 0.0014 8.055e-09 0 8.169e-09 0 8.172e-09 0.0014 8.175e-09 0 8.289e-09 0 8.292e-09 0.0014 8.295e-09 0 8.409e-09 0 8.412e-09 0.0014 8.415e-09 0 8.529e-09 0 8.532e-09 0.0014 8.535e-09 0 8.649e-09 0 8.652e-09 0.0014 8.655e-09 0 8.769e-09 0 8.772e-09 0.0014 8.775e-09 0 8.889e-09 0 8.892e-09 0.0014 8.895e-09 0 9.009e-09 0 9.012e-09 0.0014 9.015e-09 0 9.129e-09 0 9.132e-09 0.0014 9.135e-09 0 9.249e-09 0 9.252e-09 0.0014 9.255e-09 0 9.369e-09 0 9.372e-09 0.0014 9.375e-09 0 9.489e-09 0 9.492e-09 0.0014 9.495e-09 0 9.609e-09 0 9.612e-09 0.0014 9.615e-09 0 9.729e-09 0 9.732e-09 0.0014 9.735e-09 0 9.849e-09 0 9.852e-09 0.0014 9.855e-09 0 9.969e-09 0 9.972e-09 0.0014 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0014 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0014 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0014 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0014 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0014 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0014 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0014 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0014 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0014 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0014 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0014 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0014 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0014 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0014 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0014 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0014 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0014 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0014 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0014 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0014 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0014 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0014 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0014 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0014 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0014 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0014 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0014 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0014 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0014 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0014 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0014 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0014 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0014 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0014 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0014 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0014 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0014 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0014 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0014 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0014 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0014 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0014 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0014 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0014 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0014 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0014 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0014 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0014 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0014 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0014 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0014 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0014 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0014 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0014 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0014 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0014 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0014 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0014 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0014 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0014 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0014 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0014 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0014 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0014 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0014 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0014 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0014 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0014 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0014 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0014 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0014 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0014 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0014 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0014 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0014 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0014 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0014 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0014 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0014 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0014 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0014 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0014 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0014 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0014 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0014 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0014 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0014 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0014 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0014 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0014 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0014 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0014 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0014 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0014 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0014 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0014 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0014 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0014 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0014 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0014 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0014 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0014 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0014 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0014 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0014 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0014 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0014 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0014 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0014 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0014 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0014 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0014 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0014 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0014 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0014 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0014 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0014 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0014 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0014 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0014 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0014 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0014 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0014 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0014 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0014 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0014 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0014 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0014 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0014 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0014 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0014 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0014 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0014 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0014 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0014 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0014 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0014 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0014 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0014 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0014 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0014 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0014 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0014 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0014 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0014 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0014 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0014 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0014 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0014 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0014 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0014 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0014 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0014 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0014 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0014 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0014 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0014 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0014 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0014 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0014 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0014 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0014 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0014 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0014 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0014 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0014 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0014 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0014 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0014 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0014 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0014 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0014 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0014 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0014 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0014 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0014 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0014 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0014 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0014 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0014 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0014 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0014 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0014 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0014 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0014 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0014 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0014 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0014 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0014 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0014 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0014 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0014 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0014 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0014 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0014 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0014 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0014 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0014 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0014 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0014 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0014 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0014 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0014 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0014 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0014 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0014 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0014 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0014 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0014 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0014 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0014 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0014 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0014 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0014 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0014 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0014 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0014 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0014 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0014 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0014 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0014 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0014 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0014 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0014 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0014 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0014 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0014 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0014 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0014 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0014 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0014 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0014 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0014 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0014 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0014 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0014 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0014 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0014 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0014 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0014 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0014 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0014 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0014 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0014 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0014 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0014 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0014 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0014 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0014 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0014 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0014 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0014 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0014 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0014 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0014 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0014 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0014 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0014 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0014 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0014 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0014 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0014 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0014 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0014 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0014 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0014 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0014 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0014 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0014 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0014 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0014 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0014 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0014 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0014 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0014 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0014 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0014 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0014 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0014 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0014 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0014 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0014 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0014 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0014 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0014 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0014 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0014 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0014 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0014 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0014 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0014 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0014 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0014 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0014 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0014 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0014 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0014 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0014 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0014 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0014 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0014 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0014 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0014 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0014 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0014 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0014 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0014 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0014 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0014 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0014 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0014 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0014 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0014 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0014 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0014 4.7775e-08 0)
ID11|T 0 D11  PWL(0 0 9e-12 0 1.2e-11 0.0007 1.5e-11 0 1.29e-10 0 1.32e-10 0.0007 1.35e-10 0 2.49e-10 0 2.52e-10 0.0007 2.55e-10 0 3.69e-10 0 3.72e-10 0.0007 3.75e-10 0 4.89e-10 0 4.92e-10 0.0007 4.95e-10 0 6.09e-10 0 6.12e-10 0.0007 6.15e-10 0 7.29e-10 0 7.32e-10 0.0007 7.35e-10 0 8.49e-10 0 8.52e-10 0.0007 8.55e-10 0 9.69e-10 0 9.72e-10 0.0007 9.75e-10 0 1.089e-09 0 1.092e-09 0.0007 1.095e-09 0 1.209e-09 0 1.212e-09 0.0007 1.215e-09 0 1.329e-09 0 1.332e-09 0.0007 1.335e-09 0 1.449e-09 0 1.452e-09 0.0007 1.455e-09 0 1.569e-09 0 1.572e-09 0.0007 1.575e-09 0 1.689e-09 0 1.692e-09 0.0007 1.695e-09 0 1.809e-09 0 1.812e-09 0.0007 1.815e-09 0 1.929e-09 0 1.932e-09 0.0007 1.935e-09 0 2.049e-09 0 2.052e-09 0.0007 2.055e-09 0 2.169e-09 0 2.172e-09 0.0007 2.175e-09 0 2.289e-09 0 2.292e-09 0.0007 2.295e-09 0 2.409e-09 0 2.412e-09 0.0007 2.415e-09 0 2.529e-09 0 2.532e-09 0.0007 2.535e-09 0 2.649e-09 0 2.652e-09 0.0007 2.655e-09 0 2.769e-09 0 2.772e-09 0.0007 2.775e-09 0 2.889e-09 0 2.892e-09 0.0007 2.895e-09 0 3.009e-09 0 3.012e-09 0.0007 3.015e-09 0 3.129e-09 0 3.132e-09 0.0007 3.135e-09 0 3.249e-09 0 3.252e-09 0.0007 3.255e-09 0 3.369e-09 0 3.372e-09 0.0007 3.375e-09 0 3.489e-09 0 3.492e-09 0.0007 3.495e-09 0 3.609e-09 0 3.612e-09 0.0007 3.615e-09 0 3.729e-09 0 3.732e-09 0.0007 3.735e-09 0 3.849e-09 0 3.852e-09 0.0007 3.855e-09 0 3.969e-09 0 3.972e-09 0.0007 3.975e-09 0 4.089e-09 0 4.092e-09 0.0007 4.095e-09 0 4.209e-09 0 4.212e-09 0.0007 4.215e-09 0 4.329e-09 0 4.332e-09 0.0007 4.335e-09 0 4.449e-09 0 4.452e-09 0.0007 4.455e-09 0 4.569e-09 0 4.572e-09 0.0007 4.575e-09 0 4.689e-09 0 4.692e-09 0.0007 4.695e-09 0 4.809e-09 0 4.812e-09 0.0007 4.815e-09 0 4.929e-09 0 4.932e-09 0.0007 4.935e-09 0 5.049e-09 0 5.052e-09 0.0007 5.055e-09 0 5.169e-09 0 5.172e-09 0.0007 5.175e-09 0 5.289e-09 0 5.292e-09 0.0007 5.295e-09 0 5.409e-09 0 5.412e-09 0.0007 5.415e-09 0 5.529e-09 0 5.532e-09 0.0007 5.535e-09 0 5.649e-09 0 5.652e-09 0.0007 5.655e-09 0 5.769e-09 0 5.772e-09 0.0007 5.775e-09 0 5.889e-09 0 5.892e-09 0.0007 5.895e-09 0 6.009e-09 0 6.012e-09 0.0007 6.015e-09 0 6.129e-09 0 6.132e-09 0.0007 6.135e-09 0 6.249e-09 0 6.252e-09 0.0007 6.255e-09 0 6.369e-09 0 6.372e-09 0.0007 6.375e-09 0 6.489e-09 0 6.492e-09 0.0007 6.495e-09 0 6.609e-09 0 6.612e-09 0.0007 6.615e-09 0 6.729e-09 0 6.732e-09 0.0007 6.735e-09 0 6.849e-09 0 6.852e-09 0.0007 6.855e-09 0 6.969e-09 0 6.972e-09 0.0007 6.975e-09 0 7.089e-09 0 7.092e-09 0.0007 7.095e-09 0 7.209e-09 0 7.212e-09 0.0007 7.215e-09 0 7.329e-09 0 7.332e-09 0.0007 7.335e-09 0 7.449e-09 0 7.452e-09 0.0007 7.455e-09 0 7.569e-09 0 7.572e-09 0.0007 7.575e-09 0 7.689e-09 0 7.692e-09 0.0007 7.695e-09 0 7.809e-09 0 7.812e-09 0.0007 7.815e-09 0 7.929e-09 0 7.932e-09 0.0007 7.935e-09 0 8.049e-09 0 8.052e-09 0.0007 8.055e-09 0 8.169e-09 0 8.172e-09 0.0007 8.175e-09 0 8.289e-09 0 8.292e-09 0.0007 8.295e-09 0 8.409e-09 0 8.412e-09 0.0007 8.415e-09 0 8.529e-09 0 8.532e-09 0.0007 8.535e-09 0 8.649e-09 0 8.652e-09 0.0007 8.655e-09 0 8.769e-09 0 8.772e-09 0.0007 8.775e-09 0 8.889e-09 0 8.892e-09 0.0007 8.895e-09 0 9.009e-09 0 9.012e-09 0.0007 9.015e-09 0 9.129e-09 0 9.132e-09 0.0007 9.135e-09 0 9.249e-09 0 9.252e-09 0.0007 9.255e-09 0 9.369e-09 0 9.372e-09 0.0007 9.375e-09 0 9.489e-09 0 9.492e-09 0.0007 9.495e-09 0 9.609e-09 0 9.612e-09 0.0007 9.615e-09 0 9.729e-09 0 9.732e-09 0.0007 9.735e-09 0 9.849e-09 0 9.852e-09 0.0007 9.855e-09 0 9.969e-09 0 9.972e-09 0.0007 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0007 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0007 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0007 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0007 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0007 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0007 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0007 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0007 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0007 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0007 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0007 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0007 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0007 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0007 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0007 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0007 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0007 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0007 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0007 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0007 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0007 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0007 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0007 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0007 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0007 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0007 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0007 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0007 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0007 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0007 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0007 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0007 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0007 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0007 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0007 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0007 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0007 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0007 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0007 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0007 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0007 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0007 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0007 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0007 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0007 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0007 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0007 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0007 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0007 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0007 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0007 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0007 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0007 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0007 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0007 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0007 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0007 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0007 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0007 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0007 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0007 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0007 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0007 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0007 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0007 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0007 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0007 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0007 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0007 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0007 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0007 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0007 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0007 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0007 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0007 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0007 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0007 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0007 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0007 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0007 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0007 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0007 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0007 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0007 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0007 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0007 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0007 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0007 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0007 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0007 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0007 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0007 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0007 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0007 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0007 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0007 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0007 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0007 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0007 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0007 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0007 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0007 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0007 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0007 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0007 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0007 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0007 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0007 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0007 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0007 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0007 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0007 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0007 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0007 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0007 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0007 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0007 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0007 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0007 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0007 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0007 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0007 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0007 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0007 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0007 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0007 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0007 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0007 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0007 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0007 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0007 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0007 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0007 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0007 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0007 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0007 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0007 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0007 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0007 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0007 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0007 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0007 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0007 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0007 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0007 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0007 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0007 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0007 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0007 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0007 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0007 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0007 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0007 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0007 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0007 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0007 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0007 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0007 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0007 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0007 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0007 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0007 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0007 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0007 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0007 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0007 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0007 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0007 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0007 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0007 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0007 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0007 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0007 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0007 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0007 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0007 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0007 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0007 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0007 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0007 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0007 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0007 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0007 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0007 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0007 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0007 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0007 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0007 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0007 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0007 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0007 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0007 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0007 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0007 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0007 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0007 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0007 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0007 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0007 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0007 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0007 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0007 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0007 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0007 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0007 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0007 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0007 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0007 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0007 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0007 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0007 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0007 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0007 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0007 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0007 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0007 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0007 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0007 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0007 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0007 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0007 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0007 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0007 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0007 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0007 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0007 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0007 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0007 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0007 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0007 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0007 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0007 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0007 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0007 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0007 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0007 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0007 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0007 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0007 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0007 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0007 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0007 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0007 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0007 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0007 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0007 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0007 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0007 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0007 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0007 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0007 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0007 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0007 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0007 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0007 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0007 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0007 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0007 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0007 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0007 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0007 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0007 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0007 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0007 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0007 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0007 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0007 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0007 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0007 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0007 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0007 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0007 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0007 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0007 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0007 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0007 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0007 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0007 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0007 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0007 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0007 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0007 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0007 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0007 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0007 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0007 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0007 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0007 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0007 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0007 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0007 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0007 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0007 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0007 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0007 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0007 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0007 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0007 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0007 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0007 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0007 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0007 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0007 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0007 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0007 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0007 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0007 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0007 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0007 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0007 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0007 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0007 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0007 4.7775e-08 0)
L_DFF_IP1_12|1 IP1_1_OUT_RX _DFF_IP1_12|A1  2.067833848e-12
L_DFF_IP1_12|2 _DFF_IP1_12|A1 _DFF_IP1_12|A2  4.135667696e-12
L_DFF_IP1_12|3 _DFF_IP1_12|A3 _DFF_IP1_12|A4  8.271335392e-12
L_DFF_IP1_12|T D11 _DFF_IP1_12|T1  2.067833848e-12
L_DFF_IP1_12|4 _DFF_IP1_12|T1 _DFF_IP1_12|T2  4.135667696e-12
L_DFF_IP1_12|5 _DFF_IP1_12|A4 _DFF_IP1_12|Q1  4.135667696e-12
L_DFF_IP1_12|6 _DFF_IP1_12|Q1 IP1_2_OUT  2.067833848e-12
ID12|T 0 D12  PWL(0 0 9e-12 0 1.2e-11 0.0007 1.5e-11 0 1.29e-10 0 1.32e-10 0.0007 1.35e-10 0 2.49e-10 0 2.52e-10 0.0007 2.55e-10 0 3.69e-10 0 3.72e-10 0.0007 3.75e-10 0 4.89e-10 0 4.92e-10 0.0007 4.95e-10 0 6.09e-10 0 6.12e-10 0.0007 6.15e-10 0 7.29e-10 0 7.32e-10 0.0007 7.35e-10 0 8.49e-10 0 8.52e-10 0.0007 8.55e-10 0 9.69e-10 0 9.72e-10 0.0007 9.75e-10 0 1.089e-09 0 1.092e-09 0.0007 1.095e-09 0 1.209e-09 0 1.212e-09 0.0007 1.215e-09 0 1.329e-09 0 1.332e-09 0.0007 1.335e-09 0 1.449e-09 0 1.452e-09 0.0007 1.455e-09 0 1.569e-09 0 1.572e-09 0.0007 1.575e-09 0 1.689e-09 0 1.692e-09 0.0007 1.695e-09 0 1.809e-09 0 1.812e-09 0.0007 1.815e-09 0 1.929e-09 0 1.932e-09 0.0007 1.935e-09 0 2.049e-09 0 2.052e-09 0.0007 2.055e-09 0 2.169e-09 0 2.172e-09 0.0007 2.175e-09 0 2.289e-09 0 2.292e-09 0.0007 2.295e-09 0 2.409e-09 0 2.412e-09 0.0007 2.415e-09 0 2.529e-09 0 2.532e-09 0.0007 2.535e-09 0 2.649e-09 0 2.652e-09 0.0007 2.655e-09 0 2.769e-09 0 2.772e-09 0.0007 2.775e-09 0 2.889e-09 0 2.892e-09 0.0007 2.895e-09 0 3.009e-09 0 3.012e-09 0.0007 3.015e-09 0 3.129e-09 0 3.132e-09 0.0007 3.135e-09 0 3.249e-09 0 3.252e-09 0.0007 3.255e-09 0 3.369e-09 0 3.372e-09 0.0007 3.375e-09 0 3.489e-09 0 3.492e-09 0.0007 3.495e-09 0 3.609e-09 0 3.612e-09 0.0007 3.615e-09 0 3.729e-09 0 3.732e-09 0.0007 3.735e-09 0 3.849e-09 0 3.852e-09 0.0007 3.855e-09 0 3.969e-09 0 3.972e-09 0.0007 3.975e-09 0 4.089e-09 0 4.092e-09 0.0007 4.095e-09 0 4.209e-09 0 4.212e-09 0.0007 4.215e-09 0 4.329e-09 0 4.332e-09 0.0007 4.335e-09 0 4.449e-09 0 4.452e-09 0.0007 4.455e-09 0 4.569e-09 0 4.572e-09 0.0007 4.575e-09 0 4.689e-09 0 4.692e-09 0.0007 4.695e-09 0 4.809e-09 0 4.812e-09 0.0007 4.815e-09 0 4.929e-09 0 4.932e-09 0.0007 4.935e-09 0 5.049e-09 0 5.052e-09 0.0007 5.055e-09 0 5.169e-09 0 5.172e-09 0.0007 5.175e-09 0 5.289e-09 0 5.292e-09 0.0007 5.295e-09 0 5.409e-09 0 5.412e-09 0.0007 5.415e-09 0 5.529e-09 0 5.532e-09 0.0007 5.535e-09 0 5.649e-09 0 5.652e-09 0.0007 5.655e-09 0 5.769e-09 0 5.772e-09 0.0007 5.775e-09 0 5.889e-09 0 5.892e-09 0.0007 5.895e-09 0 6.009e-09 0 6.012e-09 0.0007 6.015e-09 0 6.129e-09 0 6.132e-09 0.0007 6.135e-09 0 6.249e-09 0 6.252e-09 0.0007 6.255e-09 0 6.369e-09 0 6.372e-09 0.0007 6.375e-09 0 6.489e-09 0 6.492e-09 0.0007 6.495e-09 0 6.609e-09 0 6.612e-09 0.0007 6.615e-09 0 6.729e-09 0 6.732e-09 0.0007 6.735e-09 0 6.849e-09 0 6.852e-09 0.0007 6.855e-09 0 6.969e-09 0 6.972e-09 0.0007 6.975e-09 0 7.089e-09 0 7.092e-09 0.0007 7.095e-09 0 7.209e-09 0 7.212e-09 0.0007 7.215e-09 0 7.329e-09 0 7.332e-09 0.0007 7.335e-09 0 7.449e-09 0 7.452e-09 0.0007 7.455e-09 0 7.569e-09 0 7.572e-09 0.0007 7.575e-09 0 7.689e-09 0 7.692e-09 0.0007 7.695e-09 0 7.809e-09 0 7.812e-09 0.0007 7.815e-09 0 7.929e-09 0 7.932e-09 0.0007 7.935e-09 0 8.049e-09 0 8.052e-09 0.0007 8.055e-09 0 8.169e-09 0 8.172e-09 0.0007 8.175e-09 0 8.289e-09 0 8.292e-09 0.0007 8.295e-09 0 8.409e-09 0 8.412e-09 0.0007 8.415e-09 0 8.529e-09 0 8.532e-09 0.0007 8.535e-09 0 8.649e-09 0 8.652e-09 0.0007 8.655e-09 0 8.769e-09 0 8.772e-09 0.0007 8.775e-09 0 8.889e-09 0 8.892e-09 0.0007 8.895e-09 0 9.009e-09 0 9.012e-09 0.0007 9.015e-09 0 9.129e-09 0 9.132e-09 0.0007 9.135e-09 0 9.249e-09 0 9.252e-09 0.0007 9.255e-09 0 9.369e-09 0 9.372e-09 0.0007 9.375e-09 0 9.489e-09 0 9.492e-09 0.0007 9.495e-09 0 9.609e-09 0 9.612e-09 0.0007 9.615e-09 0 9.729e-09 0 9.732e-09 0.0007 9.735e-09 0 9.849e-09 0 9.852e-09 0.0007 9.855e-09 0 9.969e-09 0 9.972e-09 0.0007 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0007 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0007 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0007 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0007 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0007 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0007 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0007 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0007 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0007 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0007 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0007 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0007 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0007 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0007 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0007 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0007 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0007 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0007 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0007 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0007 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0007 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0007 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0007 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0007 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0007 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0007 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0007 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0007 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0007 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0007 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0007 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0007 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0007 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0007 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0007 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0007 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0007 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0007 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0007 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0007 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0007 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0007 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0007 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0007 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0007 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0007 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0007 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0007 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0007 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0007 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0007 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0007 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0007 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0007 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0007 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0007 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0007 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0007 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0007 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0007 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0007 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0007 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0007 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0007 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0007 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0007 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0007 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0007 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0007 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0007 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0007 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0007 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0007 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0007 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0007 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0007 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0007 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0007 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0007 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0007 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0007 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0007 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0007 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0007 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0007 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0007 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0007 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0007 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0007 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0007 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0007 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0007 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0007 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0007 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0007 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0007 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0007 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0007 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0007 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0007 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0007 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0007 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0007 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0007 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0007 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0007 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0007 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0007 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0007 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0007 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0007 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0007 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0007 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0007 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0007 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0007 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0007 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0007 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0007 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0007 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0007 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0007 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0007 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0007 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0007 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0007 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0007 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0007 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0007 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0007 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0007 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0007 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0007 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0007 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0007 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0007 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0007 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0007 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0007 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0007 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0007 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0007 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0007 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0007 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0007 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0007 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0007 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0007 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0007 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0007 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0007 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0007 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0007 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0007 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0007 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0007 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0007 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0007 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0007 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0007 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0007 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0007 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0007 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0007 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0007 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0007 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0007 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0007 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0007 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0007 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0007 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0007 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0007 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0007 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0007 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0007 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0007 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0007 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0007 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0007 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0007 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0007 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0007 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0007 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0007 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0007 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0007 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0007 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0007 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0007 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0007 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0007 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0007 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0007 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0007 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0007 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0007 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0007 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0007 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0007 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0007 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0007 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0007 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0007 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0007 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0007 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0007 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0007 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0007 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0007 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0007 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0007 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0007 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0007 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0007 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0007 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0007 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0007 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0007 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0007 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0007 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0007 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0007 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0007 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0007 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0007 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0007 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0007 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0007 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0007 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0007 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0007 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0007 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0007 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0007 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0007 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0007 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0007 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0007 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0007 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0007 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0007 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0007 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0007 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0007 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0007 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0007 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0007 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0007 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0007 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0007 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0007 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0007 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0007 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0007 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0007 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0007 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0007 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0007 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0007 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0007 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0007 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0007 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0007 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0007 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0007 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0007 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0007 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0007 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0007 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0007 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0007 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0007 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0007 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0007 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0007 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0007 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0007 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0007 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0007 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0007 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0007 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0007 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0007 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0007 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0007 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0007 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0007 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0007 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0007 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0007 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0007 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0007 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0007 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0007 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0007 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0007 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0007 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0007 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0007 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0007 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0007 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0007 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0007 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0007 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0007 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0007 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0007 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0007 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0007 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0007 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0007 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0007 4.7775e-08 0)
L_DFF_IP2_12|1 IP2_1_OUT_RX _DFF_IP2_12|A1  2.067833848e-12
L_DFF_IP2_12|2 _DFF_IP2_12|A1 _DFF_IP2_12|A2  4.135667696e-12
L_DFF_IP2_12|3 _DFF_IP2_12|A3 _DFF_IP2_12|A4  8.271335392e-12
L_DFF_IP2_12|T D12 _DFF_IP2_12|T1  2.067833848e-12
L_DFF_IP2_12|4 _DFF_IP2_12|T1 _DFF_IP2_12|T2  4.135667696e-12
L_DFF_IP2_12|5 _DFF_IP2_12|A4 _DFF_IP2_12|Q1  4.135667696e-12
L_DFF_IP2_12|6 _DFF_IP2_12|Q1 IP2_2_OUT  2.067833848e-12
ID13|T 0 D13  PWL(0 0 9e-12 0 1.2e-11 0.0007 1.5e-11 0 1.29e-10 0 1.32e-10 0.0007 1.35e-10 0 2.49e-10 0 2.52e-10 0.0007 2.55e-10 0 3.69e-10 0 3.72e-10 0.0007 3.75e-10 0 4.89e-10 0 4.92e-10 0.0007 4.95e-10 0 6.09e-10 0 6.12e-10 0.0007 6.15e-10 0 7.29e-10 0 7.32e-10 0.0007 7.35e-10 0 8.49e-10 0 8.52e-10 0.0007 8.55e-10 0 9.69e-10 0 9.72e-10 0.0007 9.75e-10 0 1.089e-09 0 1.092e-09 0.0007 1.095e-09 0 1.209e-09 0 1.212e-09 0.0007 1.215e-09 0 1.329e-09 0 1.332e-09 0.0007 1.335e-09 0 1.449e-09 0 1.452e-09 0.0007 1.455e-09 0 1.569e-09 0 1.572e-09 0.0007 1.575e-09 0 1.689e-09 0 1.692e-09 0.0007 1.695e-09 0 1.809e-09 0 1.812e-09 0.0007 1.815e-09 0 1.929e-09 0 1.932e-09 0.0007 1.935e-09 0 2.049e-09 0 2.052e-09 0.0007 2.055e-09 0 2.169e-09 0 2.172e-09 0.0007 2.175e-09 0 2.289e-09 0 2.292e-09 0.0007 2.295e-09 0 2.409e-09 0 2.412e-09 0.0007 2.415e-09 0 2.529e-09 0 2.532e-09 0.0007 2.535e-09 0 2.649e-09 0 2.652e-09 0.0007 2.655e-09 0 2.769e-09 0 2.772e-09 0.0007 2.775e-09 0 2.889e-09 0 2.892e-09 0.0007 2.895e-09 0 3.009e-09 0 3.012e-09 0.0007 3.015e-09 0 3.129e-09 0 3.132e-09 0.0007 3.135e-09 0 3.249e-09 0 3.252e-09 0.0007 3.255e-09 0 3.369e-09 0 3.372e-09 0.0007 3.375e-09 0 3.489e-09 0 3.492e-09 0.0007 3.495e-09 0 3.609e-09 0 3.612e-09 0.0007 3.615e-09 0 3.729e-09 0 3.732e-09 0.0007 3.735e-09 0 3.849e-09 0 3.852e-09 0.0007 3.855e-09 0 3.969e-09 0 3.972e-09 0.0007 3.975e-09 0 4.089e-09 0 4.092e-09 0.0007 4.095e-09 0 4.209e-09 0 4.212e-09 0.0007 4.215e-09 0 4.329e-09 0 4.332e-09 0.0007 4.335e-09 0 4.449e-09 0 4.452e-09 0.0007 4.455e-09 0 4.569e-09 0 4.572e-09 0.0007 4.575e-09 0 4.689e-09 0 4.692e-09 0.0007 4.695e-09 0 4.809e-09 0 4.812e-09 0.0007 4.815e-09 0 4.929e-09 0 4.932e-09 0.0007 4.935e-09 0 5.049e-09 0 5.052e-09 0.0007 5.055e-09 0 5.169e-09 0 5.172e-09 0.0007 5.175e-09 0 5.289e-09 0 5.292e-09 0.0007 5.295e-09 0 5.409e-09 0 5.412e-09 0.0007 5.415e-09 0 5.529e-09 0 5.532e-09 0.0007 5.535e-09 0 5.649e-09 0 5.652e-09 0.0007 5.655e-09 0 5.769e-09 0 5.772e-09 0.0007 5.775e-09 0 5.889e-09 0 5.892e-09 0.0007 5.895e-09 0 6.009e-09 0 6.012e-09 0.0007 6.015e-09 0 6.129e-09 0 6.132e-09 0.0007 6.135e-09 0 6.249e-09 0 6.252e-09 0.0007 6.255e-09 0 6.369e-09 0 6.372e-09 0.0007 6.375e-09 0 6.489e-09 0 6.492e-09 0.0007 6.495e-09 0 6.609e-09 0 6.612e-09 0.0007 6.615e-09 0 6.729e-09 0 6.732e-09 0.0007 6.735e-09 0 6.849e-09 0 6.852e-09 0.0007 6.855e-09 0 6.969e-09 0 6.972e-09 0.0007 6.975e-09 0 7.089e-09 0 7.092e-09 0.0007 7.095e-09 0 7.209e-09 0 7.212e-09 0.0007 7.215e-09 0 7.329e-09 0 7.332e-09 0.0007 7.335e-09 0 7.449e-09 0 7.452e-09 0.0007 7.455e-09 0 7.569e-09 0 7.572e-09 0.0007 7.575e-09 0 7.689e-09 0 7.692e-09 0.0007 7.695e-09 0 7.809e-09 0 7.812e-09 0.0007 7.815e-09 0 7.929e-09 0 7.932e-09 0.0007 7.935e-09 0 8.049e-09 0 8.052e-09 0.0007 8.055e-09 0 8.169e-09 0 8.172e-09 0.0007 8.175e-09 0 8.289e-09 0 8.292e-09 0.0007 8.295e-09 0 8.409e-09 0 8.412e-09 0.0007 8.415e-09 0 8.529e-09 0 8.532e-09 0.0007 8.535e-09 0 8.649e-09 0 8.652e-09 0.0007 8.655e-09 0 8.769e-09 0 8.772e-09 0.0007 8.775e-09 0 8.889e-09 0 8.892e-09 0.0007 8.895e-09 0 9.009e-09 0 9.012e-09 0.0007 9.015e-09 0 9.129e-09 0 9.132e-09 0.0007 9.135e-09 0 9.249e-09 0 9.252e-09 0.0007 9.255e-09 0 9.369e-09 0 9.372e-09 0.0007 9.375e-09 0 9.489e-09 0 9.492e-09 0.0007 9.495e-09 0 9.609e-09 0 9.612e-09 0.0007 9.615e-09 0 9.729e-09 0 9.732e-09 0.0007 9.735e-09 0 9.849e-09 0 9.852e-09 0.0007 9.855e-09 0 9.969e-09 0 9.972e-09 0.0007 9.975e-09 0 1.0089e-08 0 1.0092e-08 0.0007 1.0095e-08 0 1.0209e-08 0 1.0212e-08 0.0007 1.0215e-08 0 1.0329e-08 0 1.0332e-08 0.0007 1.0335e-08 0 1.0449e-08 0 1.0452e-08 0.0007 1.0455e-08 0 1.0569e-08 0 1.0572e-08 0.0007 1.0575e-08 0 1.0689e-08 0 1.0692e-08 0.0007 1.0695e-08 0 1.0809e-08 0 1.0812e-08 0.0007 1.0815e-08 0 1.0929e-08 0 1.0932e-08 0.0007 1.0935e-08 0 1.1049e-08 0 1.1052e-08 0.0007 1.1055e-08 0 1.1169e-08 0 1.1172e-08 0.0007 1.1175e-08 0 1.1289e-08 0 1.1292e-08 0.0007 1.1295e-08 0 1.1409e-08 0 1.1412e-08 0.0007 1.1415e-08 0 1.1529e-08 0 1.1532e-08 0.0007 1.1535e-08 0 1.1649e-08 0 1.1652e-08 0.0007 1.1655e-08 0 1.1769e-08 0 1.1772e-08 0.0007 1.1775e-08 0 1.1889e-08 0 1.1892e-08 0.0007 1.1895e-08 0 1.2009e-08 0 1.2012e-08 0.0007 1.2015e-08 0 1.2129e-08 0 1.2132e-08 0.0007 1.2135e-08 0 1.2249e-08 0 1.2252e-08 0.0007 1.2255e-08 0 1.2369e-08 0 1.2372e-08 0.0007 1.2375e-08 0 1.2489e-08 0 1.2492e-08 0.0007 1.2495e-08 0 1.2609e-08 0 1.2612e-08 0.0007 1.2615e-08 0 1.2729e-08 0 1.2732e-08 0.0007 1.2735e-08 0 1.2849e-08 0 1.2852e-08 0.0007 1.2855e-08 0 1.2969e-08 0 1.2972e-08 0.0007 1.2975e-08 0 1.3089e-08 0 1.3092e-08 0.0007 1.3095e-08 0 1.3209e-08 0 1.3212e-08 0.0007 1.3215e-08 0 1.3329e-08 0 1.3332e-08 0.0007 1.3335e-08 0 1.3449e-08 0 1.3452e-08 0.0007 1.3455e-08 0 1.3569e-08 0 1.3572e-08 0.0007 1.3575e-08 0 1.3689e-08 0 1.3692e-08 0.0007 1.3695e-08 0 1.3809e-08 0 1.3812e-08 0.0007 1.3815e-08 0 1.3929e-08 0 1.3932e-08 0.0007 1.3935e-08 0 1.4049e-08 0 1.4052e-08 0.0007 1.4055e-08 0 1.4169e-08 0 1.4172e-08 0.0007 1.4175e-08 0 1.4289e-08 0 1.4292e-08 0.0007 1.4295e-08 0 1.4409e-08 0 1.4412e-08 0.0007 1.4415e-08 0 1.4529e-08 0 1.4532e-08 0.0007 1.4535e-08 0 1.4649e-08 0 1.4652e-08 0.0007 1.4655e-08 0 1.4769e-08 0 1.4772e-08 0.0007 1.4775e-08 0 1.4889e-08 0 1.4892e-08 0.0007 1.4895e-08 0 1.5009e-08 0 1.5012e-08 0.0007 1.5015e-08 0 1.5129e-08 0 1.5132e-08 0.0007 1.5135e-08 0 1.5249e-08 0 1.5252e-08 0.0007 1.5255e-08 0 1.5369e-08 0 1.5372e-08 0.0007 1.5375e-08 0 1.5489e-08 0 1.5492e-08 0.0007 1.5495e-08 0 1.5609e-08 0 1.5612e-08 0.0007 1.5615e-08 0 1.5729e-08 0 1.5732e-08 0.0007 1.5735e-08 0 1.5849e-08 0 1.5852e-08 0.0007 1.5855e-08 0 1.5969e-08 0 1.5972e-08 0.0007 1.5975e-08 0 1.6089e-08 0 1.6092e-08 0.0007 1.6095e-08 0 1.6209e-08 0 1.6212e-08 0.0007 1.6215e-08 0 1.6329e-08 0 1.6332e-08 0.0007 1.6335e-08 0 1.6449e-08 0 1.6452e-08 0.0007 1.6455e-08 0 1.6569e-08 0 1.6572e-08 0.0007 1.6575e-08 0 1.6689e-08 0 1.6692e-08 0.0007 1.6695e-08 0 1.6809e-08 0 1.6812e-08 0.0007 1.6815e-08 0 1.6929e-08 0 1.6932e-08 0.0007 1.6935e-08 0 1.7049e-08 0 1.7052e-08 0.0007 1.7055e-08 0 1.7169e-08 0 1.7172e-08 0.0007 1.7175e-08 0 1.7289e-08 0 1.7292e-08 0.0007 1.7295e-08 0 1.7409e-08 0 1.7412e-08 0.0007 1.7415e-08 0 1.7529e-08 0 1.7532e-08 0.0007 1.7535e-08 0 1.7649e-08 0 1.7652e-08 0.0007 1.7655e-08 0 1.7769e-08 0 1.7772e-08 0.0007 1.7775e-08 0 1.7889e-08 0 1.7892e-08 0.0007 1.7895e-08 0 1.8009e-08 0 1.8012e-08 0.0007 1.8015e-08 0 1.8129e-08 0 1.8132e-08 0.0007 1.8135e-08 0 1.8249e-08 0 1.8252e-08 0.0007 1.8255e-08 0 1.8369e-08 0 1.8372e-08 0.0007 1.8375e-08 0 1.8489e-08 0 1.8492e-08 0.0007 1.8495e-08 0 1.8609e-08 0 1.8612e-08 0.0007 1.8615e-08 0 1.8729e-08 0 1.8732e-08 0.0007 1.8735e-08 0 1.8849e-08 0 1.8852e-08 0.0007 1.8855e-08 0 1.8969e-08 0 1.8972e-08 0.0007 1.8975e-08 0 1.9089e-08 0 1.9092e-08 0.0007 1.9095e-08 0 1.9209e-08 0 1.9212e-08 0.0007 1.9215e-08 0 1.9329e-08 0 1.9332e-08 0.0007 1.9335e-08 0 1.9449e-08 0 1.9452e-08 0.0007 1.9455e-08 0 1.9569e-08 0 1.9572e-08 0.0007 1.9575e-08 0 1.9689e-08 0 1.9692e-08 0.0007 1.9695e-08 0 1.9809e-08 0 1.9812e-08 0.0007 1.9815e-08 0 1.9929e-08 0 1.9932e-08 0.0007 1.9935e-08 0 2.0049e-08 0 2.0052e-08 0.0007 2.0055e-08 0 2.0169e-08 0 2.0172e-08 0.0007 2.0175e-08 0 2.0289e-08 0 2.0292e-08 0.0007 2.0295e-08 0 2.0409e-08 0 2.0412e-08 0.0007 2.0415e-08 0 2.0529e-08 0 2.0532e-08 0.0007 2.0535e-08 0 2.0649e-08 0 2.0652e-08 0.0007 2.0655e-08 0 2.0769e-08 0 2.0772e-08 0.0007 2.0775e-08 0 2.0889e-08 0 2.0892e-08 0.0007 2.0895e-08 0 2.1009e-08 0 2.1012e-08 0.0007 2.1015e-08 0 2.1129e-08 0 2.1132e-08 0.0007 2.1135e-08 0 2.1249e-08 0 2.1252e-08 0.0007 2.1255e-08 0 2.1369e-08 0 2.1372e-08 0.0007 2.1375e-08 0 2.1489e-08 0 2.1492e-08 0.0007 2.1495e-08 0 2.1609e-08 0 2.1612e-08 0.0007 2.1615e-08 0 2.1729e-08 0 2.1732e-08 0.0007 2.1735e-08 0 2.1849e-08 0 2.1852e-08 0.0007 2.1855e-08 0 2.1969e-08 0 2.1972e-08 0.0007 2.1975e-08 0 2.2089e-08 0 2.2092e-08 0.0007 2.2095e-08 0 2.2209e-08 0 2.2212e-08 0.0007 2.2215e-08 0 2.2329e-08 0 2.2332e-08 0.0007 2.2335e-08 0 2.2449e-08 0 2.2452e-08 0.0007 2.2455e-08 0 2.2569e-08 0 2.2572e-08 0.0007 2.2575e-08 0 2.2689e-08 0 2.2692e-08 0.0007 2.2695e-08 0 2.2809e-08 0 2.2812e-08 0.0007 2.2815e-08 0 2.2929e-08 0 2.2932e-08 0.0007 2.2935e-08 0 2.3049e-08 0 2.3052e-08 0.0007 2.3055e-08 0 2.3169e-08 0 2.3172e-08 0.0007 2.3175e-08 0 2.3289e-08 0 2.3292e-08 0.0007 2.3295e-08 0 2.3409e-08 0 2.3412e-08 0.0007 2.3415e-08 0 2.3529e-08 0 2.3532e-08 0.0007 2.3535e-08 0 2.3649e-08 0 2.3652e-08 0.0007 2.3655e-08 0 2.3769e-08 0 2.3772e-08 0.0007 2.3775e-08 0 2.3889e-08 0 2.3892e-08 0.0007 2.3895e-08 0 2.4009e-08 0 2.4012e-08 0.0007 2.4015e-08 0 2.4129e-08 0 2.4132e-08 0.0007 2.4135e-08 0 2.4249e-08 0 2.4252e-08 0.0007 2.4255e-08 0 2.4369e-08 0 2.4372e-08 0.0007 2.4375e-08 0 2.4489e-08 0 2.4492e-08 0.0007 2.4495e-08 0 2.4609e-08 0 2.4612e-08 0.0007 2.4615e-08 0 2.4729e-08 0 2.4732e-08 0.0007 2.4735e-08 0 2.4849e-08 0 2.4852e-08 0.0007 2.4855e-08 0 2.4969e-08 0 2.4972e-08 0.0007 2.4975e-08 0 2.5089e-08 0 2.5092e-08 0.0007 2.5095e-08 0 2.5209e-08 0 2.5212e-08 0.0007 2.5215e-08 0 2.5329e-08 0 2.5332e-08 0.0007 2.5335e-08 0 2.5449e-08 0 2.5452e-08 0.0007 2.5455e-08 0 2.5569e-08 0 2.5572e-08 0.0007 2.5575e-08 0 2.5689e-08 0 2.5692e-08 0.0007 2.5695e-08 0 2.5809e-08 0 2.5812e-08 0.0007 2.5815e-08 0 2.5929e-08 0 2.5932e-08 0.0007 2.5935e-08 0 2.6049e-08 0 2.6052e-08 0.0007 2.6055e-08 0 2.6169e-08 0 2.6172e-08 0.0007 2.6175e-08 0 2.6289e-08 0 2.6292e-08 0.0007 2.6295e-08 0 2.6409e-08 0 2.6412e-08 0.0007 2.6415e-08 0 2.6529e-08 0 2.6532e-08 0.0007 2.6535e-08 0 2.6649e-08 0 2.6652e-08 0.0007 2.6655e-08 0 2.6769e-08 0 2.6772e-08 0.0007 2.6775e-08 0 2.6889e-08 0 2.6892e-08 0.0007 2.6895e-08 0 2.7009e-08 0 2.7012e-08 0.0007 2.7015e-08 0 2.7129e-08 0 2.7132e-08 0.0007 2.7135e-08 0 2.7249e-08 0 2.7252e-08 0.0007 2.7255e-08 0 2.7369e-08 0 2.7372e-08 0.0007 2.7375e-08 0 2.7489e-08 0 2.7492e-08 0.0007 2.7495e-08 0 2.7609e-08 0 2.7612e-08 0.0007 2.7615e-08 0 2.7729e-08 0 2.7732e-08 0.0007 2.7735e-08 0 2.7849e-08 0 2.7852e-08 0.0007 2.7855e-08 0 2.7969e-08 0 2.7972e-08 0.0007 2.7975e-08 0 2.8089e-08 0 2.8092e-08 0.0007 2.8095e-08 0 2.8209e-08 0 2.8212e-08 0.0007 2.8215e-08 0 2.8329e-08 0 2.8332e-08 0.0007 2.8335e-08 0 2.8449e-08 0 2.8452e-08 0.0007 2.8455e-08 0 2.8569e-08 0 2.8572e-08 0.0007 2.8575e-08 0 2.8689e-08 0 2.8692e-08 0.0007 2.8695e-08 0 2.8809e-08 0 2.8812e-08 0.0007 2.8815e-08 0 2.8929e-08 0 2.8932e-08 0.0007 2.8935e-08 0 2.9049e-08 0 2.9052e-08 0.0007 2.9055e-08 0 2.9169e-08 0 2.9172e-08 0.0007 2.9175e-08 0 2.9289e-08 0 2.9292e-08 0.0007 2.9295e-08 0 2.9409e-08 0 2.9412e-08 0.0007 2.9415e-08 0 2.9529e-08 0 2.9532e-08 0.0007 2.9535e-08 0 2.9649e-08 0 2.9652e-08 0.0007 2.9655e-08 0 2.9769e-08 0 2.9772e-08 0.0007 2.9775e-08 0 2.9889e-08 0 2.9892e-08 0.0007 2.9895e-08 0 3.0009e-08 0 3.0012e-08 0.0007 3.0015e-08 0 3.0129e-08 0 3.0132e-08 0.0007 3.0135e-08 0 3.0249e-08 0 3.0252e-08 0.0007 3.0255e-08 0 3.0369e-08 0 3.0372e-08 0.0007 3.0375e-08 0 3.0489e-08 0 3.0492e-08 0.0007 3.0495e-08 0 3.0609e-08 0 3.0612e-08 0.0007 3.0615e-08 0 3.0729e-08 0 3.0732e-08 0.0007 3.0735e-08 0 3.0849e-08 0 3.0852e-08 0.0007 3.0855e-08 0 3.0969e-08 0 3.0972e-08 0.0007 3.0975e-08 0 3.1089e-08 0 3.1092e-08 0.0007 3.1095e-08 0 3.1209e-08 0 3.1212e-08 0.0007 3.1215e-08 0 3.1329e-08 0 3.1332e-08 0.0007 3.1335e-08 0 3.1449e-08 0 3.1452e-08 0.0007 3.1455e-08 0 3.1569e-08 0 3.1572e-08 0.0007 3.1575e-08 0 3.1689e-08 0 3.1692e-08 0.0007 3.1695e-08 0 3.1809e-08 0 3.1812e-08 0.0007 3.1815e-08 0 3.1929e-08 0 3.1932e-08 0.0007 3.1935e-08 0 3.2049e-08 0 3.2052e-08 0.0007 3.2055e-08 0 3.2169e-08 0 3.2172e-08 0.0007 3.2175e-08 0 3.2289e-08 0 3.2292e-08 0.0007 3.2295e-08 0 3.2409e-08 0 3.2412e-08 0.0007 3.2415e-08 0 3.2529e-08 0 3.2532e-08 0.0007 3.2535e-08 0 3.2649e-08 0 3.2652e-08 0.0007 3.2655e-08 0 3.2769e-08 0 3.2772e-08 0.0007 3.2775e-08 0 3.2889e-08 0 3.2892e-08 0.0007 3.2895e-08 0 3.3009e-08 0 3.3012e-08 0.0007 3.3015e-08 0 3.3129e-08 0 3.3132e-08 0.0007 3.3135e-08 0 3.3249e-08 0 3.3252e-08 0.0007 3.3255e-08 0 3.3369e-08 0 3.3372e-08 0.0007 3.3375e-08 0 3.3489e-08 0 3.3492e-08 0.0007 3.3495e-08 0 3.3609e-08 0 3.3612e-08 0.0007 3.3615e-08 0 3.3729e-08 0 3.3732e-08 0.0007 3.3735e-08 0 3.3849e-08 0 3.3852e-08 0.0007 3.3855e-08 0 3.3969e-08 0 3.3972e-08 0.0007 3.3975e-08 0 3.4089e-08 0 3.4092e-08 0.0007 3.4095e-08 0 3.4209e-08 0 3.4212e-08 0.0007 3.4215e-08 0 3.4329e-08 0 3.4332e-08 0.0007 3.4335e-08 0 3.4449e-08 0 3.4452e-08 0.0007 3.4455e-08 0 3.4569e-08 0 3.4572e-08 0.0007 3.4575e-08 0 3.4689e-08 0 3.4692e-08 0.0007 3.4695e-08 0 3.4809e-08 0 3.4812e-08 0.0007 3.4815e-08 0 3.4929e-08 0 3.4932e-08 0.0007 3.4935e-08 0 3.5049e-08 0 3.5052e-08 0.0007 3.5055e-08 0 3.5169e-08 0 3.5172e-08 0.0007 3.5175e-08 0 3.5289e-08 0 3.5292e-08 0.0007 3.5295e-08 0 3.5409e-08 0 3.5412e-08 0.0007 3.5415e-08 0 3.5529e-08 0 3.5532e-08 0.0007 3.5535e-08 0 3.5649e-08 0 3.5652e-08 0.0007 3.5655e-08 0 3.5769e-08 0 3.5772e-08 0.0007 3.5775e-08 0 3.5889e-08 0 3.5892e-08 0.0007 3.5895e-08 0 3.6009e-08 0 3.6012e-08 0.0007 3.6015e-08 0 3.6129e-08 0 3.6132e-08 0.0007 3.6135e-08 0 3.6249e-08 0 3.6252e-08 0.0007 3.6255e-08 0 3.6369e-08 0 3.6372e-08 0.0007 3.6375e-08 0 3.6489e-08 0 3.6492e-08 0.0007 3.6495e-08 0 3.6609e-08 0 3.6612e-08 0.0007 3.6615e-08 0 3.6729e-08 0 3.6732e-08 0.0007 3.6735e-08 0 3.6849e-08 0 3.6852e-08 0.0007 3.6855e-08 0 3.6969e-08 0 3.6972e-08 0.0007 3.6975e-08 0 3.7089e-08 0 3.7092e-08 0.0007 3.7095e-08 0 3.7209e-08 0 3.7212e-08 0.0007 3.7215e-08 0 3.7329e-08 0 3.7332e-08 0.0007 3.7335e-08 0 3.7449e-08 0 3.7452e-08 0.0007 3.7455e-08 0 3.7569e-08 0 3.7572e-08 0.0007 3.7575e-08 0 3.7689e-08 0 3.7692e-08 0.0007 3.7695e-08 0 3.7809e-08 0 3.7812e-08 0.0007 3.7815e-08 0 3.7929e-08 0 3.7932e-08 0.0007 3.7935e-08 0 3.8049e-08 0 3.8052e-08 0.0007 3.8055e-08 0 3.8169e-08 0 3.8172e-08 0.0007 3.8175e-08 0 3.8289e-08 0 3.8292e-08 0.0007 3.8295e-08 0 3.8409e-08 0 3.8412e-08 0.0007 3.8415e-08 0 3.8529e-08 0 3.8532e-08 0.0007 3.8535e-08 0 3.8649e-08 0 3.8652e-08 0.0007 3.8655e-08 0 3.8769e-08 0 3.8772e-08 0.0007 3.8775e-08 0 3.8889e-08 0 3.8892e-08 0.0007 3.8895e-08 0 3.9009e-08 0 3.9012e-08 0.0007 3.9015e-08 0 3.9129e-08 0 3.9132e-08 0.0007 3.9135e-08 0 3.9249e-08 0 3.9252e-08 0.0007 3.9255e-08 0 3.9369e-08 0 3.9372e-08 0.0007 3.9375e-08 0 3.9489e-08 0 3.9492e-08 0.0007 3.9495e-08 0 3.9609e-08 0 3.9612e-08 0.0007 3.9615e-08 0 3.9729e-08 0 3.9732e-08 0.0007 3.9735e-08 0 3.9849e-08 0 3.9852e-08 0.0007 3.9855e-08 0 3.9969e-08 0 3.9972e-08 0.0007 3.9975e-08 0 4.0089e-08 0 4.0092e-08 0.0007 4.0095e-08 0 4.0209e-08 0 4.0212e-08 0.0007 4.0215e-08 0 4.0329e-08 0 4.0332e-08 0.0007 4.0335e-08 0 4.0449e-08 0 4.0452e-08 0.0007 4.0455e-08 0 4.0569e-08 0 4.0572e-08 0.0007 4.0575e-08 0 4.0689e-08 0 4.0692e-08 0.0007 4.0695e-08 0 4.0809e-08 0 4.0812e-08 0.0007 4.0815e-08 0 4.0929e-08 0 4.0932e-08 0.0007 4.0935e-08 0 4.1049e-08 0 4.1052e-08 0.0007 4.1055e-08 0 4.1169e-08 0 4.1172e-08 0.0007 4.1175e-08 0 4.1289e-08 0 4.1292e-08 0.0007 4.1295e-08 0 4.1409e-08 0 4.1412e-08 0.0007 4.1415e-08 0 4.1529e-08 0 4.1532e-08 0.0007 4.1535e-08 0 4.1649e-08 0 4.1652e-08 0.0007 4.1655e-08 0 4.1769e-08 0 4.1772e-08 0.0007 4.1775e-08 0 4.1889e-08 0 4.1892e-08 0.0007 4.1895e-08 0 4.2009e-08 0 4.2012e-08 0.0007 4.2015e-08 0 4.2129e-08 0 4.2132e-08 0.0007 4.2135e-08 0 4.2249e-08 0 4.2252e-08 0.0007 4.2255e-08 0 4.2369e-08 0 4.2372e-08 0.0007 4.2375e-08 0 4.2489e-08 0 4.2492e-08 0.0007 4.2495e-08 0 4.2609e-08 0 4.2612e-08 0.0007 4.2615e-08 0 4.2729e-08 0 4.2732e-08 0.0007 4.2735e-08 0 4.2849e-08 0 4.2852e-08 0.0007 4.2855e-08 0 4.2969e-08 0 4.2972e-08 0.0007 4.2975e-08 0 4.3089e-08 0 4.3092e-08 0.0007 4.3095e-08 0 4.3209e-08 0 4.3212e-08 0.0007 4.3215e-08 0 4.3329e-08 0 4.3332e-08 0.0007 4.3335e-08 0 4.3449e-08 0 4.3452e-08 0.0007 4.3455e-08 0 4.3569e-08 0 4.3572e-08 0.0007 4.3575e-08 0 4.3689e-08 0 4.3692e-08 0.0007 4.3695e-08 0 4.3809e-08 0 4.3812e-08 0.0007 4.3815e-08 0 4.3929e-08 0 4.3932e-08 0.0007 4.3935e-08 0 4.4049e-08 0 4.4052e-08 0.0007 4.4055e-08 0 4.4169e-08 0 4.4172e-08 0.0007 4.4175e-08 0 4.4289e-08 0 4.4292e-08 0.0007 4.4295e-08 0 4.4409e-08 0 4.4412e-08 0.0007 4.4415e-08 0 4.4529e-08 0 4.4532e-08 0.0007 4.4535e-08 0 4.4649e-08 0 4.4652e-08 0.0007 4.4655e-08 0 4.4769e-08 0 4.4772e-08 0.0007 4.4775e-08 0 4.4889e-08 0 4.4892e-08 0.0007 4.4895e-08 0 4.5009e-08 0 4.5012e-08 0.0007 4.5015e-08 0 4.5129e-08 0 4.5132e-08 0.0007 4.5135e-08 0 4.5249e-08 0 4.5252e-08 0.0007 4.5255e-08 0 4.5369e-08 0 4.5372e-08 0.0007 4.5375e-08 0 4.5489e-08 0 4.5492e-08 0.0007 4.5495e-08 0 4.5609e-08 0 4.5612e-08 0.0007 4.5615e-08 0 4.5729e-08 0 4.5732e-08 0.0007 4.5735e-08 0 4.5849e-08 0 4.5852e-08 0.0007 4.5855e-08 0 4.5969e-08 0 4.5972e-08 0.0007 4.5975e-08 0 4.6089e-08 0 4.6092e-08 0.0007 4.6095e-08 0 4.6209e-08 0 4.6212e-08 0.0007 4.6215e-08 0 4.6329e-08 0 4.6332e-08 0.0007 4.6335e-08 0 4.6449e-08 0 4.6452e-08 0.0007 4.6455e-08 0 4.6569e-08 0 4.6572e-08 0.0007 4.6575e-08 0 4.6689e-08 0 4.6692e-08 0.0007 4.6695e-08 0 4.6809e-08 0 4.6812e-08 0.0007 4.6815e-08 0 4.6929e-08 0 4.6932e-08 0.0007 4.6935e-08 0 4.7049e-08 0 4.7052e-08 0.0007 4.7055e-08 0 4.7169e-08 0 4.7172e-08 0.0007 4.7175e-08 0 4.7289e-08 0 4.7292e-08 0.0007 4.7295e-08 0 4.7409e-08 0 4.7412e-08 0.0007 4.7415e-08 0 4.7529e-08 0 4.7532e-08 0.0007 4.7535e-08 0 4.7649e-08 0 4.7652e-08 0.0007 4.7655e-08 0 4.7769e-08 0 4.7772e-08 0.0007 4.7775e-08 0)
L_DFF_IP3_12|1 IP3_1_OUT_RX _DFF_IP3_12|A1  2.067833848e-12
L_DFF_IP3_12|2 _DFF_IP3_12|A1 _DFF_IP3_12|A2  4.135667696e-12
L_DFF_IP3_12|3 _DFF_IP3_12|A3 _DFF_IP3_12|A4  8.271335392e-12
L_DFF_IP3_12|T D13 _DFF_IP3_12|T1  2.067833848e-12
L_DFF_IP3_12|4 _DFF_IP3_12|T1 _DFF_IP3_12|T2  4.135667696e-12
L_DFF_IP3_12|5 _DFF_IP3_12|A4 _DFF_IP3_12|Q1  4.135667696e-12
L_DFF_IP3_12|6 _DFF_IP3_12|Q1 IP3_2_OUT  2.067833848e-12
IT12|T 0 T12  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0 2.4003e-08 0 2.4006e-08 0.0007 2.4009e-08 0 2.4123e-08 0 2.4126e-08 0.0007 2.4129e-08 0 2.4243e-08 0 2.4246e-08 0.0007 2.4249e-08 0 2.4363e-08 0 2.4366e-08 0.0007 2.4369e-08 0 2.4483e-08 0 2.4486e-08 0.0007 2.4489e-08 0 2.4603e-08 0 2.4606e-08 0.0007 2.4609e-08 0 2.4723e-08 0 2.4726e-08 0.0007 2.4729e-08 0 2.4843e-08 0 2.4846e-08 0.0007 2.4849e-08 0 2.4963e-08 0 2.4966e-08 0.0007 2.4969e-08 0 2.5083e-08 0 2.5086e-08 0.0007 2.5089e-08 0 2.5203e-08 0 2.5206e-08 0.0007 2.5209e-08 0 2.5323e-08 0 2.5326e-08 0.0007 2.5329e-08 0 2.5443e-08 0 2.5446e-08 0.0007 2.5449e-08 0 2.5563e-08 0 2.5566e-08 0.0007 2.5569e-08 0 2.5683e-08 0 2.5686e-08 0.0007 2.5689e-08 0 2.5803e-08 0 2.5806e-08 0.0007 2.5809e-08 0 2.5923e-08 0 2.5926e-08 0.0007 2.5929e-08 0 2.6043e-08 0 2.6046e-08 0.0007 2.6049e-08 0 2.6163e-08 0 2.6166e-08 0.0007 2.6169e-08 0 2.6283e-08 0 2.6286e-08 0.0007 2.6289e-08 0 2.6403e-08 0 2.6406e-08 0.0007 2.6409e-08 0 2.6523e-08 0 2.6526e-08 0.0007 2.6529e-08 0 2.6643e-08 0 2.6646e-08 0.0007 2.6649e-08 0 2.6763e-08 0 2.6766e-08 0.0007 2.6769e-08 0 2.6883e-08 0 2.6886e-08 0.0007 2.6889e-08 0 2.7003e-08 0 2.7006e-08 0.0007 2.7009e-08 0 2.7123e-08 0 2.7126e-08 0.0007 2.7129e-08 0 2.7243e-08 0 2.7246e-08 0.0007 2.7249e-08 0 2.7363e-08 0 2.7366e-08 0.0007 2.7369e-08 0 2.7483e-08 0 2.7486e-08 0.0007 2.7489e-08 0 2.7603e-08 0 2.7606e-08 0.0007 2.7609e-08 0 2.7723e-08 0 2.7726e-08 0.0007 2.7729e-08 0 2.7843e-08 0 2.7846e-08 0.0007 2.7849e-08 0 2.7963e-08 0 2.7966e-08 0.0007 2.7969e-08 0 2.8083e-08 0 2.8086e-08 0.0007 2.8089e-08 0 2.8203e-08 0 2.8206e-08 0.0007 2.8209e-08 0 2.8323e-08 0 2.8326e-08 0.0007 2.8329e-08 0 2.8443e-08 0 2.8446e-08 0.0007 2.8449e-08 0 2.8563e-08 0 2.8566e-08 0.0007 2.8569e-08 0 2.8683e-08 0 2.8686e-08 0.0007 2.8689e-08 0 2.8803e-08 0 2.8806e-08 0.0007 2.8809e-08 0 2.8923e-08 0 2.8926e-08 0.0007 2.8929e-08 0 2.9043e-08 0 2.9046e-08 0.0007 2.9049e-08 0 2.9163e-08 0 2.9166e-08 0.0007 2.9169e-08 0 2.9283e-08 0 2.9286e-08 0.0007 2.9289e-08 0 2.9403e-08 0 2.9406e-08 0.0007 2.9409e-08 0 2.9523e-08 0 2.9526e-08 0.0007 2.9529e-08 0 2.9643e-08 0 2.9646e-08 0.0007 2.9649e-08 0 2.9763e-08 0 2.9766e-08 0.0007 2.9769e-08 0 2.9883e-08 0 2.9886e-08 0.0007 2.9889e-08 0 3.0003e-08 0 3.0006e-08 0.0007 3.0009e-08 0 3.0123e-08 0 3.0126e-08 0.0007 3.0129e-08 0 3.0243e-08 0 3.0246e-08 0.0007 3.0249e-08 0 3.0363e-08 0 3.0366e-08 0.0007 3.0369e-08 0 3.0483e-08 0 3.0486e-08 0.0007 3.0489e-08 0 3.0603e-08 0 3.0606e-08 0.0007 3.0609e-08 0 3.0723e-08 0 3.0726e-08 0.0007 3.0729e-08 0 3.0843e-08 0 3.0846e-08 0.0007 3.0849e-08 0 3.0963e-08 0 3.0966e-08 0.0007 3.0969e-08 0 3.1083e-08 0 3.1086e-08 0.0007 3.1089e-08 0 3.1203e-08 0 3.1206e-08 0.0007 3.1209e-08 0 3.1323e-08 0 3.1326e-08 0.0007 3.1329e-08 0 3.1443e-08 0 3.1446e-08 0.0007 3.1449e-08 0 3.1563e-08 0 3.1566e-08 0.0007 3.1569e-08 0 3.1683e-08 0 3.1686e-08 0.0007 3.1689e-08 0 3.1803e-08 0 3.1806e-08 0.0007 3.1809e-08 0 3.1923e-08 0 3.1926e-08 0.0007 3.1929e-08 0 3.2043e-08 0 3.2046e-08 0.0007 3.2049e-08 0 3.2163e-08 0 3.2166e-08 0.0007 3.2169e-08 0 3.2283e-08 0 3.2286e-08 0.0007 3.2289e-08 0 3.2403e-08 0 3.2406e-08 0.0007 3.2409e-08 0 3.2523e-08 0 3.2526e-08 0.0007 3.2529e-08 0 3.2643e-08 0 3.2646e-08 0.0007 3.2649e-08 0 3.2763e-08 0 3.2766e-08 0.0007 3.2769e-08 0 3.2883e-08 0 3.2886e-08 0.0007 3.2889e-08 0 3.3003e-08 0 3.3006e-08 0.0007 3.3009e-08 0 3.3123e-08 0 3.3126e-08 0.0007 3.3129e-08 0 3.3243e-08 0 3.3246e-08 0.0007 3.3249e-08 0 3.3363e-08 0 3.3366e-08 0.0007 3.3369e-08 0 3.3483e-08 0 3.3486e-08 0.0007 3.3489e-08 0 3.3603e-08 0 3.3606e-08 0.0007 3.3609e-08 0 3.3723e-08 0 3.3726e-08 0.0007 3.3729e-08 0 3.3843e-08 0 3.3846e-08 0.0007 3.3849e-08 0 3.3963e-08 0 3.3966e-08 0.0007 3.3969e-08 0 3.4083e-08 0 3.4086e-08 0.0007 3.4089e-08 0 3.4203e-08 0 3.4206e-08 0.0007 3.4209e-08 0 3.4323e-08 0 3.4326e-08 0.0007 3.4329e-08 0 3.4443e-08 0 3.4446e-08 0.0007 3.4449e-08 0 3.4563e-08 0 3.4566e-08 0.0007 3.4569e-08 0 3.4683e-08 0 3.4686e-08 0.0007 3.4689e-08 0 3.4803e-08 0 3.4806e-08 0.0007 3.4809e-08 0 3.4923e-08 0 3.4926e-08 0.0007 3.4929e-08 0 3.5043e-08 0 3.5046e-08 0.0007 3.5049e-08 0 3.5163e-08 0 3.5166e-08 0.0007 3.5169e-08 0 3.5283e-08 0 3.5286e-08 0.0007 3.5289e-08 0 3.5403e-08 0 3.5406e-08 0.0007 3.5409e-08 0 3.5523e-08 0 3.5526e-08 0.0007 3.5529e-08 0 3.5643e-08 0 3.5646e-08 0.0007 3.5649e-08 0 3.5763e-08 0 3.5766e-08 0.0007 3.5769e-08 0 3.5883e-08 0 3.5886e-08 0.0007 3.5889e-08 0 3.6003e-08 0 3.6006e-08 0.0007 3.6009e-08 0 3.6123e-08 0 3.6126e-08 0.0007 3.6129e-08 0 3.6243e-08 0 3.6246e-08 0.0007 3.6249e-08 0 3.6363e-08 0 3.6366e-08 0.0007 3.6369e-08 0 3.6483e-08 0 3.6486e-08 0.0007 3.6489e-08 0 3.6603e-08 0 3.6606e-08 0.0007 3.6609e-08 0 3.6723e-08 0 3.6726e-08 0.0007 3.6729e-08 0 3.6843e-08 0 3.6846e-08 0.0007 3.6849e-08 0 3.6963e-08 0 3.6966e-08 0.0007 3.6969e-08 0 3.7083e-08 0 3.7086e-08 0.0007 3.7089e-08 0 3.7203e-08 0 3.7206e-08 0.0007 3.7209e-08 0 3.7323e-08 0 3.7326e-08 0.0007 3.7329e-08 0 3.7443e-08 0 3.7446e-08 0.0007 3.7449e-08 0 3.7563e-08 0 3.7566e-08 0.0007 3.7569e-08 0 3.7683e-08 0 3.7686e-08 0.0007 3.7689e-08 0 3.7803e-08 0 3.7806e-08 0.0007 3.7809e-08 0 3.7923e-08 0 3.7926e-08 0.0007 3.7929e-08 0 3.8043e-08 0 3.8046e-08 0.0007 3.8049e-08 0 3.8163e-08 0 3.8166e-08 0.0007 3.8169e-08 0 3.8283e-08 0 3.8286e-08 0.0007 3.8289e-08 0 3.8403e-08 0 3.8406e-08 0.0007 3.8409e-08 0 3.8523e-08 0 3.8526e-08 0.0007 3.8529e-08 0 3.8643e-08 0 3.8646e-08 0.0007 3.8649e-08 0 3.8763e-08 0 3.8766e-08 0.0007 3.8769e-08 0 3.8883e-08 0 3.8886e-08 0.0007 3.8889e-08 0 3.9003e-08 0 3.9006e-08 0.0007 3.9009e-08 0 3.9123e-08 0 3.9126e-08 0.0007 3.9129e-08 0 3.9243e-08 0 3.9246e-08 0.0007 3.9249e-08 0 3.9363e-08 0 3.9366e-08 0.0007 3.9369e-08 0 3.9483e-08 0 3.9486e-08 0.0007 3.9489e-08 0 3.9603e-08 0 3.9606e-08 0.0007 3.9609e-08 0 3.9723e-08 0 3.9726e-08 0.0007 3.9729e-08 0 3.9843e-08 0 3.9846e-08 0.0007 3.9849e-08 0 3.9963e-08 0 3.9966e-08 0.0007 3.9969e-08 0 4.0083e-08 0 4.0086e-08 0.0007 4.0089e-08 0 4.0203e-08 0 4.0206e-08 0.0007 4.0209e-08 0 4.0323e-08 0 4.0326e-08 0.0007 4.0329e-08 0 4.0443e-08 0 4.0446e-08 0.0007 4.0449e-08 0 4.0563e-08 0 4.0566e-08 0.0007 4.0569e-08 0 4.0683e-08 0 4.0686e-08 0.0007 4.0689e-08 0 4.0803e-08 0 4.0806e-08 0.0007 4.0809e-08 0 4.0923e-08 0 4.0926e-08 0.0007 4.0929e-08 0 4.1043e-08 0 4.1046e-08 0.0007 4.1049e-08 0 4.1163e-08 0 4.1166e-08 0.0007 4.1169e-08 0 4.1283e-08 0 4.1286e-08 0.0007 4.1289e-08 0 4.1403e-08 0 4.1406e-08 0.0007 4.1409e-08 0 4.1523e-08 0 4.1526e-08 0.0007 4.1529e-08 0 4.1643e-08 0 4.1646e-08 0.0007 4.1649e-08 0 4.1763e-08 0 4.1766e-08 0.0007 4.1769e-08 0 4.1883e-08 0 4.1886e-08 0.0007 4.1889e-08 0 4.2003e-08 0 4.2006e-08 0.0007 4.2009e-08 0 4.2123e-08 0 4.2126e-08 0.0007 4.2129e-08 0 4.2243e-08 0 4.2246e-08 0.0007 4.2249e-08 0 4.2363e-08 0 4.2366e-08 0.0007 4.2369e-08 0 4.2483e-08 0 4.2486e-08 0.0007 4.2489e-08 0 4.2603e-08 0 4.2606e-08 0.0007 4.2609e-08 0 4.2723e-08 0 4.2726e-08 0.0007 4.2729e-08 0 4.2843e-08 0 4.2846e-08 0.0007 4.2849e-08 0 4.2963e-08 0 4.2966e-08 0.0007 4.2969e-08 0 4.3083e-08 0 4.3086e-08 0.0007 4.3089e-08 0 4.3203e-08 0 4.3206e-08 0.0007 4.3209e-08 0 4.3323e-08 0 4.3326e-08 0.0007 4.3329e-08 0 4.3443e-08 0 4.3446e-08 0.0007 4.3449e-08 0 4.3563e-08 0 4.3566e-08 0.0007 4.3569e-08 0 4.3683e-08 0 4.3686e-08 0.0007 4.3689e-08 0 4.3803e-08 0 4.3806e-08 0.0007 4.3809e-08 0 4.3923e-08 0 4.3926e-08 0.0007 4.3929e-08 0 4.4043e-08 0 4.4046e-08 0.0007 4.4049e-08 0 4.4163e-08 0 4.4166e-08 0.0007 4.4169e-08 0 4.4283e-08 0 4.4286e-08 0.0007 4.4289e-08 0 4.4403e-08 0 4.4406e-08 0.0007 4.4409e-08 0 4.4523e-08 0 4.4526e-08 0.0007 4.4529e-08 0 4.4643e-08 0 4.4646e-08 0.0007 4.4649e-08 0 4.4763e-08 0 4.4766e-08 0.0007 4.4769e-08 0 4.4883e-08 0 4.4886e-08 0.0007 4.4889e-08 0 4.5003e-08 0 4.5006e-08 0.0007 4.5009e-08 0 4.5123e-08 0 4.5126e-08 0.0007 4.5129e-08 0 4.5243e-08 0 4.5246e-08 0.0007 4.5249e-08 0 4.5363e-08 0 4.5366e-08 0.0007 4.5369e-08 0 4.5483e-08 0 4.5486e-08 0.0007 4.5489e-08 0 4.5603e-08 0 4.5606e-08 0.0007 4.5609e-08 0 4.5723e-08 0 4.5726e-08 0.0007 4.5729e-08 0 4.5843e-08 0 4.5846e-08 0.0007 4.5849e-08 0 4.5963e-08 0 4.5966e-08 0.0007 4.5969e-08 0 4.6083e-08 0 4.6086e-08 0.0007 4.6089e-08 0 4.6203e-08 0 4.6206e-08 0.0007 4.6209e-08 0 4.6323e-08 0 4.6326e-08 0.0007 4.6329e-08 0 4.6443e-08 0 4.6446e-08 0.0007 4.6449e-08 0 4.6563e-08 0 4.6566e-08 0.0007 4.6569e-08 0 4.6683e-08 0 4.6686e-08 0.0007 4.6689e-08 0 4.6803e-08 0 4.6806e-08 0.0007 4.6809e-08 0 4.6923e-08 0 4.6926e-08 0.0007 4.6929e-08 0 4.7043e-08 0 4.7046e-08 0.0007 4.7049e-08 0 4.7163e-08 0 4.7166e-08 0.0007 4.7169e-08 0 4.7283e-08 0 4.7286e-08 0.0007 4.7289e-08 0 4.7403e-08 0 4.7406e-08 0.0007 4.7409e-08 0 4.7523e-08 0 4.7526e-08 0.0007 4.7529e-08 0 4.7643e-08 0 4.7646e-08 0.0007 4.7649e-08 0 4.7763e-08 0 4.7766e-08 0.0007 4.7769e-08 0)
L_S0|1 P0_2_RX _S0|A1  2.067833848e-12
L_S0|2 _S0|A1 _S0|A2  4.135667696e-12
L_S0|3 _S0|A3 _S0|A4  8.271335392e-12
L_S0|T T12 _S0|T1  2.067833848e-12
L_S0|4 _S0|T1 _S0|T2  4.135667696e-12
L_S0|5 _S0|A4 _S0|Q1  4.135667696e-12
L_S0|6 _S0|Q1 S0  2.067833848e-12
IT13|T 0 T13  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0 2.4003e-08 0 2.4006e-08 0.0007 2.4009e-08 0 2.4123e-08 0 2.4126e-08 0.0007 2.4129e-08 0 2.4243e-08 0 2.4246e-08 0.0007 2.4249e-08 0 2.4363e-08 0 2.4366e-08 0.0007 2.4369e-08 0 2.4483e-08 0 2.4486e-08 0.0007 2.4489e-08 0 2.4603e-08 0 2.4606e-08 0.0007 2.4609e-08 0 2.4723e-08 0 2.4726e-08 0.0007 2.4729e-08 0 2.4843e-08 0 2.4846e-08 0.0007 2.4849e-08 0 2.4963e-08 0 2.4966e-08 0.0007 2.4969e-08 0 2.5083e-08 0 2.5086e-08 0.0007 2.5089e-08 0 2.5203e-08 0 2.5206e-08 0.0007 2.5209e-08 0 2.5323e-08 0 2.5326e-08 0.0007 2.5329e-08 0 2.5443e-08 0 2.5446e-08 0.0007 2.5449e-08 0 2.5563e-08 0 2.5566e-08 0.0007 2.5569e-08 0 2.5683e-08 0 2.5686e-08 0.0007 2.5689e-08 0 2.5803e-08 0 2.5806e-08 0.0007 2.5809e-08 0 2.5923e-08 0 2.5926e-08 0.0007 2.5929e-08 0 2.6043e-08 0 2.6046e-08 0.0007 2.6049e-08 0 2.6163e-08 0 2.6166e-08 0.0007 2.6169e-08 0 2.6283e-08 0 2.6286e-08 0.0007 2.6289e-08 0 2.6403e-08 0 2.6406e-08 0.0007 2.6409e-08 0 2.6523e-08 0 2.6526e-08 0.0007 2.6529e-08 0 2.6643e-08 0 2.6646e-08 0.0007 2.6649e-08 0 2.6763e-08 0 2.6766e-08 0.0007 2.6769e-08 0 2.6883e-08 0 2.6886e-08 0.0007 2.6889e-08 0 2.7003e-08 0 2.7006e-08 0.0007 2.7009e-08 0 2.7123e-08 0 2.7126e-08 0.0007 2.7129e-08 0 2.7243e-08 0 2.7246e-08 0.0007 2.7249e-08 0 2.7363e-08 0 2.7366e-08 0.0007 2.7369e-08 0 2.7483e-08 0 2.7486e-08 0.0007 2.7489e-08 0 2.7603e-08 0 2.7606e-08 0.0007 2.7609e-08 0 2.7723e-08 0 2.7726e-08 0.0007 2.7729e-08 0 2.7843e-08 0 2.7846e-08 0.0007 2.7849e-08 0 2.7963e-08 0 2.7966e-08 0.0007 2.7969e-08 0 2.8083e-08 0 2.8086e-08 0.0007 2.8089e-08 0 2.8203e-08 0 2.8206e-08 0.0007 2.8209e-08 0 2.8323e-08 0 2.8326e-08 0.0007 2.8329e-08 0 2.8443e-08 0 2.8446e-08 0.0007 2.8449e-08 0 2.8563e-08 0 2.8566e-08 0.0007 2.8569e-08 0 2.8683e-08 0 2.8686e-08 0.0007 2.8689e-08 0 2.8803e-08 0 2.8806e-08 0.0007 2.8809e-08 0 2.8923e-08 0 2.8926e-08 0.0007 2.8929e-08 0 2.9043e-08 0 2.9046e-08 0.0007 2.9049e-08 0 2.9163e-08 0 2.9166e-08 0.0007 2.9169e-08 0 2.9283e-08 0 2.9286e-08 0.0007 2.9289e-08 0 2.9403e-08 0 2.9406e-08 0.0007 2.9409e-08 0 2.9523e-08 0 2.9526e-08 0.0007 2.9529e-08 0 2.9643e-08 0 2.9646e-08 0.0007 2.9649e-08 0 2.9763e-08 0 2.9766e-08 0.0007 2.9769e-08 0 2.9883e-08 0 2.9886e-08 0.0007 2.9889e-08 0 3.0003e-08 0 3.0006e-08 0.0007 3.0009e-08 0 3.0123e-08 0 3.0126e-08 0.0007 3.0129e-08 0 3.0243e-08 0 3.0246e-08 0.0007 3.0249e-08 0 3.0363e-08 0 3.0366e-08 0.0007 3.0369e-08 0 3.0483e-08 0 3.0486e-08 0.0007 3.0489e-08 0 3.0603e-08 0 3.0606e-08 0.0007 3.0609e-08 0 3.0723e-08 0 3.0726e-08 0.0007 3.0729e-08 0 3.0843e-08 0 3.0846e-08 0.0007 3.0849e-08 0 3.0963e-08 0 3.0966e-08 0.0007 3.0969e-08 0 3.1083e-08 0 3.1086e-08 0.0007 3.1089e-08 0 3.1203e-08 0 3.1206e-08 0.0007 3.1209e-08 0 3.1323e-08 0 3.1326e-08 0.0007 3.1329e-08 0 3.1443e-08 0 3.1446e-08 0.0007 3.1449e-08 0 3.1563e-08 0 3.1566e-08 0.0007 3.1569e-08 0 3.1683e-08 0 3.1686e-08 0.0007 3.1689e-08 0 3.1803e-08 0 3.1806e-08 0.0007 3.1809e-08 0 3.1923e-08 0 3.1926e-08 0.0007 3.1929e-08 0 3.2043e-08 0 3.2046e-08 0.0007 3.2049e-08 0 3.2163e-08 0 3.2166e-08 0.0007 3.2169e-08 0 3.2283e-08 0 3.2286e-08 0.0007 3.2289e-08 0 3.2403e-08 0 3.2406e-08 0.0007 3.2409e-08 0 3.2523e-08 0 3.2526e-08 0.0007 3.2529e-08 0 3.2643e-08 0 3.2646e-08 0.0007 3.2649e-08 0 3.2763e-08 0 3.2766e-08 0.0007 3.2769e-08 0 3.2883e-08 0 3.2886e-08 0.0007 3.2889e-08 0 3.3003e-08 0 3.3006e-08 0.0007 3.3009e-08 0 3.3123e-08 0 3.3126e-08 0.0007 3.3129e-08 0 3.3243e-08 0 3.3246e-08 0.0007 3.3249e-08 0 3.3363e-08 0 3.3366e-08 0.0007 3.3369e-08 0 3.3483e-08 0 3.3486e-08 0.0007 3.3489e-08 0 3.3603e-08 0 3.3606e-08 0.0007 3.3609e-08 0 3.3723e-08 0 3.3726e-08 0.0007 3.3729e-08 0 3.3843e-08 0 3.3846e-08 0.0007 3.3849e-08 0 3.3963e-08 0 3.3966e-08 0.0007 3.3969e-08 0 3.4083e-08 0 3.4086e-08 0.0007 3.4089e-08 0 3.4203e-08 0 3.4206e-08 0.0007 3.4209e-08 0 3.4323e-08 0 3.4326e-08 0.0007 3.4329e-08 0 3.4443e-08 0 3.4446e-08 0.0007 3.4449e-08 0 3.4563e-08 0 3.4566e-08 0.0007 3.4569e-08 0 3.4683e-08 0 3.4686e-08 0.0007 3.4689e-08 0 3.4803e-08 0 3.4806e-08 0.0007 3.4809e-08 0 3.4923e-08 0 3.4926e-08 0.0007 3.4929e-08 0 3.5043e-08 0 3.5046e-08 0.0007 3.5049e-08 0 3.5163e-08 0 3.5166e-08 0.0007 3.5169e-08 0 3.5283e-08 0 3.5286e-08 0.0007 3.5289e-08 0 3.5403e-08 0 3.5406e-08 0.0007 3.5409e-08 0 3.5523e-08 0 3.5526e-08 0.0007 3.5529e-08 0 3.5643e-08 0 3.5646e-08 0.0007 3.5649e-08 0 3.5763e-08 0 3.5766e-08 0.0007 3.5769e-08 0 3.5883e-08 0 3.5886e-08 0.0007 3.5889e-08 0 3.6003e-08 0 3.6006e-08 0.0007 3.6009e-08 0 3.6123e-08 0 3.6126e-08 0.0007 3.6129e-08 0 3.6243e-08 0 3.6246e-08 0.0007 3.6249e-08 0 3.6363e-08 0 3.6366e-08 0.0007 3.6369e-08 0 3.6483e-08 0 3.6486e-08 0.0007 3.6489e-08 0 3.6603e-08 0 3.6606e-08 0.0007 3.6609e-08 0 3.6723e-08 0 3.6726e-08 0.0007 3.6729e-08 0 3.6843e-08 0 3.6846e-08 0.0007 3.6849e-08 0 3.6963e-08 0 3.6966e-08 0.0007 3.6969e-08 0 3.7083e-08 0 3.7086e-08 0.0007 3.7089e-08 0 3.7203e-08 0 3.7206e-08 0.0007 3.7209e-08 0 3.7323e-08 0 3.7326e-08 0.0007 3.7329e-08 0 3.7443e-08 0 3.7446e-08 0.0007 3.7449e-08 0 3.7563e-08 0 3.7566e-08 0.0007 3.7569e-08 0 3.7683e-08 0 3.7686e-08 0.0007 3.7689e-08 0 3.7803e-08 0 3.7806e-08 0.0007 3.7809e-08 0 3.7923e-08 0 3.7926e-08 0.0007 3.7929e-08 0 3.8043e-08 0 3.8046e-08 0.0007 3.8049e-08 0 3.8163e-08 0 3.8166e-08 0.0007 3.8169e-08 0 3.8283e-08 0 3.8286e-08 0.0007 3.8289e-08 0 3.8403e-08 0 3.8406e-08 0.0007 3.8409e-08 0 3.8523e-08 0 3.8526e-08 0.0007 3.8529e-08 0 3.8643e-08 0 3.8646e-08 0.0007 3.8649e-08 0 3.8763e-08 0 3.8766e-08 0.0007 3.8769e-08 0 3.8883e-08 0 3.8886e-08 0.0007 3.8889e-08 0 3.9003e-08 0 3.9006e-08 0.0007 3.9009e-08 0 3.9123e-08 0 3.9126e-08 0.0007 3.9129e-08 0 3.9243e-08 0 3.9246e-08 0.0007 3.9249e-08 0 3.9363e-08 0 3.9366e-08 0.0007 3.9369e-08 0 3.9483e-08 0 3.9486e-08 0.0007 3.9489e-08 0 3.9603e-08 0 3.9606e-08 0.0007 3.9609e-08 0 3.9723e-08 0 3.9726e-08 0.0007 3.9729e-08 0 3.9843e-08 0 3.9846e-08 0.0007 3.9849e-08 0 3.9963e-08 0 3.9966e-08 0.0007 3.9969e-08 0 4.0083e-08 0 4.0086e-08 0.0007 4.0089e-08 0 4.0203e-08 0 4.0206e-08 0.0007 4.0209e-08 0 4.0323e-08 0 4.0326e-08 0.0007 4.0329e-08 0 4.0443e-08 0 4.0446e-08 0.0007 4.0449e-08 0 4.0563e-08 0 4.0566e-08 0.0007 4.0569e-08 0 4.0683e-08 0 4.0686e-08 0.0007 4.0689e-08 0 4.0803e-08 0 4.0806e-08 0.0007 4.0809e-08 0 4.0923e-08 0 4.0926e-08 0.0007 4.0929e-08 0 4.1043e-08 0 4.1046e-08 0.0007 4.1049e-08 0 4.1163e-08 0 4.1166e-08 0.0007 4.1169e-08 0 4.1283e-08 0 4.1286e-08 0.0007 4.1289e-08 0 4.1403e-08 0 4.1406e-08 0.0007 4.1409e-08 0 4.1523e-08 0 4.1526e-08 0.0007 4.1529e-08 0 4.1643e-08 0 4.1646e-08 0.0007 4.1649e-08 0 4.1763e-08 0 4.1766e-08 0.0007 4.1769e-08 0 4.1883e-08 0 4.1886e-08 0.0007 4.1889e-08 0 4.2003e-08 0 4.2006e-08 0.0007 4.2009e-08 0 4.2123e-08 0 4.2126e-08 0.0007 4.2129e-08 0 4.2243e-08 0 4.2246e-08 0.0007 4.2249e-08 0 4.2363e-08 0 4.2366e-08 0.0007 4.2369e-08 0 4.2483e-08 0 4.2486e-08 0.0007 4.2489e-08 0 4.2603e-08 0 4.2606e-08 0.0007 4.2609e-08 0 4.2723e-08 0 4.2726e-08 0.0007 4.2729e-08 0 4.2843e-08 0 4.2846e-08 0.0007 4.2849e-08 0 4.2963e-08 0 4.2966e-08 0.0007 4.2969e-08 0 4.3083e-08 0 4.3086e-08 0.0007 4.3089e-08 0 4.3203e-08 0 4.3206e-08 0.0007 4.3209e-08 0 4.3323e-08 0 4.3326e-08 0.0007 4.3329e-08 0 4.3443e-08 0 4.3446e-08 0.0007 4.3449e-08 0 4.3563e-08 0 4.3566e-08 0.0007 4.3569e-08 0 4.3683e-08 0 4.3686e-08 0.0007 4.3689e-08 0 4.3803e-08 0 4.3806e-08 0.0007 4.3809e-08 0 4.3923e-08 0 4.3926e-08 0.0007 4.3929e-08 0 4.4043e-08 0 4.4046e-08 0.0007 4.4049e-08 0 4.4163e-08 0 4.4166e-08 0.0007 4.4169e-08 0 4.4283e-08 0 4.4286e-08 0.0007 4.4289e-08 0 4.4403e-08 0 4.4406e-08 0.0007 4.4409e-08 0 4.4523e-08 0 4.4526e-08 0.0007 4.4529e-08 0 4.4643e-08 0 4.4646e-08 0.0007 4.4649e-08 0 4.4763e-08 0 4.4766e-08 0.0007 4.4769e-08 0 4.4883e-08 0 4.4886e-08 0.0007 4.4889e-08 0 4.5003e-08 0 4.5006e-08 0.0007 4.5009e-08 0 4.5123e-08 0 4.5126e-08 0.0007 4.5129e-08 0 4.5243e-08 0 4.5246e-08 0.0007 4.5249e-08 0 4.5363e-08 0 4.5366e-08 0.0007 4.5369e-08 0 4.5483e-08 0 4.5486e-08 0.0007 4.5489e-08 0 4.5603e-08 0 4.5606e-08 0.0007 4.5609e-08 0 4.5723e-08 0 4.5726e-08 0.0007 4.5729e-08 0 4.5843e-08 0 4.5846e-08 0.0007 4.5849e-08 0 4.5963e-08 0 4.5966e-08 0.0007 4.5969e-08 0 4.6083e-08 0 4.6086e-08 0.0007 4.6089e-08 0 4.6203e-08 0 4.6206e-08 0.0007 4.6209e-08 0 4.6323e-08 0 4.6326e-08 0.0007 4.6329e-08 0 4.6443e-08 0 4.6446e-08 0.0007 4.6449e-08 0 4.6563e-08 0 4.6566e-08 0.0007 4.6569e-08 0 4.6683e-08 0 4.6686e-08 0.0007 4.6689e-08 0 4.6803e-08 0 4.6806e-08 0.0007 4.6809e-08 0 4.6923e-08 0 4.6926e-08 0.0007 4.6929e-08 0 4.7043e-08 0 4.7046e-08 0.0007 4.7049e-08 0 4.7163e-08 0 4.7166e-08 0.0007 4.7169e-08 0 4.7283e-08 0 4.7286e-08 0.0007 4.7289e-08 0 4.7403e-08 0 4.7406e-08 0.0007 4.7409e-08 0 4.7523e-08 0 4.7526e-08 0.0007 4.7529e-08 0 4.7643e-08 0 4.7646e-08 0.0007 4.7649e-08 0 4.7763e-08 0 4.7766e-08 0.0007 4.7769e-08 0)
L_S1|A1 G0_2_RX _S1|A1  2.067833848e-12
L_S1|A2 _S1|A1 _S1|A2  4.135667696e-12
L_S1|A3 _S1|A3 _S1|AB  8.271335392e-12
L_S1|B1 IP1_2_OUT_RX _S1|B1  2.067833848e-12
L_S1|B2 _S1|B1 _S1|B2  4.135667696e-12
L_S1|B3 _S1|B3 _S1|AB  8.271335392e-12
L_S1|T1 T13 _S1|T1  2.067833848e-12
L_S1|T2 _S1|T1 _S1|T2  4.135667696e-12
L_S1|Q2 _S1|ABTQ _S1|Q1  4.135667696e-12
L_S1|Q1 _S1|Q1 S1  2.067833848e-12
IT14|T 0 T14  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0 2.4003e-08 0 2.4006e-08 0.0007 2.4009e-08 0 2.4123e-08 0 2.4126e-08 0.0007 2.4129e-08 0 2.4243e-08 0 2.4246e-08 0.0007 2.4249e-08 0 2.4363e-08 0 2.4366e-08 0.0007 2.4369e-08 0 2.4483e-08 0 2.4486e-08 0.0007 2.4489e-08 0 2.4603e-08 0 2.4606e-08 0.0007 2.4609e-08 0 2.4723e-08 0 2.4726e-08 0.0007 2.4729e-08 0 2.4843e-08 0 2.4846e-08 0.0007 2.4849e-08 0 2.4963e-08 0 2.4966e-08 0.0007 2.4969e-08 0 2.5083e-08 0 2.5086e-08 0.0007 2.5089e-08 0 2.5203e-08 0 2.5206e-08 0.0007 2.5209e-08 0 2.5323e-08 0 2.5326e-08 0.0007 2.5329e-08 0 2.5443e-08 0 2.5446e-08 0.0007 2.5449e-08 0 2.5563e-08 0 2.5566e-08 0.0007 2.5569e-08 0 2.5683e-08 0 2.5686e-08 0.0007 2.5689e-08 0 2.5803e-08 0 2.5806e-08 0.0007 2.5809e-08 0 2.5923e-08 0 2.5926e-08 0.0007 2.5929e-08 0 2.6043e-08 0 2.6046e-08 0.0007 2.6049e-08 0 2.6163e-08 0 2.6166e-08 0.0007 2.6169e-08 0 2.6283e-08 0 2.6286e-08 0.0007 2.6289e-08 0 2.6403e-08 0 2.6406e-08 0.0007 2.6409e-08 0 2.6523e-08 0 2.6526e-08 0.0007 2.6529e-08 0 2.6643e-08 0 2.6646e-08 0.0007 2.6649e-08 0 2.6763e-08 0 2.6766e-08 0.0007 2.6769e-08 0 2.6883e-08 0 2.6886e-08 0.0007 2.6889e-08 0 2.7003e-08 0 2.7006e-08 0.0007 2.7009e-08 0 2.7123e-08 0 2.7126e-08 0.0007 2.7129e-08 0 2.7243e-08 0 2.7246e-08 0.0007 2.7249e-08 0 2.7363e-08 0 2.7366e-08 0.0007 2.7369e-08 0 2.7483e-08 0 2.7486e-08 0.0007 2.7489e-08 0 2.7603e-08 0 2.7606e-08 0.0007 2.7609e-08 0 2.7723e-08 0 2.7726e-08 0.0007 2.7729e-08 0 2.7843e-08 0 2.7846e-08 0.0007 2.7849e-08 0 2.7963e-08 0 2.7966e-08 0.0007 2.7969e-08 0 2.8083e-08 0 2.8086e-08 0.0007 2.8089e-08 0 2.8203e-08 0 2.8206e-08 0.0007 2.8209e-08 0 2.8323e-08 0 2.8326e-08 0.0007 2.8329e-08 0 2.8443e-08 0 2.8446e-08 0.0007 2.8449e-08 0 2.8563e-08 0 2.8566e-08 0.0007 2.8569e-08 0 2.8683e-08 0 2.8686e-08 0.0007 2.8689e-08 0 2.8803e-08 0 2.8806e-08 0.0007 2.8809e-08 0 2.8923e-08 0 2.8926e-08 0.0007 2.8929e-08 0 2.9043e-08 0 2.9046e-08 0.0007 2.9049e-08 0 2.9163e-08 0 2.9166e-08 0.0007 2.9169e-08 0 2.9283e-08 0 2.9286e-08 0.0007 2.9289e-08 0 2.9403e-08 0 2.9406e-08 0.0007 2.9409e-08 0 2.9523e-08 0 2.9526e-08 0.0007 2.9529e-08 0 2.9643e-08 0 2.9646e-08 0.0007 2.9649e-08 0 2.9763e-08 0 2.9766e-08 0.0007 2.9769e-08 0 2.9883e-08 0 2.9886e-08 0.0007 2.9889e-08 0 3.0003e-08 0 3.0006e-08 0.0007 3.0009e-08 0 3.0123e-08 0 3.0126e-08 0.0007 3.0129e-08 0 3.0243e-08 0 3.0246e-08 0.0007 3.0249e-08 0 3.0363e-08 0 3.0366e-08 0.0007 3.0369e-08 0 3.0483e-08 0 3.0486e-08 0.0007 3.0489e-08 0 3.0603e-08 0 3.0606e-08 0.0007 3.0609e-08 0 3.0723e-08 0 3.0726e-08 0.0007 3.0729e-08 0 3.0843e-08 0 3.0846e-08 0.0007 3.0849e-08 0 3.0963e-08 0 3.0966e-08 0.0007 3.0969e-08 0 3.1083e-08 0 3.1086e-08 0.0007 3.1089e-08 0 3.1203e-08 0 3.1206e-08 0.0007 3.1209e-08 0 3.1323e-08 0 3.1326e-08 0.0007 3.1329e-08 0 3.1443e-08 0 3.1446e-08 0.0007 3.1449e-08 0 3.1563e-08 0 3.1566e-08 0.0007 3.1569e-08 0 3.1683e-08 0 3.1686e-08 0.0007 3.1689e-08 0 3.1803e-08 0 3.1806e-08 0.0007 3.1809e-08 0 3.1923e-08 0 3.1926e-08 0.0007 3.1929e-08 0 3.2043e-08 0 3.2046e-08 0.0007 3.2049e-08 0 3.2163e-08 0 3.2166e-08 0.0007 3.2169e-08 0 3.2283e-08 0 3.2286e-08 0.0007 3.2289e-08 0 3.2403e-08 0 3.2406e-08 0.0007 3.2409e-08 0 3.2523e-08 0 3.2526e-08 0.0007 3.2529e-08 0 3.2643e-08 0 3.2646e-08 0.0007 3.2649e-08 0 3.2763e-08 0 3.2766e-08 0.0007 3.2769e-08 0 3.2883e-08 0 3.2886e-08 0.0007 3.2889e-08 0 3.3003e-08 0 3.3006e-08 0.0007 3.3009e-08 0 3.3123e-08 0 3.3126e-08 0.0007 3.3129e-08 0 3.3243e-08 0 3.3246e-08 0.0007 3.3249e-08 0 3.3363e-08 0 3.3366e-08 0.0007 3.3369e-08 0 3.3483e-08 0 3.3486e-08 0.0007 3.3489e-08 0 3.3603e-08 0 3.3606e-08 0.0007 3.3609e-08 0 3.3723e-08 0 3.3726e-08 0.0007 3.3729e-08 0 3.3843e-08 0 3.3846e-08 0.0007 3.3849e-08 0 3.3963e-08 0 3.3966e-08 0.0007 3.3969e-08 0 3.4083e-08 0 3.4086e-08 0.0007 3.4089e-08 0 3.4203e-08 0 3.4206e-08 0.0007 3.4209e-08 0 3.4323e-08 0 3.4326e-08 0.0007 3.4329e-08 0 3.4443e-08 0 3.4446e-08 0.0007 3.4449e-08 0 3.4563e-08 0 3.4566e-08 0.0007 3.4569e-08 0 3.4683e-08 0 3.4686e-08 0.0007 3.4689e-08 0 3.4803e-08 0 3.4806e-08 0.0007 3.4809e-08 0 3.4923e-08 0 3.4926e-08 0.0007 3.4929e-08 0 3.5043e-08 0 3.5046e-08 0.0007 3.5049e-08 0 3.5163e-08 0 3.5166e-08 0.0007 3.5169e-08 0 3.5283e-08 0 3.5286e-08 0.0007 3.5289e-08 0 3.5403e-08 0 3.5406e-08 0.0007 3.5409e-08 0 3.5523e-08 0 3.5526e-08 0.0007 3.5529e-08 0 3.5643e-08 0 3.5646e-08 0.0007 3.5649e-08 0 3.5763e-08 0 3.5766e-08 0.0007 3.5769e-08 0 3.5883e-08 0 3.5886e-08 0.0007 3.5889e-08 0 3.6003e-08 0 3.6006e-08 0.0007 3.6009e-08 0 3.6123e-08 0 3.6126e-08 0.0007 3.6129e-08 0 3.6243e-08 0 3.6246e-08 0.0007 3.6249e-08 0 3.6363e-08 0 3.6366e-08 0.0007 3.6369e-08 0 3.6483e-08 0 3.6486e-08 0.0007 3.6489e-08 0 3.6603e-08 0 3.6606e-08 0.0007 3.6609e-08 0 3.6723e-08 0 3.6726e-08 0.0007 3.6729e-08 0 3.6843e-08 0 3.6846e-08 0.0007 3.6849e-08 0 3.6963e-08 0 3.6966e-08 0.0007 3.6969e-08 0 3.7083e-08 0 3.7086e-08 0.0007 3.7089e-08 0 3.7203e-08 0 3.7206e-08 0.0007 3.7209e-08 0 3.7323e-08 0 3.7326e-08 0.0007 3.7329e-08 0 3.7443e-08 0 3.7446e-08 0.0007 3.7449e-08 0 3.7563e-08 0 3.7566e-08 0.0007 3.7569e-08 0 3.7683e-08 0 3.7686e-08 0.0007 3.7689e-08 0 3.7803e-08 0 3.7806e-08 0.0007 3.7809e-08 0 3.7923e-08 0 3.7926e-08 0.0007 3.7929e-08 0 3.8043e-08 0 3.8046e-08 0.0007 3.8049e-08 0 3.8163e-08 0 3.8166e-08 0.0007 3.8169e-08 0 3.8283e-08 0 3.8286e-08 0.0007 3.8289e-08 0 3.8403e-08 0 3.8406e-08 0.0007 3.8409e-08 0 3.8523e-08 0 3.8526e-08 0.0007 3.8529e-08 0 3.8643e-08 0 3.8646e-08 0.0007 3.8649e-08 0 3.8763e-08 0 3.8766e-08 0.0007 3.8769e-08 0 3.8883e-08 0 3.8886e-08 0.0007 3.8889e-08 0 3.9003e-08 0 3.9006e-08 0.0007 3.9009e-08 0 3.9123e-08 0 3.9126e-08 0.0007 3.9129e-08 0 3.9243e-08 0 3.9246e-08 0.0007 3.9249e-08 0 3.9363e-08 0 3.9366e-08 0.0007 3.9369e-08 0 3.9483e-08 0 3.9486e-08 0.0007 3.9489e-08 0 3.9603e-08 0 3.9606e-08 0.0007 3.9609e-08 0 3.9723e-08 0 3.9726e-08 0.0007 3.9729e-08 0 3.9843e-08 0 3.9846e-08 0.0007 3.9849e-08 0 3.9963e-08 0 3.9966e-08 0.0007 3.9969e-08 0 4.0083e-08 0 4.0086e-08 0.0007 4.0089e-08 0 4.0203e-08 0 4.0206e-08 0.0007 4.0209e-08 0 4.0323e-08 0 4.0326e-08 0.0007 4.0329e-08 0 4.0443e-08 0 4.0446e-08 0.0007 4.0449e-08 0 4.0563e-08 0 4.0566e-08 0.0007 4.0569e-08 0 4.0683e-08 0 4.0686e-08 0.0007 4.0689e-08 0 4.0803e-08 0 4.0806e-08 0.0007 4.0809e-08 0 4.0923e-08 0 4.0926e-08 0.0007 4.0929e-08 0 4.1043e-08 0 4.1046e-08 0.0007 4.1049e-08 0 4.1163e-08 0 4.1166e-08 0.0007 4.1169e-08 0 4.1283e-08 0 4.1286e-08 0.0007 4.1289e-08 0 4.1403e-08 0 4.1406e-08 0.0007 4.1409e-08 0 4.1523e-08 0 4.1526e-08 0.0007 4.1529e-08 0 4.1643e-08 0 4.1646e-08 0.0007 4.1649e-08 0 4.1763e-08 0 4.1766e-08 0.0007 4.1769e-08 0 4.1883e-08 0 4.1886e-08 0.0007 4.1889e-08 0 4.2003e-08 0 4.2006e-08 0.0007 4.2009e-08 0 4.2123e-08 0 4.2126e-08 0.0007 4.2129e-08 0 4.2243e-08 0 4.2246e-08 0.0007 4.2249e-08 0 4.2363e-08 0 4.2366e-08 0.0007 4.2369e-08 0 4.2483e-08 0 4.2486e-08 0.0007 4.2489e-08 0 4.2603e-08 0 4.2606e-08 0.0007 4.2609e-08 0 4.2723e-08 0 4.2726e-08 0.0007 4.2729e-08 0 4.2843e-08 0 4.2846e-08 0.0007 4.2849e-08 0 4.2963e-08 0 4.2966e-08 0.0007 4.2969e-08 0 4.3083e-08 0 4.3086e-08 0.0007 4.3089e-08 0 4.3203e-08 0 4.3206e-08 0.0007 4.3209e-08 0 4.3323e-08 0 4.3326e-08 0.0007 4.3329e-08 0 4.3443e-08 0 4.3446e-08 0.0007 4.3449e-08 0 4.3563e-08 0 4.3566e-08 0.0007 4.3569e-08 0 4.3683e-08 0 4.3686e-08 0.0007 4.3689e-08 0 4.3803e-08 0 4.3806e-08 0.0007 4.3809e-08 0 4.3923e-08 0 4.3926e-08 0.0007 4.3929e-08 0 4.4043e-08 0 4.4046e-08 0.0007 4.4049e-08 0 4.4163e-08 0 4.4166e-08 0.0007 4.4169e-08 0 4.4283e-08 0 4.4286e-08 0.0007 4.4289e-08 0 4.4403e-08 0 4.4406e-08 0.0007 4.4409e-08 0 4.4523e-08 0 4.4526e-08 0.0007 4.4529e-08 0 4.4643e-08 0 4.4646e-08 0.0007 4.4649e-08 0 4.4763e-08 0 4.4766e-08 0.0007 4.4769e-08 0 4.4883e-08 0 4.4886e-08 0.0007 4.4889e-08 0 4.5003e-08 0 4.5006e-08 0.0007 4.5009e-08 0 4.5123e-08 0 4.5126e-08 0.0007 4.5129e-08 0 4.5243e-08 0 4.5246e-08 0.0007 4.5249e-08 0 4.5363e-08 0 4.5366e-08 0.0007 4.5369e-08 0 4.5483e-08 0 4.5486e-08 0.0007 4.5489e-08 0 4.5603e-08 0 4.5606e-08 0.0007 4.5609e-08 0 4.5723e-08 0 4.5726e-08 0.0007 4.5729e-08 0 4.5843e-08 0 4.5846e-08 0.0007 4.5849e-08 0 4.5963e-08 0 4.5966e-08 0.0007 4.5969e-08 0 4.6083e-08 0 4.6086e-08 0.0007 4.6089e-08 0 4.6203e-08 0 4.6206e-08 0.0007 4.6209e-08 0 4.6323e-08 0 4.6326e-08 0.0007 4.6329e-08 0 4.6443e-08 0 4.6446e-08 0.0007 4.6449e-08 0 4.6563e-08 0 4.6566e-08 0.0007 4.6569e-08 0 4.6683e-08 0 4.6686e-08 0.0007 4.6689e-08 0 4.6803e-08 0 4.6806e-08 0.0007 4.6809e-08 0 4.6923e-08 0 4.6926e-08 0.0007 4.6929e-08 0 4.7043e-08 0 4.7046e-08 0.0007 4.7049e-08 0 4.7163e-08 0 4.7166e-08 0.0007 4.7169e-08 0 4.7283e-08 0 4.7286e-08 0.0007 4.7289e-08 0 4.7403e-08 0 4.7406e-08 0.0007 4.7409e-08 0 4.7523e-08 0 4.7526e-08 0.0007 4.7529e-08 0 4.7643e-08 0 4.7646e-08 0.0007 4.7649e-08 0 4.7763e-08 0 4.7766e-08 0.0007 4.7769e-08 0)
L_S2|A1 G1_2_RX _S2|A1  2.067833848e-12
L_S2|A2 _S2|A1 _S2|A2  4.135667696e-12
L_S2|A3 _S2|A3 _S2|AB  8.271335392e-12
L_S2|B1 IP2_2_OUT_RX _S2|B1  2.067833848e-12
L_S2|B2 _S2|B1 _S2|B2  4.135667696e-12
L_S2|B3 _S2|B3 _S2|AB  8.271335392e-12
L_S2|T1 T14 _S2|T1  2.067833848e-12
L_S2|T2 _S2|T1 _S2|T2  4.135667696e-12
L_S2|Q2 _S2|ABTQ _S2|Q1  4.135667696e-12
L_S2|Q1 _S2|Q1 S2  2.067833848e-12
IT15|T 0 T15  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0 2.4003e-08 0 2.4006e-08 0.0007 2.4009e-08 0 2.4123e-08 0 2.4126e-08 0.0007 2.4129e-08 0 2.4243e-08 0 2.4246e-08 0.0007 2.4249e-08 0 2.4363e-08 0 2.4366e-08 0.0007 2.4369e-08 0 2.4483e-08 0 2.4486e-08 0.0007 2.4489e-08 0 2.4603e-08 0 2.4606e-08 0.0007 2.4609e-08 0 2.4723e-08 0 2.4726e-08 0.0007 2.4729e-08 0 2.4843e-08 0 2.4846e-08 0.0007 2.4849e-08 0 2.4963e-08 0 2.4966e-08 0.0007 2.4969e-08 0 2.5083e-08 0 2.5086e-08 0.0007 2.5089e-08 0 2.5203e-08 0 2.5206e-08 0.0007 2.5209e-08 0 2.5323e-08 0 2.5326e-08 0.0007 2.5329e-08 0 2.5443e-08 0 2.5446e-08 0.0007 2.5449e-08 0 2.5563e-08 0 2.5566e-08 0.0007 2.5569e-08 0 2.5683e-08 0 2.5686e-08 0.0007 2.5689e-08 0 2.5803e-08 0 2.5806e-08 0.0007 2.5809e-08 0 2.5923e-08 0 2.5926e-08 0.0007 2.5929e-08 0 2.6043e-08 0 2.6046e-08 0.0007 2.6049e-08 0 2.6163e-08 0 2.6166e-08 0.0007 2.6169e-08 0 2.6283e-08 0 2.6286e-08 0.0007 2.6289e-08 0 2.6403e-08 0 2.6406e-08 0.0007 2.6409e-08 0 2.6523e-08 0 2.6526e-08 0.0007 2.6529e-08 0 2.6643e-08 0 2.6646e-08 0.0007 2.6649e-08 0 2.6763e-08 0 2.6766e-08 0.0007 2.6769e-08 0 2.6883e-08 0 2.6886e-08 0.0007 2.6889e-08 0 2.7003e-08 0 2.7006e-08 0.0007 2.7009e-08 0 2.7123e-08 0 2.7126e-08 0.0007 2.7129e-08 0 2.7243e-08 0 2.7246e-08 0.0007 2.7249e-08 0 2.7363e-08 0 2.7366e-08 0.0007 2.7369e-08 0 2.7483e-08 0 2.7486e-08 0.0007 2.7489e-08 0 2.7603e-08 0 2.7606e-08 0.0007 2.7609e-08 0 2.7723e-08 0 2.7726e-08 0.0007 2.7729e-08 0 2.7843e-08 0 2.7846e-08 0.0007 2.7849e-08 0 2.7963e-08 0 2.7966e-08 0.0007 2.7969e-08 0 2.8083e-08 0 2.8086e-08 0.0007 2.8089e-08 0 2.8203e-08 0 2.8206e-08 0.0007 2.8209e-08 0 2.8323e-08 0 2.8326e-08 0.0007 2.8329e-08 0 2.8443e-08 0 2.8446e-08 0.0007 2.8449e-08 0 2.8563e-08 0 2.8566e-08 0.0007 2.8569e-08 0 2.8683e-08 0 2.8686e-08 0.0007 2.8689e-08 0 2.8803e-08 0 2.8806e-08 0.0007 2.8809e-08 0 2.8923e-08 0 2.8926e-08 0.0007 2.8929e-08 0 2.9043e-08 0 2.9046e-08 0.0007 2.9049e-08 0 2.9163e-08 0 2.9166e-08 0.0007 2.9169e-08 0 2.9283e-08 0 2.9286e-08 0.0007 2.9289e-08 0 2.9403e-08 0 2.9406e-08 0.0007 2.9409e-08 0 2.9523e-08 0 2.9526e-08 0.0007 2.9529e-08 0 2.9643e-08 0 2.9646e-08 0.0007 2.9649e-08 0 2.9763e-08 0 2.9766e-08 0.0007 2.9769e-08 0 2.9883e-08 0 2.9886e-08 0.0007 2.9889e-08 0 3.0003e-08 0 3.0006e-08 0.0007 3.0009e-08 0 3.0123e-08 0 3.0126e-08 0.0007 3.0129e-08 0 3.0243e-08 0 3.0246e-08 0.0007 3.0249e-08 0 3.0363e-08 0 3.0366e-08 0.0007 3.0369e-08 0 3.0483e-08 0 3.0486e-08 0.0007 3.0489e-08 0 3.0603e-08 0 3.0606e-08 0.0007 3.0609e-08 0 3.0723e-08 0 3.0726e-08 0.0007 3.0729e-08 0 3.0843e-08 0 3.0846e-08 0.0007 3.0849e-08 0 3.0963e-08 0 3.0966e-08 0.0007 3.0969e-08 0 3.1083e-08 0 3.1086e-08 0.0007 3.1089e-08 0 3.1203e-08 0 3.1206e-08 0.0007 3.1209e-08 0 3.1323e-08 0 3.1326e-08 0.0007 3.1329e-08 0 3.1443e-08 0 3.1446e-08 0.0007 3.1449e-08 0 3.1563e-08 0 3.1566e-08 0.0007 3.1569e-08 0 3.1683e-08 0 3.1686e-08 0.0007 3.1689e-08 0 3.1803e-08 0 3.1806e-08 0.0007 3.1809e-08 0 3.1923e-08 0 3.1926e-08 0.0007 3.1929e-08 0 3.2043e-08 0 3.2046e-08 0.0007 3.2049e-08 0 3.2163e-08 0 3.2166e-08 0.0007 3.2169e-08 0 3.2283e-08 0 3.2286e-08 0.0007 3.2289e-08 0 3.2403e-08 0 3.2406e-08 0.0007 3.2409e-08 0 3.2523e-08 0 3.2526e-08 0.0007 3.2529e-08 0 3.2643e-08 0 3.2646e-08 0.0007 3.2649e-08 0 3.2763e-08 0 3.2766e-08 0.0007 3.2769e-08 0 3.2883e-08 0 3.2886e-08 0.0007 3.2889e-08 0 3.3003e-08 0 3.3006e-08 0.0007 3.3009e-08 0 3.3123e-08 0 3.3126e-08 0.0007 3.3129e-08 0 3.3243e-08 0 3.3246e-08 0.0007 3.3249e-08 0 3.3363e-08 0 3.3366e-08 0.0007 3.3369e-08 0 3.3483e-08 0 3.3486e-08 0.0007 3.3489e-08 0 3.3603e-08 0 3.3606e-08 0.0007 3.3609e-08 0 3.3723e-08 0 3.3726e-08 0.0007 3.3729e-08 0 3.3843e-08 0 3.3846e-08 0.0007 3.3849e-08 0 3.3963e-08 0 3.3966e-08 0.0007 3.3969e-08 0 3.4083e-08 0 3.4086e-08 0.0007 3.4089e-08 0 3.4203e-08 0 3.4206e-08 0.0007 3.4209e-08 0 3.4323e-08 0 3.4326e-08 0.0007 3.4329e-08 0 3.4443e-08 0 3.4446e-08 0.0007 3.4449e-08 0 3.4563e-08 0 3.4566e-08 0.0007 3.4569e-08 0 3.4683e-08 0 3.4686e-08 0.0007 3.4689e-08 0 3.4803e-08 0 3.4806e-08 0.0007 3.4809e-08 0 3.4923e-08 0 3.4926e-08 0.0007 3.4929e-08 0 3.5043e-08 0 3.5046e-08 0.0007 3.5049e-08 0 3.5163e-08 0 3.5166e-08 0.0007 3.5169e-08 0 3.5283e-08 0 3.5286e-08 0.0007 3.5289e-08 0 3.5403e-08 0 3.5406e-08 0.0007 3.5409e-08 0 3.5523e-08 0 3.5526e-08 0.0007 3.5529e-08 0 3.5643e-08 0 3.5646e-08 0.0007 3.5649e-08 0 3.5763e-08 0 3.5766e-08 0.0007 3.5769e-08 0 3.5883e-08 0 3.5886e-08 0.0007 3.5889e-08 0 3.6003e-08 0 3.6006e-08 0.0007 3.6009e-08 0 3.6123e-08 0 3.6126e-08 0.0007 3.6129e-08 0 3.6243e-08 0 3.6246e-08 0.0007 3.6249e-08 0 3.6363e-08 0 3.6366e-08 0.0007 3.6369e-08 0 3.6483e-08 0 3.6486e-08 0.0007 3.6489e-08 0 3.6603e-08 0 3.6606e-08 0.0007 3.6609e-08 0 3.6723e-08 0 3.6726e-08 0.0007 3.6729e-08 0 3.6843e-08 0 3.6846e-08 0.0007 3.6849e-08 0 3.6963e-08 0 3.6966e-08 0.0007 3.6969e-08 0 3.7083e-08 0 3.7086e-08 0.0007 3.7089e-08 0 3.7203e-08 0 3.7206e-08 0.0007 3.7209e-08 0 3.7323e-08 0 3.7326e-08 0.0007 3.7329e-08 0 3.7443e-08 0 3.7446e-08 0.0007 3.7449e-08 0 3.7563e-08 0 3.7566e-08 0.0007 3.7569e-08 0 3.7683e-08 0 3.7686e-08 0.0007 3.7689e-08 0 3.7803e-08 0 3.7806e-08 0.0007 3.7809e-08 0 3.7923e-08 0 3.7926e-08 0.0007 3.7929e-08 0 3.8043e-08 0 3.8046e-08 0.0007 3.8049e-08 0 3.8163e-08 0 3.8166e-08 0.0007 3.8169e-08 0 3.8283e-08 0 3.8286e-08 0.0007 3.8289e-08 0 3.8403e-08 0 3.8406e-08 0.0007 3.8409e-08 0 3.8523e-08 0 3.8526e-08 0.0007 3.8529e-08 0 3.8643e-08 0 3.8646e-08 0.0007 3.8649e-08 0 3.8763e-08 0 3.8766e-08 0.0007 3.8769e-08 0 3.8883e-08 0 3.8886e-08 0.0007 3.8889e-08 0 3.9003e-08 0 3.9006e-08 0.0007 3.9009e-08 0 3.9123e-08 0 3.9126e-08 0.0007 3.9129e-08 0 3.9243e-08 0 3.9246e-08 0.0007 3.9249e-08 0 3.9363e-08 0 3.9366e-08 0.0007 3.9369e-08 0 3.9483e-08 0 3.9486e-08 0.0007 3.9489e-08 0 3.9603e-08 0 3.9606e-08 0.0007 3.9609e-08 0 3.9723e-08 0 3.9726e-08 0.0007 3.9729e-08 0 3.9843e-08 0 3.9846e-08 0.0007 3.9849e-08 0 3.9963e-08 0 3.9966e-08 0.0007 3.9969e-08 0 4.0083e-08 0 4.0086e-08 0.0007 4.0089e-08 0 4.0203e-08 0 4.0206e-08 0.0007 4.0209e-08 0 4.0323e-08 0 4.0326e-08 0.0007 4.0329e-08 0 4.0443e-08 0 4.0446e-08 0.0007 4.0449e-08 0 4.0563e-08 0 4.0566e-08 0.0007 4.0569e-08 0 4.0683e-08 0 4.0686e-08 0.0007 4.0689e-08 0 4.0803e-08 0 4.0806e-08 0.0007 4.0809e-08 0 4.0923e-08 0 4.0926e-08 0.0007 4.0929e-08 0 4.1043e-08 0 4.1046e-08 0.0007 4.1049e-08 0 4.1163e-08 0 4.1166e-08 0.0007 4.1169e-08 0 4.1283e-08 0 4.1286e-08 0.0007 4.1289e-08 0 4.1403e-08 0 4.1406e-08 0.0007 4.1409e-08 0 4.1523e-08 0 4.1526e-08 0.0007 4.1529e-08 0 4.1643e-08 0 4.1646e-08 0.0007 4.1649e-08 0 4.1763e-08 0 4.1766e-08 0.0007 4.1769e-08 0 4.1883e-08 0 4.1886e-08 0.0007 4.1889e-08 0 4.2003e-08 0 4.2006e-08 0.0007 4.2009e-08 0 4.2123e-08 0 4.2126e-08 0.0007 4.2129e-08 0 4.2243e-08 0 4.2246e-08 0.0007 4.2249e-08 0 4.2363e-08 0 4.2366e-08 0.0007 4.2369e-08 0 4.2483e-08 0 4.2486e-08 0.0007 4.2489e-08 0 4.2603e-08 0 4.2606e-08 0.0007 4.2609e-08 0 4.2723e-08 0 4.2726e-08 0.0007 4.2729e-08 0 4.2843e-08 0 4.2846e-08 0.0007 4.2849e-08 0 4.2963e-08 0 4.2966e-08 0.0007 4.2969e-08 0 4.3083e-08 0 4.3086e-08 0.0007 4.3089e-08 0 4.3203e-08 0 4.3206e-08 0.0007 4.3209e-08 0 4.3323e-08 0 4.3326e-08 0.0007 4.3329e-08 0 4.3443e-08 0 4.3446e-08 0.0007 4.3449e-08 0 4.3563e-08 0 4.3566e-08 0.0007 4.3569e-08 0 4.3683e-08 0 4.3686e-08 0.0007 4.3689e-08 0 4.3803e-08 0 4.3806e-08 0.0007 4.3809e-08 0 4.3923e-08 0 4.3926e-08 0.0007 4.3929e-08 0 4.4043e-08 0 4.4046e-08 0.0007 4.4049e-08 0 4.4163e-08 0 4.4166e-08 0.0007 4.4169e-08 0 4.4283e-08 0 4.4286e-08 0.0007 4.4289e-08 0 4.4403e-08 0 4.4406e-08 0.0007 4.4409e-08 0 4.4523e-08 0 4.4526e-08 0.0007 4.4529e-08 0 4.4643e-08 0 4.4646e-08 0.0007 4.4649e-08 0 4.4763e-08 0 4.4766e-08 0.0007 4.4769e-08 0 4.4883e-08 0 4.4886e-08 0.0007 4.4889e-08 0 4.5003e-08 0 4.5006e-08 0.0007 4.5009e-08 0 4.5123e-08 0 4.5126e-08 0.0007 4.5129e-08 0 4.5243e-08 0 4.5246e-08 0.0007 4.5249e-08 0 4.5363e-08 0 4.5366e-08 0.0007 4.5369e-08 0 4.5483e-08 0 4.5486e-08 0.0007 4.5489e-08 0 4.5603e-08 0 4.5606e-08 0.0007 4.5609e-08 0 4.5723e-08 0 4.5726e-08 0.0007 4.5729e-08 0 4.5843e-08 0 4.5846e-08 0.0007 4.5849e-08 0 4.5963e-08 0 4.5966e-08 0.0007 4.5969e-08 0 4.6083e-08 0 4.6086e-08 0.0007 4.6089e-08 0 4.6203e-08 0 4.6206e-08 0.0007 4.6209e-08 0 4.6323e-08 0 4.6326e-08 0.0007 4.6329e-08 0 4.6443e-08 0 4.6446e-08 0.0007 4.6449e-08 0 4.6563e-08 0 4.6566e-08 0.0007 4.6569e-08 0 4.6683e-08 0 4.6686e-08 0.0007 4.6689e-08 0 4.6803e-08 0 4.6806e-08 0.0007 4.6809e-08 0 4.6923e-08 0 4.6926e-08 0.0007 4.6929e-08 0 4.7043e-08 0 4.7046e-08 0.0007 4.7049e-08 0 4.7163e-08 0 4.7166e-08 0.0007 4.7169e-08 0 4.7283e-08 0 4.7286e-08 0.0007 4.7289e-08 0 4.7403e-08 0 4.7406e-08 0.0007 4.7409e-08 0 4.7523e-08 0 4.7526e-08 0.0007 4.7529e-08 0 4.7643e-08 0 4.7646e-08 0.0007 4.7649e-08 0 4.7763e-08 0 4.7766e-08 0.0007 4.7769e-08 0)
L_S3|A1 G2_2_RX _S3|A1  2.067833848e-12
L_S3|A2 _S3|A1 _S3|A2  4.135667696e-12
L_S3|A3 _S3|A3 _S3|AB  8.271335392e-12
L_S3|B1 IP3_2_OUT_RX _S3|B1  2.067833848e-12
L_S3|B2 _S3|B1 _S3|B2  4.135667696e-12
L_S3|B3 _S3|B3 _S3|AB  8.271335392e-12
L_S3|T1 T15 _S3|T1  2.067833848e-12
L_S3|T2 _S3|T1 _S3|T2  4.135667696e-12
L_S3|Q2 _S3|ABTQ _S3|Q1  4.135667696e-12
L_S3|Q1 _S3|Q1 S3  2.067833848e-12
IT16|T 0 T16  PWL(0 0 3e-12 0 6e-12 0.0007 9e-12 0 1.23e-10 0 1.26e-10 0.0007 1.29e-10 0 2.43e-10 0 2.46e-10 0.0007 2.49e-10 0 3.63e-10 0 3.66e-10 0.0007 3.69e-10 0 4.83e-10 0 4.86e-10 0.0007 4.89e-10 0 6.03e-10 0 6.06e-10 0.0007 6.09e-10 0 7.23e-10 0 7.26e-10 0.0007 7.29e-10 0 8.43e-10 0 8.46e-10 0.0007 8.49e-10 0 9.63e-10 0 9.66e-10 0.0007 9.69e-10 0 1.083e-09 0 1.086e-09 0.0007 1.089e-09 0 1.203e-09 0 1.206e-09 0.0007 1.209e-09 0 1.323e-09 0 1.326e-09 0.0007 1.329e-09 0 1.443e-09 0 1.446e-09 0.0007 1.449e-09 0 1.563e-09 0 1.566e-09 0.0007 1.569e-09 0 1.683e-09 0 1.686e-09 0.0007 1.689e-09 0 1.803e-09 0 1.806e-09 0.0007 1.809e-09 0 1.923e-09 0 1.926e-09 0.0007 1.929e-09 0 2.043e-09 0 2.046e-09 0.0007 2.049e-09 0 2.163e-09 0 2.166e-09 0.0007 2.169e-09 0 2.283e-09 0 2.286e-09 0.0007 2.289e-09 0 2.403e-09 0 2.406e-09 0.0007 2.409e-09 0 2.523e-09 0 2.526e-09 0.0007 2.529e-09 0 2.643e-09 0 2.646e-09 0.0007 2.649e-09 0 2.763e-09 0 2.766e-09 0.0007 2.769e-09 0 2.883e-09 0 2.886e-09 0.0007 2.889e-09 0 3.003e-09 0 3.006e-09 0.0007 3.009e-09 0 3.123e-09 0 3.126e-09 0.0007 3.129e-09 0 3.243e-09 0 3.246e-09 0.0007 3.249e-09 0 3.363e-09 0 3.366e-09 0.0007 3.369e-09 0 3.483e-09 0 3.486e-09 0.0007 3.489e-09 0 3.603e-09 0 3.606e-09 0.0007 3.609e-09 0 3.723e-09 0 3.726e-09 0.0007 3.729e-09 0 3.843e-09 0 3.846e-09 0.0007 3.849e-09 0 3.963e-09 0 3.966e-09 0.0007 3.969e-09 0 4.083e-09 0 4.086e-09 0.0007 4.089e-09 0 4.203e-09 0 4.206e-09 0.0007 4.209e-09 0 4.323e-09 0 4.326e-09 0.0007 4.329e-09 0 4.443e-09 0 4.446e-09 0.0007 4.449e-09 0 4.563e-09 0 4.566e-09 0.0007 4.569e-09 0 4.683e-09 0 4.686e-09 0.0007 4.689e-09 0 4.803e-09 0 4.806e-09 0.0007 4.809e-09 0 4.923e-09 0 4.926e-09 0.0007 4.929e-09 0 5.043e-09 0 5.046e-09 0.0007 5.049e-09 0 5.163e-09 0 5.166e-09 0.0007 5.169e-09 0 5.283e-09 0 5.286e-09 0.0007 5.289e-09 0 5.403e-09 0 5.406e-09 0.0007 5.409e-09 0 5.523e-09 0 5.526e-09 0.0007 5.529e-09 0 5.643e-09 0 5.646e-09 0.0007 5.649e-09 0 5.763e-09 0 5.766e-09 0.0007 5.769e-09 0 5.883e-09 0 5.886e-09 0.0007 5.889e-09 0 6.003e-09 0 6.006e-09 0.0007 6.009e-09 0 6.123e-09 0 6.126e-09 0.0007 6.129e-09 0 6.243e-09 0 6.246e-09 0.0007 6.249e-09 0 6.363e-09 0 6.366e-09 0.0007 6.369e-09 0 6.483e-09 0 6.486e-09 0.0007 6.489e-09 0 6.603e-09 0 6.606e-09 0.0007 6.609e-09 0 6.723e-09 0 6.726e-09 0.0007 6.729e-09 0 6.843e-09 0 6.846e-09 0.0007 6.849e-09 0 6.963e-09 0 6.966e-09 0.0007 6.969e-09 0 7.083e-09 0 7.086e-09 0.0007 7.089e-09 0 7.203e-09 0 7.206e-09 0.0007 7.209e-09 0 7.323e-09 0 7.326e-09 0.0007 7.329e-09 0 7.443e-09 0 7.446e-09 0.0007 7.449e-09 0 7.563e-09 0 7.566e-09 0.0007 7.569e-09 0 7.683e-09 0 7.686e-09 0.0007 7.689e-09 0 7.803e-09 0 7.806e-09 0.0007 7.809e-09 0 7.923e-09 0 7.926e-09 0.0007 7.929e-09 0 8.043e-09 0 8.046e-09 0.0007 8.049e-09 0 8.163e-09 0 8.166e-09 0.0007 8.169e-09 0 8.283e-09 0 8.286e-09 0.0007 8.289e-09 0 8.403e-09 0 8.406e-09 0.0007 8.409e-09 0 8.523e-09 0 8.526e-09 0.0007 8.529e-09 0 8.643e-09 0 8.646e-09 0.0007 8.649e-09 0 8.763e-09 0 8.766e-09 0.0007 8.769e-09 0 8.883e-09 0 8.886e-09 0.0007 8.889e-09 0 9.003e-09 0 9.006e-09 0.0007 9.009e-09 0 9.123e-09 0 9.126e-09 0.0007 9.129e-09 0 9.243e-09 0 9.246e-09 0.0007 9.249e-09 0 9.363e-09 0 9.366e-09 0.0007 9.369e-09 0 9.483e-09 0 9.486e-09 0.0007 9.489e-09 0 9.603e-09 0 9.606e-09 0.0007 9.609e-09 0 9.723e-09 0 9.726e-09 0.0007 9.729e-09 0 9.843e-09 0 9.846e-09 0.0007 9.849e-09 0 9.963e-09 0 9.966e-09 0.0007 9.969e-09 0 1.0083e-08 0 1.0086e-08 0.0007 1.0089e-08 0 1.0203e-08 0 1.0206e-08 0.0007 1.0209e-08 0 1.0323e-08 0 1.0326e-08 0.0007 1.0329e-08 0 1.0443e-08 0 1.0446e-08 0.0007 1.0449e-08 0 1.0563e-08 0 1.0566e-08 0.0007 1.0569e-08 0 1.0683e-08 0 1.0686e-08 0.0007 1.0689e-08 0 1.0803e-08 0 1.0806e-08 0.0007 1.0809e-08 0 1.0923e-08 0 1.0926e-08 0.0007 1.0929e-08 0 1.1043e-08 0 1.1046e-08 0.0007 1.1049e-08 0 1.1163e-08 0 1.1166e-08 0.0007 1.1169e-08 0 1.1283e-08 0 1.1286e-08 0.0007 1.1289e-08 0 1.1403e-08 0 1.1406e-08 0.0007 1.1409e-08 0 1.1523e-08 0 1.1526e-08 0.0007 1.1529e-08 0 1.1643e-08 0 1.1646e-08 0.0007 1.1649e-08 0 1.1763e-08 0 1.1766e-08 0.0007 1.1769e-08 0 1.1883e-08 0 1.1886e-08 0.0007 1.1889e-08 0 1.2003e-08 0 1.2006e-08 0.0007 1.2009e-08 0 1.2123e-08 0 1.2126e-08 0.0007 1.2129e-08 0 1.2243e-08 0 1.2246e-08 0.0007 1.2249e-08 0 1.2363e-08 0 1.2366e-08 0.0007 1.2369e-08 0 1.2483e-08 0 1.2486e-08 0.0007 1.2489e-08 0 1.2603e-08 0 1.2606e-08 0.0007 1.2609e-08 0 1.2723e-08 0 1.2726e-08 0.0007 1.2729e-08 0 1.2843e-08 0 1.2846e-08 0.0007 1.2849e-08 0 1.2963e-08 0 1.2966e-08 0.0007 1.2969e-08 0 1.3083e-08 0 1.3086e-08 0.0007 1.3089e-08 0 1.3203e-08 0 1.3206e-08 0.0007 1.3209e-08 0 1.3323e-08 0 1.3326e-08 0.0007 1.3329e-08 0 1.3443e-08 0 1.3446e-08 0.0007 1.3449e-08 0 1.3563e-08 0 1.3566e-08 0.0007 1.3569e-08 0 1.3683e-08 0 1.3686e-08 0.0007 1.3689e-08 0 1.3803e-08 0 1.3806e-08 0.0007 1.3809e-08 0 1.3923e-08 0 1.3926e-08 0.0007 1.3929e-08 0 1.4043e-08 0 1.4046e-08 0.0007 1.4049e-08 0 1.4163e-08 0 1.4166e-08 0.0007 1.4169e-08 0 1.4283e-08 0 1.4286e-08 0.0007 1.4289e-08 0 1.4403e-08 0 1.4406e-08 0.0007 1.4409e-08 0 1.4523e-08 0 1.4526e-08 0.0007 1.4529e-08 0 1.4643e-08 0 1.4646e-08 0.0007 1.4649e-08 0 1.4763e-08 0 1.4766e-08 0.0007 1.4769e-08 0 1.4883e-08 0 1.4886e-08 0.0007 1.4889e-08 0 1.5003e-08 0 1.5006e-08 0.0007 1.5009e-08 0 1.5123e-08 0 1.5126e-08 0.0007 1.5129e-08 0 1.5243e-08 0 1.5246e-08 0.0007 1.5249e-08 0 1.5363e-08 0 1.5366e-08 0.0007 1.5369e-08 0 1.5483e-08 0 1.5486e-08 0.0007 1.5489e-08 0 1.5603e-08 0 1.5606e-08 0.0007 1.5609e-08 0 1.5723e-08 0 1.5726e-08 0.0007 1.5729e-08 0 1.5843e-08 0 1.5846e-08 0.0007 1.5849e-08 0 1.5963e-08 0 1.5966e-08 0.0007 1.5969e-08 0 1.6083e-08 0 1.6086e-08 0.0007 1.6089e-08 0 1.6203e-08 0 1.6206e-08 0.0007 1.6209e-08 0 1.6323e-08 0 1.6326e-08 0.0007 1.6329e-08 0 1.6443e-08 0 1.6446e-08 0.0007 1.6449e-08 0 1.6563e-08 0 1.6566e-08 0.0007 1.6569e-08 0 1.6683e-08 0 1.6686e-08 0.0007 1.6689e-08 0 1.6803e-08 0 1.6806e-08 0.0007 1.6809e-08 0 1.6923e-08 0 1.6926e-08 0.0007 1.6929e-08 0 1.7043e-08 0 1.7046e-08 0.0007 1.7049e-08 0 1.7163e-08 0 1.7166e-08 0.0007 1.7169e-08 0 1.7283e-08 0 1.7286e-08 0.0007 1.7289e-08 0 1.7403e-08 0 1.7406e-08 0.0007 1.7409e-08 0 1.7523e-08 0 1.7526e-08 0.0007 1.7529e-08 0 1.7643e-08 0 1.7646e-08 0.0007 1.7649e-08 0 1.7763e-08 0 1.7766e-08 0.0007 1.7769e-08 0 1.7883e-08 0 1.7886e-08 0.0007 1.7889e-08 0 1.8003e-08 0 1.8006e-08 0.0007 1.8009e-08 0 1.8123e-08 0 1.8126e-08 0.0007 1.8129e-08 0 1.8243e-08 0 1.8246e-08 0.0007 1.8249e-08 0 1.8363e-08 0 1.8366e-08 0.0007 1.8369e-08 0 1.8483e-08 0 1.8486e-08 0.0007 1.8489e-08 0 1.8603e-08 0 1.8606e-08 0.0007 1.8609e-08 0 1.8723e-08 0 1.8726e-08 0.0007 1.8729e-08 0 1.8843e-08 0 1.8846e-08 0.0007 1.8849e-08 0 1.8963e-08 0 1.8966e-08 0.0007 1.8969e-08 0 1.9083e-08 0 1.9086e-08 0.0007 1.9089e-08 0 1.9203e-08 0 1.9206e-08 0.0007 1.9209e-08 0 1.9323e-08 0 1.9326e-08 0.0007 1.9329e-08 0 1.9443e-08 0 1.9446e-08 0.0007 1.9449e-08 0 1.9563e-08 0 1.9566e-08 0.0007 1.9569e-08 0 1.9683e-08 0 1.9686e-08 0.0007 1.9689e-08 0 1.9803e-08 0 1.9806e-08 0.0007 1.9809e-08 0 1.9923e-08 0 1.9926e-08 0.0007 1.9929e-08 0 2.0043e-08 0 2.0046e-08 0.0007 2.0049e-08 0 2.0163e-08 0 2.0166e-08 0.0007 2.0169e-08 0 2.0283e-08 0 2.0286e-08 0.0007 2.0289e-08 0 2.0403e-08 0 2.0406e-08 0.0007 2.0409e-08 0 2.0523e-08 0 2.0526e-08 0.0007 2.0529e-08 0 2.0643e-08 0 2.0646e-08 0.0007 2.0649e-08 0 2.0763e-08 0 2.0766e-08 0.0007 2.0769e-08 0 2.0883e-08 0 2.0886e-08 0.0007 2.0889e-08 0 2.1003e-08 0 2.1006e-08 0.0007 2.1009e-08 0 2.1123e-08 0 2.1126e-08 0.0007 2.1129e-08 0 2.1243e-08 0 2.1246e-08 0.0007 2.1249e-08 0 2.1363e-08 0 2.1366e-08 0.0007 2.1369e-08 0 2.1483e-08 0 2.1486e-08 0.0007 2.1489e-08 0 2.1603e-08 0 2.1606e-08 0.0007 2.1609e-08 0 2.1723e-08 0 2.1726e-08 0.0007 2.1729e-08 0 2.1843e-08 0 2.1846e-08 0.0007 2.1849e-08 0 2.1963e-08 0 2.1966e-08 0.0007 2.1969e-08 0 2.2083e-08 0 2.2086e-08 0.0007 2.2089e-08 0 2.2203e-08 0 2.2206e-08 0.0007 2.2209e-08 0 2.2323e-08 0 2.2326e-08 0.0007 2.2329e-08 0 2.2443e-08 0 2.2446e-08 0.0007 2.2449e-08 0 2.2563e-08 0 2.2566e-08 0.0007 2.2569e-08 0 2.2683e-08 0 2.2686e-08 0.0007 2.2689e-08 0 2.2803e-08 0 2.2806e-08 0.0007 2.2809e-08 0 2.2923e-08 0 2.2926e-08 0.0007 2.2929e-08 0 2.3043e-08 0 2.3046e-08 0.0007 2.3049e-08 0 2.3163e-08 0 2.3166e-08 0.0007 2.3169e-08 0 2.3283e-08 0 2.3286e-08 0.0007 2.3289e-08 0 2.3403e-08 0 2.3406e-08 0.0007 2.3409e-08 0 2.3523e-08 0 2.3526e-08 0.0007 2.3529e-08 0 2.3643e-08 0 2.3646e-08 0.0007 2.3649e-08 0 2.3763e-08 0 2.3766e-08 0.0007 2.3769e-08 0 2.3883e-08 0 2.3886e-08 0.0007 2.3889e-08 0 2.4003e-08 0 2.4006e-08 0.0007 2.4009e-08 0 2.4123e-08 0 2.4126e-08 0.0007 2.4129e-08 0 2.4243e-08 0 2.4246e-08 0.0007 2.4249e-08 0 2.4363e-08 0 2.4366e-08 0.0007 2.4369e-08 0 2.4483e-08 0 2.4486e-08 0.0007 2.4489e-08 0 2.4603e-08 0 2.4606e-08 0.0007 2.4609e-08 0 2.4723e-08 0 2.4726e-08 0.0007 2.4729e-08 0 2.4843e-08 0 2.4846e-08 0.0007 2.4849e-08 0 2.4963e-08 0 2.4966e-08 0.0007 2.4969e-08 0 2.5083e-08 0 2.5086e-08 0.0007 2.5089e-08 0 2.5203e-08 0 2.5206e-08 0.0007 2.5209e-08 0 2.5323e-08 0 2.5326e-08 0.0007 2.5329e-08 0 2.5443e-08 0 2.5446e-08 0.0007 2.5449e-08 0 2.5563e-08 0 2.5566e-08 0.0007 2.5569e-08 0 2.5683e-08 0 2.5686e-08 0.0007 2.5689e-08 0 2.5803e-08 0 2.5806e-08 0.0007 2.5809e-08 0 2.5923e-08 0 2.5926e-08 0.0007 2.5929e-08 0 2.6043e-08 0 2.6046e-08 0.0007 2.6049e-08 0 2.6163e-08 0 2.6166e-08 0.0007 2.6169e-08 0 2.6283e-08 0 2.6286e-08 0.0007 2.6289e-08 0 2.6403e-08 0 2.6406e-08 0.0007 2.6409e-08 0 2.6523e-08 0 2.6526e-08 0.0007 2.6529e-08 0 2.6643e-08 0 2.6646e-08 0.0007 2.6649e-08 0 2.6763e-08 0 2.6766e-08 0.0007 2.6769e-08 0 2.6883e-08 0 2.6886e-08 0.0007 2.6889e-08 0 2.7003e-08 0 2.7006e-08 0.0007 2.7009e-08 0 2.7123e-08 0 2.7126e-08 0.0007 2.7129e-08 0 2.7243e-08 0 2.7246e-08 0.0007 2.7249e-08 0 2.7363e-08 0 2.7366e-08 0.0007 2.7369e-08 0 2.7483e-08 0 2.7486e-08 0.0007 2.7489e-08 0 2.7603e-08 0 2.7606e-08 0.0007 2.7609e-08 0 2.7723e-08 0 2.7726e-08 0.0007 2.7729e-08 0 2.7843e-08 0 2.7846e-08 0.0007 2.7849e-08 0 2.7963e-08 0 2.7966e-08 0.0007 2.7969e-08 0 2.8083e-08 0 2.8086e-08 0.0007 2.8089e-08 0 2.8203e-08 0 2.8206e-08 0.0007 2.8209e-08 0 2.8323e-08 0 2.8326e-08 0.0007 2.8329e-08 0 2.8443e-08 0 2.8446e-08 0.0007 2.8449e-08 0 2.8563e-08 0 2.8566e-08 0.0007 2.8569e-08 0 2.8683e-08 0 2.8686e-08 0.0007 2.8689e-08 0 2.8803e-08 0 2.8806e-08 0.0007 2.8809e-08 0 2.8923e-08 0 2.8926e-08 0.0007 2.8929e-08 0 2.9043e-08 0 2.9046e-08 0.0007 2.9049e-08 0 2.9163e-08 0 2.9166e-08 0.0007 2.9169e-08 0 2.9283e-08 0 2.9286e-08 0.0007 2.9289e-08 0 2.9403e-08 0 2.9406e-08 0.0007 2.9409e-08 0 2.9523e-08 0 2.9526e-08 0.0007 2.9529e-08 0 2.9643e-08 0 2.9646e-08 0.0007 2.9649e-08 0 2.9763e-08 0 2.9766e-08 0.0007 2.9769e-08 0 2.9883e-08 0 2.9886e-08 0.0007 2.9889e-08 0 3.0003e-08 0 3.0006e-08 0.0007 3.0009e-08 0 3.0123e-08 0 3.0126e-08 0.0007 3.0129e-08 0 3.0243e-08 0 3.0246e-08 0.0007 3.0249e-08 0 3.0363e-08 0 3.0366e-08 0.0007 3.0369e-08 0 3.0483e-08 0 3.0486e-08 0.0007 3.0489e-08 0 3.0603e-08 0 3.0606e-08 0.0007 3.0609e-08 0 3.0723e-08 0 3.0726e-08 0.0007 3.0729e-08 0 3.0843e-08 0 3.0846e-08 0.0007 3.0849e-08 0 3.0963e-08 0 3.0966e-08 0.0007 3.0969e-08 0 3.1083e-08 0 3.1086e-08 0.0007 3.1089e-08 0 3.1203e-08 0 3.1206e-08 0.0007 3.1209e-08 0 3.1323e-08 0 3.1326e-08 0.0007 3.1329e-08 0 3.1443e-08 0 3.1446e-08 0.0007 3.1449e-08 0 3.1563e-08 0 3.1566e-08 0.0007 3.1569e-08 0 3.1683e-08 0 3.1686e-08 0.0007 3.1689e-08 0 3.1803e-08 0 3.1806e-08 0.0007 3.1809e-08 0 3.1923e-08 0 3.1926e-08 0.0007 3.1929e-08 0 3.2043e-08 0 3.2046e-08 0.0007 3.2049e-08 0 3.2163e-08 0 3.2166e-08 0.0007 3.2169e-08 0 3.2283e-08 0 3.2286e-08 0.0007 3.2289e-08 0 3.2403e-08 0 3.2406e-08 0.0007 3.2409e-08 0 3.2523e-08 0 3.2526e-08 0.0007 3.2529e-08 0 3.2643e-08 0 3.2646e-08 0.0007 3.2649e-08 0 3.2763e-08 0 3.2766e-08 0.0007 3.2769e-08 0 3.2883e-08 0 3.2886e-08 0.0007 3.2889e-08 0 3.3003e-08 0 3.3006e-08 0.0007 3.3009e-08 0 3.3123e-08 0 3.3126e-08 0.0007 3.3129e-08 0 3.3243e-08 0 3.3246e-08 0.0007 3.3249e-08 0 3.3363e-08 0 3.3366e-08 0.0007 3.3369e-08 0 3.3483e-08 0 3.3486e-08 0.0007 3.3489e-08 0 3.3603e-08 0 3.3606e-08 0.0007 3.3609e-08 0 3.3723e-08 0 3.3726e-08 0.0007 3.3729e-08 0 3.3843e-08 0 3.3846e-08 0.0007 3.3849e-08 0 3.3963e-08 0 3.3966e-08 0.0007 3.3969e-08 0 3.4083e-08 0 3.4086e-08 0.0007 3.4089e-08 0 3.4203e-08 0 3.4206e-08 0.0007 3.4209e-08 0 3.4323e-08 0 3.4326e-08 0.0007 3.4329e-08 0 3.4443e-08 0 3.4446e-08 0.0007 3.4449e-08 0 3.4563e-08 0 3.4566e-08 0.0007 3.4569e-08 0 3.4683e-08 0 3.4686e-08 0.0007 3.4689e-08 0 3.4803e-08 0 3.4806e-08 0.0007 3.4809e-08 0 3.4923e-08 0 3.4926e-08 0.0007 3.4929e-08 0 3.5043e-08 0 3.5046e-08 0.0007 3.5049e-08 0 3.5163e-08 0 3.5166e-08 0.0007 3.5169e-08 0 3.5283e-08 0 3.5286e-08 0.0007 3.5289e-08 0 3.5403e-08 0 3.5406e-08 0.0007 3.5409e-08 0 3.5523e-08 0 3.5526e-08 0.0007 3.5529e-08 0 3.5643e-08 0 3.5646e-08 0.0007 3.5649e-08 0 3.5763e-08 0 3.5766e-08 0.0007 3.5769e-08 0 3.5883e-08 0 3.5886e-08 0.0007 3.5889e-08 0 3.6003e-08 0 3.6006e-08 0.0007 3.6009e-08 0 3.6123e-08 0 3.6126e-08 0.0007 3.6129e-08 0 3.6243e-08 0 3.6246e-08 0.0007 3.6249e-08 0 3.6363e-08 0 3.6366e-08 0.0007 3.6369e-08 0 3.6483e-08 0 3.6486e-08 0.0007 3.6489e-08 0 3.6603e-08 0 3.6606e-08 0.0007 3.6609e-08 0 3.6723e-08 0 3.6726e-08 0.0007 3.6729e-08 0 3.6843e-08 0 3.6846e-08 0.0007 3.6849e-08 0 3.6963e-08 0 3.6966e-08 0.0007 3.6969e-08 0 3.7083e-08 0 3.7086e-08 0.0007 3.7089e-08 0 3.7203e-08 0 3.7206e-08 0.0007 3.7209e-08 0 3.7323e-08 0 3.7326e-08 0.0007 3.7329e-08 0 3.7443e-08 0 3.7446e-08 0.0007 3.7449e-08 0 3.7563e-08 0 3.7566e-08 0.0007 3.7569e-08 0 3.7683e-08 0 3.7686e-08 0.0007 3.7689e-08 0 3.7803e-08 0 3.7806e-08 0.0007 3.7809e-08 0 3.7923e-08 0 3.7926e-08 0.0007 3.7929e-08 0 3.8043e-08 0 3.8046e-08 0.0007 3.8049e-08 0 3.8163e-08 0 3.8166e-08 0.0007 3.8169e-08 0 3.8283e-08 0 3.8286e-08 0.0007 3.8289e-08 0 3.8403e-08 0 3.8406e-08 0.0007 3.8409e-08 0 3.8523e-08 0 3.8526e-08 0.0007 3.8529e-08 0 3.8643e-08 0 3.8646e-08 0.0007 3.8649e-08 0 3.8763e-08 0 3.8766e-08 0.0007 3.8769e-08 0 3.8883e-08 0 3.8886e-08 0.0007 3.8889e-08 0 3.9003e-08 0 3.9006e-08 0.0007 3.9009e-08 0 3.9123e-08 0 3.9126e-08 0.0007 3.9129e-08 0 3.9243e-08 0 3.9246e-08 0.0007 3.9249e-08 0 3.9363e-08 0 3.9366e-08 0.0007 3.9369e-08 0 3.9483e-08 0 3.9486e-08 0.0007 3.9489e-08 0 3.9603e-08 0 3.9606e-08 0.0007 3.9609e-08 0 3.9723e-08 0 3.9726e-08 0.0007 3.9729e-08 0 3.9843e-08 0 3.9846e-08 0.0007 3.9849e-08 0 3.9963e-08 0 3.9966e-08 0.0007 3.9969e-08 0 4.0083e-08 0 4.0086e-08 0.0007 4.0089e-08 0 4.0203e-08 0 4.0206e-08 0.0007 4.0209e-08 0 4.0323e-08 0 4.0326e-08 0.0007 4.0329e-08 0 4.0443e-08 0 4.0446e-08 0.0007 4.0449e-08 0 4.0563e-08 0 4.0566e-08 0.0007 4.0569e-08 0 4.0683e-08 0 4.0686e-08 0.0007 4.0689e-08 0 4.0803e-08 0 4.0806e-08 0.0007 4.0809e-08 0 4.0923e-08 0 4.0926e-08 0.0007 4.0929e-08 0 4.1043e-08 0 4.1046e-08 0.0007 4.1049e-08 0 4.1163e-08 0 4.1166e-08 0.0007 4.1169e-08 0 4.1283e-08 0 4.1286e-08 0.0007 4.1289e-08 0 4.1403e-08 0 4.1406e-08 0.0007 4.1409e-08 0 4.1523e-08 0 4.1526e-08 0.0007 4.1529e-08 0 4.1643e-08 0 4.1646e-08 0.0007 4.1649e-08 0 4.1763e-08 0 4.1766e-08 0.0007 4.1769e-08 0 4.1883e-08 0 4.1886e-08 0.0007 4.1889e-08 0 4.2003e-08 0 4.2006e-08 0.0007 4.2009e-08 0 4.2123e-08 0 4.2126e-08 0.0007 4.2129e-08 0 4.2243e-08 0 4.2246e-08 0.0007 4.2249e-08 0 4.2363e-08 0 4.2366e-08 0.0007 4.2369e-08 0 4.2483e-08 0 4.2486e-08 0.0007 4.2489e-08 0 4.2603e-08 0 4.2606e-08 0.0007 4.2609e-08 0 4.2723e-08 0 4.2726e-08 0.0007 4.2729e-08 0 4.2843e-08 0 4.2846e-08 0.0007 4.2849e-08 0 4.2963e-08 0 4.2966e-08 0.0007 4.2969e-08 0 4.3083e-08 0 4.3086e-08 0.0007 4.3089e-08 0 4.3203e-08 0 4.3206e-08 0.0007 4.3209e-08 0 4.3323e-08 0 4.3326e-08 0.0007 4.3329e-08 0 4.3443e-08 0 4.3446e-08 0.0007 4.3449e-08 0 4.3563e-08 0 4.3566e-08 0.0007 4.3569e-08 0 4.3683e-08 0 4.3686e-08 0.0007 4.3689e-08 0 4.3803e-08 0 4.3806e-08 0.0007 4.3809e-08 0 4.3923e-08 0 4.3926e-08 0.0007 4.3929e-08 0 4.4043e-08 0 4.4046e-08 0.0007 4.4049e-08 0 4.4163e-08 0 4.4166e-08 0.0007 4.4169e-08 0 4.4283e-08 0 4.4286e-08 0.0007 4.4289e-08 0 4.4403e-08 0 4.4406e-08 0.0007 4.4409e-08 0 4.4523e-08 0 4.4526e-08 0.0007 4.4529e-08 0 4.4643e-08 0 4.4646e-08 0.0007 4.4649e-08 0 4.4763e-08 0 4.4766e-08 0.0007 4.4769e-08 0 4.4883e-08 0 4.4886e-08 0.0007 4.4889e-08 0 4.5003e-08 0 4.5006e-08 0.0007 4.5009e-08 0 4.5123e-08 0 4.5126e-08 0.0007 4.5129e-08 0 4.5243e-08 0 4.5246e-08 0.0007 4.5249e-08 0 4.5363e-08 0 4.5366e-08 0.0007 4.5369e-08 0 4.5483e-08 0 4.5486e-08 0.0007 4.5489e-08 0 4.5603e-08 0 4.5606e-08 0.0007 4.5609e-08 0 4.5723e-08 0 4.5726e-08 0.0007 4.5729e-08 0 4.5843e-08 0 4.5846e-08 0.0007 4.5849e-08 0 4.5963e-08 0 4.5966e-08 0.0007 4.5969e-08 0 4.6083e-08 0 4.6086e-08 0.0007 4.6089e-08 0 4.6203e-08 0 4.6206e-08 0.0007 4.6209e-08 0 4.6323e-08 0 4.6326e-08 0.0007 4.6329e-08 0 4.6443e-08 0 4.6446e-08 0.0007 4.6449e-08 0 4.6563e-08 0 4.6566e-08 0.0007 4.6569e-08 0 4.6683e-08 0 4.6686e-08 0.0007 4.6689e-08 0 4.6803e-08 0 4.6806e-08 0.0007 4.6809e-08 0 4.6923e-08 0 4.6926e-08 0.0007 4.6929e-08 0 4.7043e-08 0 4.7046e-08 0.0007 4.7049e-08 0 4.7163e-08 0 4.7166e-08 0.0007 4.7169e-08 0 4.7283e-08 0 4.7286e-08 0.0007 4.7289e-08 0 4.7403e-08 0 4.7406e-08 0.0007 4.7409e-08 0 4.7523e-08 0 4.7526e-08 0.0007 4.7529e-08 0 4.7643e-08 0 4.7646e-08 0.0007 4.7649e-08 0 4.7763e-08 0 4.7766e-08 0.0007 4.7769e-08 0)
L_S4|1 G3_2_RX _S4|A1  2.067833848e-12
L_S4|2 _S4|A1 _S4|A2  4.135667696e-12
L_S4|3 _S4|A3 _S4|A4  8.271335392e-12
L_S4|T T16 _S4|T1  2.067833848e-12
L_S4|4 _S4|T1 _S4|T2  4.135667696e-12
L_S4|5 _S4|A4 _S4|Q1  4.135667696e-12
L_S4|6 _S4|Q1 S4  2.067833848e-12
B_PTL_A0|_TX|1 _PTL_A0|_TX|1 _PTL_A0|_TX|2 JJMIT AREA=2.5
B_PTL_A0|_TX|2 _PTL_A0|_TX|4 _PTL_A0|_TX|5 JJMIT AREA=2.5
I_PTL_A0|_TX|B1 0 _PTL_A0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A0|_TX|B2 0 _PTL_A0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|3  1.684e-12
L_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|6  3.596e-12
L_PTL_A0|_TX|1 A0 _PTL_A0|_TX|1  2.063e-12
L_PTL_A0|_TX|2 _PTL_A0|_TX|1 _PTL_A0|_TX|4  4.123e-12
L_PTL_A0|_TX|3 _PTL_A0|_TX|4 _PTL_A0|_TX|7  2.193e-12
R_PTL_A0|_TX|D _PTL_A0|_TX|7 _PTL_A0|A_PTL  1.36
L_PTL_A0|_TX|P1 _PTL_A0|_TX|2 0  5.254e-13
L_PTL_A0|_TX|P2 _PTL_A0|_TX|5 0  5.141e-13
R_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|101  2.7439617672
R_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|104  2.7439617672
L_PTL_A0|_TX|RB1 _PTL_A0|_TX|101 0  1.550338398468e-12
L_PTL_A0|_TX|RB2 _PTL_A0|_TX|104 0  1.550338398468e-12
B_PTL_A0|_RX|1 _PTL_A0|_RX|1 _PTL_A0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A0|_RX|2 _PTL_A0|_RX|4 _PTL_A0|_RX|5 JJMIT AREA=2.0
B_PTL_A0|_RX|3 _PTL_A0|_RX|7 _PTL_A0|_RX|8 JJMIT AREA=2.5
I_PTL_A0|_RX|B1 0 _PTL_A0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|3  2.777e-12
I_PTL_A0|_RX|B2 0 _PTL_A0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|6  2.685e-12
I_PTL_A0|_RX|B3 0 _PTL_A0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|9  2.764e-12
L_PTL_A0|_RX|1 _PTL_A0|A_PTL _PTL_A0|_RX|1  1.346e-12
L_PTL_A0|_RX|2 _PTL_A0|_RX|1 _PTL_A0|_RX|4  6.348e-12
L_PTL_A0|_RX|3 _PTL_A0|_RX|4 _PTL_A0|_RX|7  5.197e-12
L_PTL_A0|_RX|4 _PTL_A0|_RX|7 A0_RX  2.058e-12
L_PTL_A0|_RX|P1 _PTL_A0|_RX|2 0  4.795e-13
L_PTL_A0|_RX|P2 _PTL_A0|_RX|5 0  5.431e-13
L_PTL_A0|_RX|P3 _PTL_A0|_RX|8 0  5.339e-13
R_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|101  4.225701121488
R_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|104  3.429952209
R_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|107  2.7439617672
L_PTL_A0|_RX|RB1 _PTL_A0|_RX|101 0  2.38752113364072e-12
L_PTL_A0|_RX|RB2 _PTL_A0|_RX|104 0  1.937922998085e-12
L_PTL_A0|_RX|RB3 _PTL_A0|_RX|107 0  1.550338398468e-12
B_PTL_B0|_TX|1 _PTL_B0|_TX|1 _PTL_B0|_TX|2 JJMIT AREA=2.5
B_PTL_B0|_TX|2 _PTL_B0|_TX|4 _PTL_B0|_TX|5 JJMIT AREA=2.5
I_PTL_B0|_TX|B1 0 _PTL_B0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B0|_TX|B2 0 _PTL_B0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|3  1.684e-12
L_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|6  3.596e-12
L_PTL_B0|_TX|1 B0 _PTL_B0|_TX|1  2.063e-12
L_PTL_B0|_TX|2 _PTL_B0|_TX|1 _PTL_B0|_TX|4  4.123e-12
L_PTL_B0|_TX|3 _PTL_B0|_TX|4 _PTL_B0|_TX|7  2.193e-12
R_PTL_B0|_TX|D _PTL_B0|_TX|7 _PTL_B0|A_PTL  1.36
L_PTL_B0|_TX|P1 _PTL_B0|_TX|2 0  5.254e-13
L_PTL_B0|_TX|P2 _PTL_B0|_TX|5 0  5.141e-13
R_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|101  2.7439617672
R_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|104  2.7439617672
L_PTL_B0|_TX|RB1 _PTL_B0|_TX|101 0  1.550338398468e-12
L_PTL_B0|_TX|RB2 _PTL_B0|_TX|104 0  1.550338398468e-12
B_PTL_B0|_RX|1 _PTL_B0|_RX|1 _PTL_B0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B0|_RX|2 _PTL_B0|_RX|4 _PTL_B0|_RX|5 JJMIT AREA=2.0
B_PTL_B0|_RX|3 _PTL_B0|_RX|7 _PTL_B0|_RX|8 JJMIT AREA=2.5
I_PTL_B0|_RX|B1 0 _PTL_B0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|3  2.777e-12
I_PTL_B0|_RX|B2 0 _PTL_B0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|6  2.685e-12
I_PTL_B0|_RX|B3 0 _PTL_B0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|9  2.764e-12
L_PTL_B0|_RX|1 _PTL_B0|A_PTL _PTL_B0|_RX|1  1.346e-12
L_PTL_B0|_RX|2 _PTL_B0|_RX|1 _PTL_B0|_RX|4  6.348e-12
L_PTL_B0|_RX|3 _PTL_B0|_RX|4 _PTL_B0|_RX|7  5.197e-12
L_PTL_B0|_RX|4 _PTL_B0|_RX|7 B0_RX  2.058e-12
L_PTL_B0|_RX|P1 _PTL_B0|_RX|2 0  4.795e-13
L_PTL_B0|_RX|P2 _PTL_B0|_RX|5 0  5.431e-13
L_PTL_B0|_RX|P3 _PTL_B0|_RX|8 0  5.339e-13
R_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|101  4.225701121488
R_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|104  3.429952209
R_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|107  2.7439617672
L_PTL_B0|_RX|RB1 _PTL_B0|_RX|101 0  2.38752113364072e-12
L_PTL_B0|_RX|RB2 _PTL_B0|_RX|104 0  1.937922998085e-12
L_PTL_B0|_RX|RB3 _PTL_B0|_RX|107 0  1.550338398468e-12
B_PTL_A1|_TX|1 _PTL_A1|_TX|1 _PTL_A1|_TX|2 JJMIT AREA=2.5
B_PTL_A1|_TX|2 _PTL_A1|_TX|4 _PTL_A1|_TX|5 JJMIT AREA=2.5
I_PTL_A1|_TX|B1 0 _PTL_A1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A1|_TX|B2 0 _PTL_A1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|3  1.684e-12
L_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|6  3.596e-12
L_PTL_A1|_TX|1 A1 _PTL_A1|_TX|1  2.063e-12
L_PTL_A1|_TX|2 _PTL_A1|_TX|1 _PTL_A1|_TX|4  4.123e-12
L_PTL_A1|_TX|3 _PTL_A1|_TX|4 _PTL_A1|_TX|7  2.193e-12
R_PTL_A1|_TX|D _PTL_A1|_TX|7 _PTL_A1|A_PTL  1.36
L_PTL_A1|_TX|P1 _PTL_A1|_TX|2 0  5.254e-13
L_PTL_A1|_TX|P2 _PTL_A1|_TX|5 0  5.141e-13
R_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|101  2.7439617672
R_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|104  2.7439617672
L_PTL_A1|_TX|RB1 _PTL_A1|_TX|101 0  1.550338398468e-12
L_PTL_A1|_TX|RB2 _PTL_A1|_TX|104 0  1.550338398468e-12
B_PTL_A1|_RX|1 _PTL_A1|_RX|1 _PTL_A1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A1|_RX|2 _PTL_A1|_RX|4 _PTL_A1|_RX|5 JJMIT AREA=2.0
B_PTL_A1|_RX|3 _PTL_A1|_RX|7 _PTL_A1|_RX|8 JJMIT AREA=2.5
I_PTL_A1|_RX|B1 0 _PTL_A1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|3  2.777e-12
I_PTL_A1|_RX|B2 0 _PTL_A1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|6  2.685e-12
I_PTL_A1|_RX|B3 0 _PTL_A1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|9  2.764e-12
L_PTL_A1|_RX|1 _PTL_A1|A_PTL _PTL_A1|_RX|1  1.346e-12
L_PTL_A1|_RX|2 _PTL_A1|_RX|1 _PTL_A1|_RX|4  6.348e-12
L_PTL_A1|_RX|3 _PTL_A1|_RX|4 _PTL_A1|_RX|7  5.197e-12
L_PTL_A1|_RX|4 _PTL_A1|_RX|7 A1_RX  2.058e-12
L_PTL_A1|_RX|P1 _PTL_A1|_RX|2 0  4.795e-13
L_PTL_A1|_RX|P2 _PTL_A1|_RX|5 0  5.431e-13
L_PTL_A1|_RX|P3 _PTL_A1|_RX|8 0  5.339e-13
R_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|101  4.225701121488
R_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|104  3.429952209
R_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|107  2.7439617672
L_PTL_A1|_RX|RB1 _PTL_A1|_RX|101 0  2.38752113364072e-12
L_PTL_A1|_RX|RB2 _PTL_A1|_RX|104 0  1.937922998085e-12
L_PTL_A1|_RX|RB3 _PTL_A1|_RX|107 0  1.550338398468e-12
B_PTL_B1|_TX|1 _PTL_B1|_TX|1 _PTL_B1|_TX|2 JJMIT AREA=2.5
B_PTL_B1|_TX|2 _PTL_B1|_TX|4 _PTL_B1|_TX|5 JJMIT AREA=2.5
I_PTL_B1|_TX|B1 0 _PTL_B1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B1|_TX|B2 0 _PTL_B1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|3  1.684e-12
L_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|6  3.596e-12
L_PTL_B1|_TX|1 B1 _PTL_B1|_TX|1  2.063e-12
L_PTL_B1|_TX|2 _PTL_B1|_TX|1 _PTL_B1|_TX|4  4.123e-12
L_PTL_B1|_TX|3 _PTL_B1|_TX|4 _PTL_B1|_TX|7  2.193e-12
R_PTL_B1|_TX|D _PTL_B1|_TX|7 _PTL_B1|A_PTL  1.36
L_PTL_B1|_TX|P1 _PTL_B1|_TX|2 0  5.254e-13
L_PTL_B1|_TX|P2 _PTL_B1|_TX|5 0  5.141e-13
R_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|101  2.7439617672
R_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|104  2.7439617672
L_PTL_B1|_TX|RB1 _PTL_B1|_TX|101 0  1.550338398468e-12
L_PTL_B1|_TX|RB2 _PTL_B1|_TX|104 0  1.550338398468e-12
B_PTL_B1|_RX|1 _PTL_B1|_RX|1 _PTL_B1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B1|_RX|2 _PTL_B1|_RX|4 _PTL_B1|_RX|5 JJMIT AREA=2.0
B_PTL_B1|_RX|3 _PTL_B1|_RX|7 _PTL_B1|_RX|8 JJMIT AREA=2.5
I_PTL_B1|_RX|B1 0 _PTL_B1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|3  2.777e-12
I_PTL_B1|_RX|B2 0 _PTL_B1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|6  2.685e-12
I_PTL_B1|_RX|B3 0 _PTL_B1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|9  2.764e-12
L_PTL_B1|_RX|1 _PTL_B1|A_PTL _PTL_B1|_RX|1  1.346e-12
L_PTL_B1|_RX|2 _PTL_B1|_RX|1 _PTL_B1|_RX|4  6.348e-12
L_PTL_B1|_RX|3 _PTL_B1|_RX|4 _PTL_B1|_RX|7  5.197e-12
L_PTL_B1|_RX|4 _PTL_B1|_RX|7 B1_RX  2.058e-12
L_PTL_B1|_RX|P1 _PTL_B1|_RX|2 0  4.795e-13
L_PTL_B1|_RX|P2 _PTL_B1|_RX|5 0  5.431e-13
L_PTL_B1|_RX|P3 _PTL_B1|_RX|8 0  5.339e-13
R_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|101  4.225701121488
R_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|104  3.429952209
R_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|107  2.7439617672
L_PTL_B1|_RX|RB1 _PTL_B1|_RX|101 0  2.38752113364072e-12
L_PTL_B1|_RX|RB2 _PTL_B1|_RX|104 0  1.937922998085e-12
L_PTL_B1|_RX|RB3 _PTL_B1|_RX|107 0  1.550338398468e-12
B_PTL_A2|_TX|1 _PTL_A2|_TX|1 _PTL_A2|_TX|2 JJMIT AREA=2.5
B_PTL_A2|_TX|2 _PTL_A2|_TX|4 _PTL_A2|_TX|5 JJMIT AREA=2.5
I_PTL_A2|_TX|B1 0 _PTL_A2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A2|_TX|B2 0 _PTL_A2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|3  1.684e-12
L_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|6  3.596e-12
L_PTL_A2|_TX|1 A2 _PTL_A2|_TX|1  2.063e-12
L_PTL_A2|_TX|2 _PTL_A2|_TX|1 _PTL_A2|_TX|4  4.123e-12
L_PTL_A2|_TX|3 _PTL_A2|_TX|4 _PTL_A2|_TX|7  2.193e-12
R_PTL_A2|_TX|D _PTL_A2|_TX|7 _PTL_A2|A_PTL  1.36
L_PTL_A2|_TX|P1 _PTL_A2|_TX|2 0  5.254e-13
L_PTL_A2|_TX|P2 _PTL_A2|_TX|5 0  5.141e-13
R_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|101  2.7439617672
R_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|104  2.7439617672
L_PTL_A2|_TX|RB1 _PTL_A2|_TX|101 0  1.550338398468e-12
L_PTL_A2|_TX|RB2 _PTL_A2|_TX|104 0  1.550338398468e-12
B_PTL_A2|_RX|1 _PTL_A2|_RX|1 _PTL_A2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A2|_RX|2 _PTL_A2|_RX|4 _PTL_A2|_RX|5 JJMIT AREA=2.0
B_PTL_A2|_RX|3 _PTL_A2|_RX|7 _PTL_A2|_RX|8 JJMIT AREA=2.5
I_PTL_A2|_RX|B1 0 _PTL_A2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|3  2.777e-12
I_PTL_A2|_RX|B2 0 _PTL_A2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|6  2.685e-12
I_PTL_A2|_RX|B3 0 _PTL_A2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|9  2.764e-12
L_PTL_A2|_RX|1 _PTL_A2|A_PTL _PTL_A2|_RX|1  1.346e-12
L_PTL_A2|_RX|2 _PTL_A2|_RX|1 _PTL_A2|_RX|4  6.348e-12
L_PTL_A2|_RX|3 _PTL_A2|_RX|4 _PTL_A2|_RX|7  5.197e-12
L_PTL_A2|_RX|4 _PTL_A2|_RX|7 A2_RX  2.058e-12
L_PTL_A2|_RX|P1 _PTL_A2|_RX|2 0  4.795e-13
L_PTL_A2|_RX|P2 _PTL_A2|_RX|5 0  5.431e-13
L_PTL_A2|_RX|P3 _PTL_A2|_RX|8 0  5.339e-13
R_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|101  4.225701121488
R_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|104  3.429952209
R_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|107  2.7439617672
L_PTL_A2|_RX|RB1 _PTL_A2|_RX|101 0  2.38752113364072e-12
L_PTL_A2|_RX|RB2 _PTL_A2|_RX|104 0  1.937922998085e-12
L_PTL_A2|_RX|RB3 _PTL_A2|_RX|107 0  1.550338398468e-12
B_PTL_B2|_TX|1 _PTL_B2|_TX|1 _PTL_B2|_TX|2 JJMIT AREA=2.5
B_PTL_B2|_TX|2 _PTL_B2|_TX|4 _PTL_B2|_TX|5 JJMIT AREA=2.5
I_PTL_B2|_TX|B1 0 _PTL_B2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B2|_TX|B2 0 _PTL_B2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|3  1.684e-12
L_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|6  3.596e-12
L_PTL_B2|_TX|1 B2 _PTL_B2|_TX|1  2.063e-12
L_PTL_B2|_TX|2 _PTL_B2|_TX|1 _PTL_B2|_TX|4  4.123e-12
L_PTL_B2|_TX|3 _PTL_B2|_TX|4 _PTL_B2|_TX|7  2.193e-12
R_PTL_B2|_TX|D _PTL_B2|_TX|7 _PTL_B2|A_PTL  1.36
L_PTL_B2|_TX|P1 _PTL_B2|_TX|2 0  5.254e-13
L_PTL_B2|_TX|P2 _PTL_B2|_TX|5 0  5.141e-13
R_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|101  2.7439617672
R_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|104  2.7439617672
L_PTL_B2|_TX|RB1 _PTL_B2|_TX|101 0  1.550338398468e-12
L_PTL_B2|_TX|RB2 _PTL_B2|_TX|104 0  1.550338398468e-12
B_PTL_B2|_RX|1 _PTL_B2|_RX|1 _PTL_B2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B2|_RX|2 _PTL_B2|_RX|4 _PTL_B2|_RX|5 JJMIT AREA=2.0
B_PTL_B2|_RX|3 _PTL_B2|_RX|7 _PTL_B2|_RX|8 JJMIT AREA=2.5
I_PTL_B2|_RX|B1 0 _PTL_B2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|3  2.777e-12
I_PTL_B2|_RX|B2 0 _PTL_B2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|6  2.685e-12
I_PTL_B2|_RX|B3 0 _PTL_B2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|9  2.764e-12
L_PTL_B2|_RX|1 _PTL_B2|A_PTL _PTL_B2|_RX|1  1.346e-12
L_PTL_B2|_RX|2 _PTL_B2|_RX|1 _PTL_B2|_RX|4  6.348e-12
L_PTL_B2|_RX|3 _PTL_B2|_RX|4 _PTL_B2|_RX|7  5.197e-12
L_PTL_B2|_RX|4 _PTL_B2|_RX|7 B2_RX  2.058e-12
L_PTL_B2|_RX|P1 _PTL_B2|_RX|2 0  4.795e-13
L_PTL_B2|_RX|P2 _PTL_B2|_RX|5 0  5.431e-13
L_PTL_B2|_RX|P3 _PTL_B2|_RX|8 0  5.339e-13
R_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|101  4.225701121488
R_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|104  3.429952209
R_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|107  2.7439617672
L_PTL_B2|_RX|RB1 _PTL_B2|_RX|101 0  2.38752113364072e-12
L_PTL_B2|_RX|RB2 _PTL_B2|_RX|104 0  1.937922998085e-12
L_PTL_B2|_RX|RB3 _PTL_B2|_RX|107 0  1.550338398468e-12
B_PTL_A3|_TX|1 _PTL_A3|_TX|1 _PTL_A3|_TX|2 JJMIT AREA=2.5
B_PTL_A3|_TX|2 _PTL_A3|_TX|4 _PTL_A3|_TX|5 JJMIT AREA=2.5
I_PTL_A3|_TX|B1 0 _PTL_A3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A3|_TX|B2 0 _PTL_A3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|3  1.684e-12
L_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|6  3.596e-12
L_PTL_A3|_TX|1 A3 _PTL_A3|_TX|1  2.063e-12
L_PTL_A3|_TX|2 _PTL_A3|_TX|1 _PTL_A3|_TX|4  4.123e-12
L_PTL_A3|_TX|3 _PTL_A3|_TX|4 _PTL_A3|_TX|7  2.193e-12
R_PTL_A3|_TX|D _PTL_A3|_TX|7 _PTL_A3|A_PTL  1.36
L_PTL_A3|_TX|P1 _PTL_A3|_TX|2 0  5.254e-13
L_PTL_A3|_TX|P2 _PTL_A3|_TX|5 0  5.141e-13
R_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|101  2.7439617672
R_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|104  2.7439617672
L_PTL_A3|_TX|RB1 _PTL_A3|_TX|101 0  1.550338398468e-12
L_PTL_A3|_TX|RB2 _PTL_A3|_TX|104 0  1.550338398468e-12
B_PTL_A3|_RX|1 _PTL_A3|_RX|1 _PTL_A3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A3|_RX|2 _PTL_A3|_RX|4 _PTL_A3|_RX|5 JJMIT AREA=2.0
B_PTL_A3|_RX|3 _PTL_A3|_RX|7 _PTL_A3|_RX|8 JJMIT AREA=2.5
I_PTL_A3|_RX|B1 0 _PTL_A3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|3  2.777e-12
I_PTL_A3|_RX|B2 0 _PTL_A3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|6  2.685e-12
I_PTL_A3|_RX|B3 0 _PTL_A3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|9  2.764e-12
L_PTL_A3|_RX|1 _PTL_A3|A_PTL _PTL_A3|_RX|1  1.346e-12
L_PTL_A3|_RX|2 _PTL_A3|_RX|1 _PTL_A3|_RX|4  6.348e-12
L_PTL_A3|_RX|3 _PTL_A3|_RX|4 _PTL_A3|_RX|7  5.197e-12
L_PTL_A3|_RX|4 _PTL_A3|_RX|7 A3_RX  2.058e-12
L_PTL_A3|_RX|P1 _PTL_A3|_RX|2 0  4.795e-13
L_PTL_A3|_RX|P2 _PTL_A3|_RX|5 0  5.431e-13
L_PTL_A3|_RX|P3 _PTL_A3|_RX|8 0  5.339e-13
R_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|101  4.225701121488
R_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|104  3.429952209
R_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|107  2.7439617672
L_PTL_A3|_RX|RB1 _PTL_A3|_RX|101 0  2.38752113364072e-12
L_PTL_A3|_RX|RB2 _PTL_A3|_RX|104 0  1.937922998085e-12
L_PTL_A3|_RX|RB3 _PTL_A3|_RX|107 0  1.550338398468e-12
B_PTL_B3|_TX|1 _PTL_B3|_TX|1 _PTL_B3|_TX|2 JJMIT AREA=2.5
B_PTL_B3|_TX|2 _PTL_B3|_TX|4 _PTL_B3|_TX|5 JJMIT AREA=2.5
I_PTL_B3|_TX|B1 0 _PTL_B3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B3|_TX|B2 0 _PTL_B3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|3  1.684e-12
L_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|6  3.596e-12
L_PTL_B3|_TX|1 B3 _PTL_B3|_TX|1  2.063e-12
L_PTL_B3|_TX|2 _PTL_B3|_TX|1 _PTL_B3|_TX|4  4.123e-12
L_PTL_B3|_TX|3 _PTL_B3|_TX|4 _PTL_B3|_TX|7  2.193e-12
R_PTL_B3|_TX|D _PTL_B3|_TX|7 _PTL_B3|A_PTL  1.36
L_PTL_B3|_TX|P1 _PTL_B3|_TX|2 0  5.254e-13
L_PTL_B3|_TX|P2 _PTL_B3|_TX|5 0  5.141e-13
R_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|101  2.7439617672
R_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|104  2.7439617672
L_PTL_B3|_TX|RB1 _PTL_B3|_TX|101 0  1.550338398468e-12
L_PTL_B3|_TX|RB2 _PTL_B3|_TX|104 0  1.550338398468e-12
B_PTL_B3|_RX|1 _PTL_B3|_RX|1 _PTL_B3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B3|_RX|2 _PTL_B3|_RX|4 _PTL_B3|_RX|5 JJMIT AREA=2.0
B_PTL_B3|_RX|3 _PTL_B3|_RX|7 _PTL_B3|_RX|8 JJMIT AREA=2.5
I_PTL_B3|_RX|B1 0 _PTL_B3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|3  2.777e-12
I_PTL_B3|_RX|B2 0 _PTL_B3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|6  2.685e-12
I_PTL_B3|_RX|B3 0 _PTL_B3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|9  2.764e-12
L_PTL_B3|_RX|1 _PTL_B3|A_PTL _PTL_B3|_RX|1  1.346e-12
L_PTL_B3|_RX|2 _PTL_B3|_RX|1 _PTL_B3|_RX|4  6.348e-12
L_PTL_B3|_RX|3 _PTL_B3|_RX|4 _PTL_B3|_RX|7  5.197e-12
L_PTL_B3|_RX|4 _PTL_B3|_RX|7 B3_RX  2.058e-12
L_PTL_B3|_RX|P1 _PTL_B3|_RX|2 0  4.795e-13
L_PTL_B3|_RX|P2 _PTL_B3|_RX|5 0  5.431e-13
L_PTL_B3|_RX|P3 _PTL_B3|_RX|8 0  5.339e-13
R_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|101  4.225701121488
R_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|104  3.429952209
R_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|107  2.7439617672
L_PTL_B3|_RX|RB1 _PTL_B3|_RX|101 0  2.38752113364072e-12
L_PTL_B3|_RX|RB2 _PTL_B3|_RX|104 0  1.937922998085e-12
L_PTL_B3|_RX|RB3 _PTL_B3|_RX|107 0  1.550338398468e-12
LI0|_SPL_A|1 A0_RX I0|_SPL_A|D1  2e-12
LI0|_SPL_A|2 I0|_SPL_A|D1 I0|_SPL_A|D2  4.135667696e-12
LI0|_SPL_A|3 I0|_SPL_A|D2 I0|_SPL_A|JCT  9.84682784761905e-13
LI0|_SPL_A|4 I0|_SPL_A|JCT I0|_SPL_A|QA1  9.84682784761905e-13
LI0|_SPL_A|5 I0|_SPL_A|QA1 I0|A1  2e-12
LI0|_SPL_A|6 I0|_SPL_A|JCT I0|_SPL_A|QB1  9.84682784761905e-13
LI0|_SPL_A|7 I0|_SPL_A|QB1 I0|A2  2e-12
LI0|_SPL_B|1 B0_RX I0|_SPL_B|D1  2e-12
LI0|_SPL_B|2 I0|_SPL_B|D1 I0|_SPL_B|D2  4.135667696e-12
LI0|_SPL_B|3 I0|_SPL_B|D2 I0|_SPL_B|JCT  9.84682784761905e-13
LI0|_SPL_B|4 I0|_SPL_B|JCT I0|_SPL_B|QA1  9.84682784761905e-13
LI0|_SPL_B|5 I0|_SPL_B|QA1 I0|B1  2e-12
LI0|_SPL_B|6 I0|_SPL_B|JCT I0|_SPL_B|QB1  9.84682784761905e-13
LI0|_SPL_B|7 I0|_SPL_B|QB1 I0|B2  2e-12
LI0|_DFF_A|1 I0|A1 I0|_DFF_A|A1  2.067833848e-12
LI0|_DFF_A|2 I0|_DFF_A|A1 I0|_DFF_A|A2  4.135667696e-12
LI0|_DFF_A|3 I0|_DFF_A|A3 I0|_DFF_A|A4  8.271335392e-12
LI0|_DFF_A|T T00 I0|_DFF_A|T1  2.067833848e-12
LI0|_DFF_A|4 I0|_DFF_A|T1 I0|_DFF_A|T2  4.135667696e-12
LI0|_DFF_A|5 I0|_DFF_A|A4 I0|_DFF_A|Q1  4.135667696e-12
LI0|_DFF_A|6 I0|_DFF_A|Q1 I0|A1_SYNC  2.067833848e-12
LI0|_DFF_B|1 I0|B1 I0|_DFF_B|A1  2.067833848e-12
LI0|_DFF_B|2 I0|_DFF_B|A1 I0|_DFF_B|A2  4.135667696e-12
LI0|_DFF_B|3 I0|_DFF_B|A3 I0|_DFF_B|A4  8.271335392e-12
LI0|_DFF_B|T T00 I0|_DFF_B|T1  2.067833848e-12
LI0|_DFF_B|4 I0|_DFF_B|T1 I0|_DFF_B|T2  4.135667696e-12
LI0|_DFF_B|5 I0|_DFF_B|A4 I0|_DFF_B|Q1  4.135667696e-12
LI0|_DFF_B|6 I0|_DFF_B|Q1 I0|B1_SYNC  2.067833848e-12
LI0|_XOR|A1 I0|A2 I0|_XOR|A1  2.067833848e-12
LI0|_XOR|A2 I0|_XOR|A1 I0|_XOR|A2  4.135667696e-12
LI0|_XOR|A3 I0|_XOR|A3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|B1 I0|B2 I0|_XOR|B1  2.067833848e-12
LI0|_XOR|B2 I0|_XOR|B1 I0|_XOR|B2  4.135667696e-12
LI0|_XOR|B3 I0|_XOR|B3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|T1 T00 I0|_XOR|T1  2.067833848e-12
LI0|_XOR|T2 I0|_XOR|T1 I0|_XOR|T2  4.135667696e-12
LI0|_XOR|Q2 I0|_XOR|ABTQ I0|_XOR|Q1  4.135667696e-12
LI0|_XOR|Q1 I0|_XOR|Q1 IP0_0  2.067833848e-12
LI0|_AND|A1 I0|A1_SYNC I0|_AND|A1  2.067833848e-12
LI0|_AND|A2 I0|_AND|A1 I0|_AND|A2  4.135667696e-12
LI0|_AND|A3 I0|_AND|A3 I0|_AND|Q3  1.2e-12
LI0|_AND|B1 I0|B1_SYNC I0|_AND|B1  2.067833848e-12
LI0|_AND|B2 I0|_AND|B1 I0|_AND|B2  4.135667696e-12
LI0|_AND|B3 I0|_AND|B3 I0|_AND|Q3  1.2e-12
LI0|_AND|Q3 I0|_AND|Q3 I0|_AND|Q2  4.135667696e-12
LI0|_AND|Q2 I0|_AND|Q2 I0|_AND|Q1  4.135667696e-12
LI0|_AND|Q1 I0|_AND|Q1 IG0_0  2.067833848e-12
LI1|_SPL_A|1 A1_RX I1|_SPL_A|D1  2e-12
LI1|_SPL_A|2 I1|_SPL_A|D1 I1|_SPL_A|D2  4.135667696e-12
LI1|_SPL_A|3 I1|_SPL_A|D2 I1|_SPL_A|JCT  9.84682784761905e-13
LI1|_SPL_A|4 I1|_SPL_A|JCT I1|_SPL_A|QA1  9.84682784761905e-13
LI1|_SPL_A|5 I1|_SPL_A|QA1 I1|A1  2e-12
LI1|_SPL_A|6 I1|_SPL_A|JCT I1|_SPL_A|QB1  9.84682784761905e-13
LI1|_SPL_A|7 I1|_SPL_A|QB1 I1|A2  2e-12
LI1|_SPL_B|1 B1_RX I1|_SPL_B|D1  2e-12
LI1|_SPL_B|2 I1|_SPL_B|D1 I1|_SPL_B|D2  4.135667696e-12
LI1|_SPL_B|3 I1|_SPL_B|D2 I1|_SPL_B|JCT  9.84682784761905e-13
LI1|_SPL_B|4 I1|_SPL_B|JCT I1|_SPL_B|QA1  9.84682784761905e-13
LI1|_SPL_B|5 I1|_SPL_B|QA1 I1|B1  2e-12
LI1|_SPL_B|6 I1|_SPL_B|JCT I1|_SPL_B|QB1  9.84682784761905e-13
LI1|_SPL_B|7 I1|_SPL_B|QB1 I1|B2  2e-12
LI1|_DFF_A|1 I1|A1 I1|_DFF_A|A1  2.067833848e-12
LI1|_DFF_A|2 I1|_DFF_A|A1 I1|_DFF_A|A2  4.135667696e-12
LI1|_DFF_A|3 I1|_DFF_A|A3 I1|_DFF_A|A4  8.271335392e-12
LI1|_DFF_A|T T01 I1|_DFF_A|T1  2.067833848e-12
LI1|_DFF_A|4 I1|_DFF_A|T1 I1|_DFF_A|T2  4.135667696e-12
LI1|_DFF_A|5 I1|_DFF_A|A4 I1|_DFF_A|Q1  4.135667696e-12
LI1|_DFF_A|6 I1|_DFF_A|Q1 I1|A1_SYNC  2.067833848e-12
LI1|_DFF_B|1 I1|B1 I1|_DFF_B|A1  2.067833848e-12
LI1|_DFF_B|2 I1|_DFF_B|A1 I1|_DFF_B|A2  4.135667696e-12
LI1|_DFF_B|3 I1|_DFF_B|A3 I1|_DFF_B|A4  8.271335392e-12
LI1|_DFF_B|T T01 I1|_DFF_B|T1  2.067833848e-12
LI1|_DFF_B|4 I1|_DFF_B|T1 I1|_DFF_B|T2  4.135667696e-12
LI1|_DFF_B|5 I1|_DFF_B|A4 I1|_DFF_B|Q1  4.135667696e-12
LI1|_DFF_B|6 I1|_DFF_B|Q1 I1|B1_SYNC  2.067833848e-12
LI1|_XOR|A1 I1|A2 I1|_XOR|A1  2.067833848e-12
LI1|_XOR|A2 I1|_XOR|A1 I1|_XOR|A2  4.135667696e-12
LI1|_XOR|A3 I1|_XOR|A3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|B1 I1|B2 I1|_XOR|B1  2.067833848e-12
LI1|_XOR|B2 I1|_XOR|B1 I1|_XOR|B2  4.135667696e-12
LI1|_XOR|B3 I1|_XOR|B3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|T1 T01 I1|_XOR|T1  2.067833848e-12
LI1|_XOR|T2 I1|_XOR|T1 I1|_XOR|T2  4.135667696e-12
LI1|_XOR|Q2 I1|_XOR|ABTQ I1|_XOR|Q1  4.135667696e-12
LI1|_XOR|Q1 I1|_XOR|Q1 IP1_0  2.067833848e-12
LI1|_AND|A1 I1|A1_SYNC I1|_AND|A1  2.067833848e-12
LI1|_AND|A2 I1|_AND|A1 I1|_AND|A2  4.135667696e-12
LI1|_AND|A3 I1|_AND|A3 I1|_AND|Q3  1.2e-12
LI1|_AND|B1 I1|B1_SYNC I1|_AND|B1  2.067833848e-12
LI1|_AND|B2 I1|_AND|B1 I1|_AND|B2  4.135667696e-12
LI1|_AND|B3 I1|_AND|B3 I1|_AND|Q3  1.2e-12
LI1|_AND|Q3 I1|_AND|Q3 I1|_AND|Q2  4.135667696e-12
LI1|_AND|Q2 I1|_AND|Q2 I1|_AND|Q1  4.135667696e-12
LI1|_AND|Q1 I1|_AND|Q1 IG1_0  2.067833848e-12
LI2|_SPL_A|1 A2_RX I2|_SPL_A|D1  2e-12
LI2|_SPL_A|2 I2|_SPL_A|D1 I2|_SPL_A|D2  4.135667696e-12
LI2|_SPL_A|3 I2|_SPL_A|D2 I2|_SPL_A|JCT  9.84682784761905e-13
LI2|_SPL_A|4 I2|_SPL_A|JCT I2|_SPL_A|QA1  9.84682784761905e-13
LI2|_SPL_A|5 I2|_SPL_A|QA1 I2|A1  2e-12
LI2|_SPL_A|6 I2|_SPL_A|JCT I2|_SPL_A|QB1  9.84682784761905e-13
LI2|_SPL_A|7 I2|_SPL_A|QB1 I2|A2  2e-12
LI2|_SPL_B|1 B2_RX I2|_SPL_B|D1  2e-12
LI2|_SPL_B|2 I2|_SPL_B|D1 I2|_SPL_B|D2  4.135667696e-12
LI2|_SPL_B|3 I2|_SPL_B|D2 I2|_SPL_B|JCT  9.84682784761905e-13
LI2|_SPL_B|4 I2|_SPL_B|JCT I2|_SPL_B|QA1  9.84682784761905e-13
LI2|_SPL_B|5 I2|_SPL_B|QA1 I2|B1  2e-12
LI2|_SPL_B|6 I2|_SPL_B|JCT I2|_SPL_B|QB1  9.84682784761905e-13
LI2|_SPL_B|7 I2|_SPL_B|QB1 I2|B2  2e-12
LI2|_DFF_A|1 I2|A1 I2|_DFF_A|A1  2.067833848e-12
LI2|_DFF_A|2 I2|_DFF_A|A1 I2|_DFF_A|A2  4.135667696e-12
LI2|_DFF_A|3 I2|_DFF_A|A3 I2|_DFF_A|A4  8.271335392e-12
LI2|_DFF_A|T T02 I2|_DFF_A|T1  2.067833848e-12
LI2|_DFF_A|4 I2|_DFF_A|T1 I2|_DFF_A|T2  4.135667696e-12
LI2|_DFF_A|5 I2|_DFF_A|A4 I2|_DFF_A|Q1  4.135667696e-12
LI2|_DFF_A|6 I2|_DFF_A|Q1 I2|A1_SYNC  2.067833848e-12
LI2|_DFF_B|1 I2|B1 I2|_DFF_B|A1  2.067833848e-12
LI2|_DFF_B|2 I2|_DFF_B|A1 I2|_DFF_B|A2  4.135667696e-12
LI2|_DFF_B|3 I2|_DFF_B|A3 I2|_DFF_B|A4  8.271335392e-12
LI2|_DFF_B|T T02 I2|_DFF_B|T1  2.067833848e-12
LI2|_DFF_B|4 I2|_DFF_B|T1 I2|_DFF_B|T2  4.135667696e-12
LI2|_DFF_B|5 I2|_DFF_B|A4 I2|_DFF_B|Q1  4.135667696e-12
LI2|_DFF_B|6 I2|_DFF_B|Q1 I2|B1_SYNC  2.067833848e-12
LI2|_XOR|A1 I2|A2 I2|_XOR|A1  2.067833848e-12
LI2|_XOR|A2 I2|_XOR|A1 I2|_XOR|A2  4.135667696e-12
LI2|_XOR|A3 I2|_XOR|A3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|B1 I2|B2 I2|_XOR|B1  2.067833848e-12
LI2|_XOR|B2 I2|_XOR|B1 I2|_XOR|B2  4.135667696e-12
LI2|_XOR|B3 I2|_XOR|B3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|T1 T02 I2|_XOR|T1  2.067833848e-12
LI2|_XOR|T2 I2|_XOR|T1 I2|_XOR|T2  4.135667696e-12
LI2|_XOR|Q2 I2|_XOR|ABTQ I2|_XOR|Q1  4.135667696e-12
LI2|_XOR|Q1 I2|_XOR|Q1 IP2_0  2.067833848e-12
LI2|_AND|A1 I2|A1_SYNC I2|_AND|A1  2.067833848e-12
LI2|_AND|A2 I2|_AND|A1 I2|_AND|A2  4.135667696e-12
LI2|_AND|A3 I2|_AND|A3 I2|_AND|Q3  1.2e-12
LI2|_AND|B1 I2|B1_SYNC I2|_AND|B1  2.067833848e-12
LI2|_AND|B2 I2|_AND|B1 I2|_AND|B2  4.135667696e-12
LI2|_AND|B3 I2|_AND|B3 I2|_AND|Q3  1.2e-12
LI2|_AND|Q3 I2|_AND|Q3 I2|_AND|Q2  4.135667696e-12
LI2|_AND|Q2 I2|_AND|Q2 I2|_AND|Q1  4.135667696e-12
LI2|_AND|Q1 I2|_AND|Q1 IG2_0  2.067833848e-12
LI3|_SPL_A|1 A3_RX I3|_SPL_A|D1  2e-12
LI3|_SPL_A|2 I3|_SPL_A|D1 I3|_SPL_A|D2  4.135667696e-12
LI3|_SPL_A|3 I3|_SPL_A|D2 I3|_SPL_A|JCT  9.84682784761905e-13
LI3|_SPL_A|4 I3|_SPL_A|JCT I3|_SPL_A|QA1  9.84682784761905e-13
LI3|_SPL_A|5 I3|_SPL_A|QA1 I3|A1  2e-12
LI3|_SPL_A|6 I3|_SPL_A|JCT I3|_SPL_A|QB1  9.84682784761905e-13
LI3|_SPL_A|7 I3|_SPL_A|QB1 I3|A2  2e-12
LI3|_SPL_B|1 B3_RX I3|_SPL_B|D1  2e-12
LI3|_SPL_B|2 I3|_SPL_B|D1 I3|_SPL_B|D2  4.135667696e-12
LI3|_SPL_B|3 I3|_SPL_B|D2 I3|_SPL_B|JCT  9.84682784761905e-13
LI3|_SPL_B|4 I3|_SPL_B|JCT I3|_SPL_B|QA1  9.84682784761905e-13
LI3|_SPL_B|5 I3|_SPL_B|QA1 I3|B1  2e-12
LI3|_SPL_B|6 I3|_SPL_B|JCT I3|_SPL_B|QB1  9.84682784761905e-13
LI3|_SPL_B|7 I3|_SPL_B|QB1 I3|B2  2e-12
LI3|_DFF_A|1 I3|A1 I3|_DFF_A|A1  2.067833848e-12
LI3|_DFF_A|2 I3|_DFF_A|A1 I3|_DFF_A|A2  4.135667696e-12
LI3|_DFF_A|3 I3|_DFF_A|A3 I3|_DFF_A|A4  8.271335392e-12
LI3|_DFF_A|T T03 I3|_DFF_A|T1  2.067833848e-12
LI3|_DFF_A|4 I3|_DFF_A|T1 I3|_DFF_A|T2  4.135667696e-12
LI3|_DFF_A|5 I3|_DFF_A|A4 I3|_DFF_A|Q1  4.135667696e-12
LI3|_DFF_A|6 I3|_DFF_A|Q1 I3|A1_SYNC  2.067833848e-12
LI3|_DFF_B|1 I3|B1 I3|_DFF_B|A1  2.067833848e-12
LI3|_DFF_B|2 I3|_DFF_B|A1 I3|_DFF_B|A2  4.135667696e-12
LI3|_DFF_B|3 I3|_DFF_B|A3 I3|_DFF_B|A4  8.271335392e-12
LI3|_DFF_B|T T03 I3|_DFF_B|T1  2.067833848e-12
LI3|_DFF_B|4 I3|_DFF_B|T1 I3|_DFF_B|T2  4.135667696e-12
LI3|_DFF_B|5 I3|_DFF_B|A4 I3|_DFF_B|Q1  4.135667696e-12
LI3|_DFF_B|6 I3|_DFF_B|Q1 I3|B1_SYNC  2.067833848e-12
LI3|_XOR|A1 I3|A2 I3|_XOR|A1  2.067833848e-12
LI3|_XOR|A2 I3|_XOR|A1 I3|_XOR|A2  4.135667696e-12
LI3|_XOR|A3 I3|_XOR|A3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|B1 I3|B2 I3|_XOR|B1  2.067833848e-12
LI3|_XOR|B2 I3|_XOR|B1 I3|_XOR|B2  4.135667696e-12
LI3|_XOR|B3 I3|_XOR|B3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|T1 T03 I3|_XOR|T1  2.067833848e-12
LI3|_XOR|T2 I3|_XOR|T1 I3|_XOR|T2  4.135667696e-12
LI3|_XOR|Q2 I3|_XOR|ABTQ I3|_XOR|Q1  4.135667696e-12
LI3|_XOR|Q1 I3|_XOR|Q1 IP3_0  2.067833848e-12
LI3|_AND|A1 I3|A1_SYNC I3|_AND|A1  2.067833848e-12
LI3|_AND|A2 I3|_AND|A1 I3|_AND|A2  4.135667696e-12
LI3|_AND|A3 I3|_AND|A3 I3|_AND|Q3  1.2e-12
LI3|_AND|B1 I3|B1_SYNC I3|_AND|B1  2.067833848e-12
LI3|_AND|B2 I3|_AND|B1 I3|_AND|B2  4.135667696e-12
LI3|_AND|B3 I3|_AND|B3 I3|_AND|Q3  1.2e-12
LI3|_AND|Q3 I3|_AND|Q3 I3|_AND|Q2  4.135667696e-12
LI3|_AND|Q2 I3|_AND|Q2 I3|_AND|Q1  4.135667696e-12
LI3|_AND|Q1 I3|_AND|Q1 IG3_0  2.067833848e-12
B_PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP0_0|_TX|B1 0 _PTL_IP0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP0_0|_TX|B2 0 _PTL_IP0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|3  1.684e-12
L_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|6  3.596e-12
L_PTL_IP0_0|_TX|1 IP0_0 _PTL_IP0_0|_TX|1  2.063e-12
L_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|4  4.123e-12
L_PTL_IP0_0|_TX|3 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|7  2.193e-12
R_PTL_IP0_0|_TX|D _PTL_IP0_0|_TX|7 _PTL_IP0_0|A_PTL  1.36
L_PTL_IP0_0|_TX|P1 _PTL_IP0_0|_TX|2 0  5.254e-13
L_PTL_IP0_0|_TX|P2 _PTL_IP0_0|_TX|5 0  5.141e-13
R_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|101  2.7439617672
R_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|104  2.7439617672
L_PTL_IP0_0|_TX|RB1 _PTL_IP0_0|_TX|101 0  1.550338398468e-12
L_PTL_IP0_0|_TX|RB2 _PTL_IP0_0|_TX|104 0  1.550338398468e-12
B_PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP0_0|_RX|B1 0 _PTL_IP0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|3  2.777e-12
I_PTL_IP0_0|_RX|B2 0 _PTL_IP0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|6  2.685e-12
I_PTL_IP0_0|_RX|B3 0 _PTL_IP0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|9  2.764e-12
L_PTL_IP0_0|_RX|1 _PTL_IP0_0|A_PTL _PTL_IP0_0|_RX|1  1.346e-12
L_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|4  6.348e-12
L_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7  5.197e-12
L_PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7 IP0_0_RX  2.058e-12
L_PTL_IP0_0|_RX|P1 _PTL_IP0_0|_RX|2 0  4.795e-13
L_PTL_IP0_0|_RX|P2 _PTL_IP0_0|_RX|5 0  5.431e-13
L_PTL_IP0_0|_RX|P3 _PTL_IP0_0|_RX|8 0  5.339e-13
R_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|101  4.225701121488
R_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|104  3.429952209
R_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|107  2.7439617672
L_PTL_IP0_0|_RX|RB1 _PTL_IP0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP0_0|_RX|RB2 _PTL_IP0_0|_RX|104 0  1.937922998085e-12
L_PTL_IP0_0|_RX|RB3 _PTL_IP0_0|_RX|107 0  1.550338398468e-12
B_PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG0_0|_TX|B1 0 _PTL_IG0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG0_0|_TX|B2 0 _PTL_IG0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|3  1.684e-12
L_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|6  3.596e-12
L_PTL_IG0_0|_TX|1 IG0_0 _PTL_IG0_0|_TX|1  2.063e-12
L_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|4  4.123e-12
L_PTL_IG0_0|_TX|3 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|7  2.193e-12
R_PTL_IG0_0|_TX|D _PTL_IG0_0|_TX|7 _PTL_IG0_0|A_PTL  1.36
L_PTL_IG0_0|_TX|P1 _PTL_IG0_0|_TX|2 0  5.254e-13
L_PTL_IG0_0|_TX|P2 _PTL_IG0_0|_TX|5 0  5.141e-13
R_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|101  2.7439617672
R_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|104  2.7439617672
L_PTL_IG0_0|_TX|RB1 _PTL_IG0_0|_TX|101 0  1.550338398468e-12
L_PTL_IG0_0|_TX|RB2 _PTL_IG0_0|_TX|104 0  1.550338398468e-12
B_PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG0_0|_RX|B1 0 _PTL_IG0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|3  2.777e-12
I_PTL_IG0_0|_RX|B2 0 _PTL_IG0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|6  2.685e-12
I_PTL_IG0_0|_RX|B3 0 _PTL_IG0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|9  2.764e-12
L_PTL_IG0_0|_RX|1 _PTL_IG0_0|A_PTL _PTL_IG0_0|_RX|1  1.346e-12
L_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|4  6.348e-12
L_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7  5.197e-12
L_PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7 IG0_0_RX  2.058e-12
L_PTL_IG0_0|_RX|P1 _PTL_IG0_0|_RX|2 0  4.795e-13
L_PTL_IG0_0|_RX|P2 _PTL_IG0_0|_RX|5 0  5.431e-13
L_PTL_IG0_0|_RX|P3 _PTL_IG0_0|_RX|8 0  5.339e-13
R_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|101  4.225701121488
R_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|104  3.429952209
R_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|107  2.7439617672
L_PTL_IG0_0|_RX|RB1 _PTL_IG0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG0_0|_RX|RB2 _PTL_IG0_0|_RX|104 0  1.937922998085e-12
L_PTL_IG0_0|_RX|RB3 _PTL_IG0_0|_RX|107 0  1.550338398468e-12
B_PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_0|_TX|B1 0 _PTL_IP1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_0|_TX|B2 0 _PTL_IP1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|3  1.684e-12
L_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|6  3.596e-12
L_PTL_IP1_0|_TX|1 IP1_0 _PTL_IP1_0|_TX|1  2.063e-12
L_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|4  4.123e-12
L_PTL_IP1_0|_TX|3 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|7  2.193e-12
R_PTL_IP1_0|_TX|D _PTL_IP1_0|_TX|7 _PTL_IP1_0|A_PTL  1.36
L_PTL_IP1_0|_TX|P1 _PTL_IP1_0|_TX|2 0  5.254e-13
L_PTL_IP1_0|_TX|P2 _PTL_IP1_0|_TX|5 0  5.141e-13
R_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|101  2.7439617672
R_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|104  2.7439617672
L_PTL_IP1_0|_TX|RB1 _PTL_IP1_0|_TX|101 0  1.550338398468e-12
L_PTL_IP1_0|_TX|RB2 _PTL_IP1_0|_TX|104 0  1.550338398468e-12
B_PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_0|_RX|B1 0 _PTL_IP1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|3  2.777e-12
I_PTL_IP1_0|_RX|B2 0 _PTL_IP1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|6  2.685e-12
I_PTL_IP1_0|_RX|B3 0 _PTL_IP1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|9  2.764e-12
L_PTL_IP1_0|_RX|1 _PTL_IP1_0|A_PTL _PTL_IP1_0|_RX|1  1.346e-12
L_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|4  6.348e-12
L_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7  5.197e-12
L_PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7 IP1_0_RX  2.058e-12
L_PTL_IP1_0|_RX|P1 _PTL_IP1_0|_RX|2 0  4.795e-13
L_PTL_IP1_0|_RX|P2 _PTL_IP1_0|_RX|5 0  5.431e-13
L_PTL_IP1_0|_RX|P3 _PTL_IP1_0|_RX|8 0  5.339e-13
R_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|101  4.225701121488
R_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|104  3.429952209
R_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|107  2.7439617672
L_PTL_IP1_0|_RX|RB1 _PTL_IP1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_0|_RX|RB2 _PTL_IP1_0|_RX|104 0  1.937922998085e-12
L_PTL_IP1_0|_RX|RB3 _PTL_IP1_0|_RX|107 0  1.550338398468e-12
B_PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG1_0|_TX|B1 0 _PTL_IG1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG1_0|_TX|B2 0 _PTL_IG1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|3  1.684e-12
L_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|6  3.596e-12
L_PTL_IG1_0|_TX|1 IG1_0 _PTL_IG1_0|_TX|1  2.063e-12
L_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|4  4.123e-12
L_PTL_IG1_0|_TX|3 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|7  2.193e-12
R_PTL_IG1_0|_TX|D _PTL_IG1_0|_TX|7 _PTL_IG1_0|A_PTL  1.36
L_PTL_IG1_0|_TX|P1 _PTL_IG1_0|_TX|2 0  5.254e-13
L_PTL_IG1_0|_TX|P2 _PTL_IG1_0|_TX|5 0  5.141e-13
R_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|101  2.7439617672
R_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|104  2.7439617672
L_PTL_IG1_0|_TX|RB1 _PTL_IG1_0|_TX|101 0  1.550338398468e-12
L_PTL_IG1_0|_TX|RB2 _PTL_IG1_0|_TX|104 0  1.550338398468e-12
B_PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG1_0|_RX|B1 0 _PTL_IG1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|3  2.777e-12
I_PTL_IG1_0|_RX|B2 0 _PTL_IG1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|6  2.685e-12
I_PTL_IG1_0|_RX|B3 0 _PTL_IG1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|9  2.764e-12
L_PTL_IG1_0|_RX|1 _PTL_IG1_0|A_PTL _PTL_IG1_0|_RX|1  1.346e-12
L_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|4  6.348e-12
L_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7  5.197e-12
L_PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7 IG1_0_RX  2.058e-12
L_PTL_IG1_0|_RX|P1 _PTL_IG1_0|_RX|2 0  4.795e-13
L_PTL_IG1_0|_RX|P2 _PTL_IG1_0|_RX|5 0  5.431e-13
L_PTL_IG1_0|_RX|P3 _PTL_IG1_0|_RX|8 0  5.339e-13
R_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|101  4.225701121488
R_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|104  3.429952209
R_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|107  2.7439617672
L_PTL_IG1_0|_RX|RB1 _PTL_IG1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG1_0|_RX|RB2 _PTL_IG1_0|_RX|104 0  1.937922998085e-12
L_PTL_IG1_0|_RX|RB3 _PTL_IG1_0|_RX|107 0  1.550338398468e-12
B_PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_0|_TX|B1 0 _PTL_IP2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_0|_TX|B2 0 _PTL_IP2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|3  1.684e-12
L_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|6  3.596e-12
L_PTL_IP2_0|_TX|1 IP2_0 _PTL_IP2_0|_TX|1  2.063e-12
L_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|4  4.123e-12
L_PTL_IP2_0|_TX|3 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|7  2.193e-12
R_PTL_IP2_0|_TX|D _PTL_IP2_0|_TX|7 _PTL_IP2_0|A_PTL  1.36
L_PTL_IP2_0|_TX|P1 _PTL_IP2_0|_TX|2 0  5.254e-13
L_PTL_IP2_0|_TX|P2 _PTL_IP2_0|_TX|5 0  5.141e-13
R_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|101  2.7439617672
R_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|104  2.7439617672
L_PTL_IP2_0|_TX|RB1 _PTL_IP2_0|_TX|101 0  1.550338398468e-12
L_PTL_IP2_0|_TX|RB2 _PTL_IP2_0|_TX|104 0  1.550338398468e-12
B_PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_0|_RX|B1 0 _PTL_IP2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|3  2.777e-12
I_PTL_IP2_0|_RX|B2 0 _PTL_IP2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|6  2.685e-12
I_PTL_IP2_0|_RX|B3 0 _PTL_IP2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|9  2.764e-12
L_PTL_IP2_0|_RX|1 _PTL_IP2_0|A_PTL _PTL_IP2_0|_RX|1  1.346e-12
L_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|4  6.348e-12
L_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7  5.197e-12
L_PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7 IP2_0_RX  2.058e-12
L_PTL_IP2_0|_RX|P1 _PTL_IP2_0|_RX|2 0  4.795e-13
L_PTL_IP2_0|_RX|P2 _PTL_IP2_0|_RX|5 0  5.431e-13
L_PTL_IP2_0|_RX|P3 _PTL_IP2_0|_RX|8 0  5.339e-13
R_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|101  4.225701121488
R_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|104  3.429952209
R_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|107  2.7439617672
L_PTL_IP2_0|_RX|RB1 _PTL_IP2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_0|_RX|RB2 _PTL_IP2_0|_RX|104 0  1.937922998085e-12
L_PTL_IP2_0|_RX|RB3 _PTL_IP2_0|_RX|107 0  1.550338398468e-12
B_PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG2_0|_TX|B1 0 _PTL_IG2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG2_0|_TX|B2 0 _PTL_IG2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|3  1.684e-12
L_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|6  3.596e-12
L_PTL_IG2_0|_TX|1 IG2_0 _PTL_IG2_0|_TX|1  2.063e-12
L_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|4  4.123e-12
L_PTL_IG2_0|_TX|3 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|7  2.193e-12
R_PTL_IG2_0|_TX|D _PTL_IG2_0|_TX|7 _PTL_IG2_0|A_PTL  1.36
L_PTL_IG2_0|_TX|P1 _PTL_IG2_0|_TX|2 0  5.254e-13
L_PTL_IG2_0|_TX|P2 _PTL_IG2_0|_TX|5 0  5.141e-13
R_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|101  2.7439617672
R_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|104  2.7439617672
L_PTL_IG2_0|_TX|RB1 _PTL_IG2_0|_TX|101 0  1.550338398468e-12
L_PTL_IG2_0|_TX|RB2 _PTL_IG2_0|_TX|104 0  1.550338398468e-12
B_PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG2_0|_RX|B1 0 _PTL_IG2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|3  2.777e-12
I_PTL_IG2_0|_RX|B2 0 _PTL_IG2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|6  2.685e-12
I_PTL_IG2_0|_RX|B3 0 _PTL_IG2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|9  2.764e-12
L_PTL_IG2_0|_RX|1 _PTL_IG2_0|A_PTL _PTL_IG2_0|_RX|1  1.346e-12
L_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|4  6.348e-12
L_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7  5.197e-12
L_PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7 IG2_0_RX  2.058e-12
L_PTL_IG2_0|_RX|P1 _PTL_IG2_0|_RX|2 0  4.795e-13
L_PTL_IG2_0|_RX|P2 _PTL_IG2_0|_RX|5 0  5.431e-13
L_PTL_IG2_0|_RX|P3 _PTL_IG2_0|_RX|8 0  5.339e-13
R_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|101  4.225701121488
R_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|104  3.429952209
R_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|107  2.7439617672
L_PTL_IG2_0|_RX|RB1 _PTL_IG2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG2_0|_RX|RB2 _PTL_IG2_0|_RX|104 0  1.937922998085e-12
L_PTL_IG2_0|_RX|RB3 _PTL_IG2_0|_RX|107 0  1.550338398468e-12
B_PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_0|_TX|B1 0 _PTL_IP3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_0|_TX|B2 0 _PTL_IP3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|3  1.684e-12
L_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|6  3.596e-12
L_PTL_IP3_0|_TX|1 IP3_0 _PTL_IP3_0|_TX|1  2.063e-12
L_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|4  4.123e-12
L_PTL_IP3_0|_TX|3 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|7  2.193e-12
R_PTL_IP3_0|_TX|D _PTL_IP3_0|_TX|7 _PTL_IP3_0|A_PTL  1.36
L_PTL_IP3_0|_TX|P1 _PTL_IP3_0|_TX|2 0  5.254e-13
L_PTL_IP3_0|_TX|P2 _PTL_IP3_0|_TX|5 0  5.141e-13
R_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|101  2.7439617672
R_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|104  2.7439617672
L_PTL_IP3_0|_TX|RB1 _PTL_IP3_0|_TX|101 0  1.550338398468e-12
L_PTL_IP3_0|_TX|RB2 _PTL_IP3_0|_TX|104 0  1.550338398468e-12
B_PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_0|_RX|B1 0 _PTL_IP3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|3  2.777e-12
I_PTL_IP3_0|_RX|B2 0 _PTL_IP3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|6  2.685e-12
I_PTL_IP3_0|_RX|B3 0 _PTL_IP3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|9  2.764e-12
L_PTL_IP3_0|_RX|1 _PTL_IP3_0|A_PTL _PTL_IP3_0|_RX|1  1.346e-12
L_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|4  6.348e-12
L_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7  5.197e-12
L_PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7 IP3_0_RX  2.058e-12
L_PTL_IP3_0|_RX|P1 _PTL_IP3_0|_RX|2 0  4.795e-13
L_PTL_IP3_0|_RX|P2 _PTL_IP3_0|_RX|5 0  5.431e-13
L_PTL_IP3_0|_RX|P3 _PTL_IP3_0|_RX|8 0  5.339e-13
R_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|101  4.225701121488
R_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|104  3.429952209
R_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|107  2.7439617672
L_PTL_IP3_0|_RX|RB1 _PTL_IP3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_0|_RX|RB2 _PTL_IP3_0|_RX|104 0  1.937922998085e-12
L_PTL_IP3_0|_RX|RB3 _PTL_IP3_0|_RX|107 0  1.550338398468e-12
B_PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG3_0|_TX|B1 0 _PTL_IG3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG3_0|_TX|B2 0 _PTL_IG3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|3  1.684e-12
L_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|6  3.596e-12
L_PTL_IG3_0|_TX|1 IG3_0 _PTL_IG3_0|_TX|1  2.063e-12
L_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|4  4.123e-12
L_PTL_IG3_0|_TX|3 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|7  2.193e-12
R_PTL_IG3_0|_TX|D _PTL_IG3_0|_TX|7 _PTL_IG3_0|A_PTL  1.36
L_PTL_IG3_0|_TX|P1 _PTL_IG3_0|_TX|2 0  5.254e-13
L_PTL_IG3_0|_TX|P2 _PTL_IG3_0|_TX|5 0  5.141e-13
R_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|101  2.7439617672
R_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|104  2.7439617672
L_PTL_IG3_0|_TX|RB1 _PTL_IG3_0|_TX|101 0  1.550338398468e-12
L_PTL_IG3_0|_TX|RB2 _PTL_IG3_0|_TX|104 0  1.550338398468e-12
B_PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG3_0|_RX|B1 0 _PTL_IG3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|3  2.777e-12
I_PTL_IG3_0|_RX|B2 0 _PTL_IG3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|6  2.685e-12
I_PTL_IG3_0|_RX|B3 0 _PTL_IG3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|9  2.764e-12
L_PTL_IG3_0|_RX|1 _PTL_IG3_0|A_PTL _PTL_IG3_0|_RX|1  1.346e-12
L_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|4  6.348e-12
L_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7  5.197e-12
L_PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7 IG3_0_RX  2.058e-12
L_PTL_IG3_0|_RX|P1 _PTL_IG3_0|_RX|2 0  4.795e-13
L_PTL_IG3_0|_RX|P2 _PTL_IG3_0|_RX|5 0  5.431e-13
L_PTL_IG3_0|_RX|P3 _PTL_IG3_0|_RX|8 0  5.339e-13
R_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|101  4.225701121488
R_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|104  3.429952209
R_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|107  2.7439617672
L_PTL_IG3_0|_RX|RB1 _PTL_IG3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG3_0|_RX|RB2 _PTL_IG3_0|_RX|104 0  1.937922998085e-12
L_PTL_IG3_0|_RX|RB3 _PTL_IG3_0|_RX|107 0  1.550338398468e-12
LSPL_IG0_0|I_D1|B SPL_IG0_0|D1 SPL_IG0_0|I_D1|MID  2e-12
ISPL_IG0_0|I_D1|B 0 SPL_IG0_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_D2|B SPL_IG0_0|D2 SPL_IG0_0|I_D2|MID  2e-12
ISPL_IG0_0|I_D2|B 0 SPL_IG0_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG0_0|I_Q1|B SPL_IG0_0|QA1 SPL_IG0_0|I_Q1|MID  2e-12
ISPL_IG0_0|I_Q1|B 0 SPL_IG0_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_Q2|B SPL_IG0_0|QB1 SPL_IG0_0|I_Q2|MID  2e-12
ISPL_IG0_0|I_Q2|B 0 SPL_IG0_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG0_0|1|1 SPL_IG0_0|D1 SPL_IG0_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|1|P SPL_IG0_0|1|MID_SERIES 0  2e-13
RSPL_IG0_0|1|B SPL_IG0_0|D1 SPL_IG0_0|1|MID_SHUNT  2.7439617672
LSPL_IG0_0|1|RB SPL_IG0_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|2|1 SPL_IG0_0|D2 SPL_IG0_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|2|P SPL_IG0_0|2|MID_SERIES 0  2e-13
RSPL_IG0_0|2|B SPL_IG0_0|D2 SPL_IG0_0|2|MID_SHUNT  2.7439617672
LSPL_IG0_0|2|RB SPL_IG0_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|A|1 SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|A|P SPL_IG0_0|A|MID_SERIES 0  2e-13
RSPL_IG0_0|A|B SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SHUNT  2.7439617672
LSPL_IG0_0|A|RB SPL_IG0_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|B|1 SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|B|P SPL_IG0_0|B|MID_SERIES 0  2e-13
RSPL_IG0_0|B|B SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SHUNT  2.7439617672
LSPL_IG0_0|B|RB SPL_IG0_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP1_0|I_D1|B SPL_IP1_0|D1 SPL_IP1_0|I_D1|MID  2e-12
ISPL_IP1_0|I_D1|B 0 SPL_IP1_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_D2|B SPL_IP1_0|D2 SPL_IP1_0|I_D2|MID  2e-12
ISPL_IP1_0|I_D2|B 0 SPL_IP1_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP1_0|I_Q1|B SPL_IP1_0|QA1 SPL_IP1_0|I_Q1|MID  2e-12
ISPL_IP1_0|I_Q1|B 0 SPL_IP1_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_Q2|B SPL_IP1_0|QB1 SPL_IP1_0|I_Q2|MID  2e-12
ISPL_IP1_0|I_Q2|B 0 SPL_IP1_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP1_0|1|1 SPL_IP1_0|D1 SPL_IP1_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|1|P SPL_IP1_0|1|MID_SERIES 0  2e-13
RSPL_IP1_0|1|B SPL_IP1_0|D1 SPL_IP1_0|1|MID_SHUNT  2.7439617672
LSPL_IP1_0|1|RB SPL_IP1_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|2|1 SPL_IP1_0|D2 SPL_IP1_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|2|P SPL_IP1_0|2|MID_SERIES 0  2e-13
RSPL_IP1_0|2|B SPL_IP1_0|D2 SPL_IP1_0|2|MID_SHUNT  2.7439617672
LSPL_IP1_0|2|RB SPL_IP1_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|A|1 SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|A|P SPL_IP1_0|A|MID_SERIES 0  2e-13
RSPL_IP1_0|A|B SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SHUNT  2.7439617672
LSPL_IP1_0|A|RB SPL_IP1_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|B|1 SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|B|P SPL_IP1_0|B|MID_SERIES 0  2e-13
RSPL_IP1_0|B|B SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SHUNT  2.7439617672
LSPL_IP1_0|B|RB SPL_IP1_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|1 IP2_0_RX SPL_IP2_0|SPL1|D1  2e-12
LSPL_IP2_0|SPL1|2 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|D2  4.135667696e-12
LSPL_IP2_0|SPL1|3 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL1|4 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL1|5 SPL_IP2_0|SPL1|QA1 IP2_0_TO2  2e-12
LSPL_IP2_0|SPL1|6 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL1|7 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|QTMP  2e-12
LSPL_IP2_0|SPL2|1 SPL_IP2_0|QTMP SPL_IP2_0|SPL2|D1  2e-12
LSPL_IP2_0|SPL2|2 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|D2  4.135667696e-12
LSPL_IP2_0|SPL2|3 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL2|4 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL2|5 SPL_IP2_0|SPL2|QA1 IP2_0_TO3  2e-12
LSPL_IP2_0|SPL2|6 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL2|7 SPL_IP2_0|SPL2|QB1 IP2_0_OUT  2e-12
LSPL_IG2_0|I_D1|B SPL_IG2_0|D1 SPL_IG2_0|I_D1|MID  2e-12
ISPL_IG2_0|I_D1|B 0 SPL_IG2_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_D2|B SPL_IG2_0|D2 SPL_IG2_0|I_D2|MID  2e-12
ISPL_IG2_0|I_D2|B 0 SPL_IG2_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG2_0|I_Q1|B SPL_IG2_0|QA1 SPL_IG2_0|I_Q1|MID  2e-12
ISPL_IG2_0|I_Q1|B 0 SPL_IG2_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_Q2|B SPL_IG2_0|QB1 SPL_IG2_0|I_Q2|MID  2e-12
ISPL_IG2_0|I_Q2|B 0 SPL_IG2_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG2_0|1|1 SPL_IG2_0|D1 SPL_IG2_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|1|P SPL_IG2_0|1|MID_SERIES 0  2e-13
RSPL_IG2_0|1|B SPL_IG2_0|D1 SPL_IG2_0|1|MID_SHUNT  2.7439617672
LSPL_IG2_0|1|RB SPL_IG2_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|2|1 SPL_IG2_0|D2 SPL_IG2_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|2|P SPL_IG2_0|2|MID_SERIES 0  2e-13
RSPL_IG2_0|2|B SPL_IG2_0|D2 SPL_IG2_0|2|MID_SHUNT  2.7439617672
LSPL_IG2_0|2|RB SPL_IG2_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|A|1 SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|A|P SPL_IG2_0|A|MID_SERIES 0  2e-13
RSPL_IG2_0|A|B SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SHUNT  2.7439617672
LSPL_IG2_0|A|RB SPL_IG2_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|B|1 SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|B|P SPL_IG2_0|B|MID_SERIES 0  2e-13
RSPL_IG2_0|B|B SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SHUNT  2.7439617672
LSPL_IG2_0|B|RB SPL_IG2_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP3_0|I_D1|B SPL_IP3_0|D1 SPL_IP3_0|I_D1|MID  2e-12
ISPL_IP3_0|I_D1|B 0 SPL_IP3_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_D2|B SPL_IP3_0|D2 SPL_IP3_0|I_D2|MID  2e-12
ISPL_IP3_0|I_D2|B 0 SPL_IP3_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP3_0|I_Q1|B SPL_IP3_0|QA1 SPL_IP3_0|I_Q1|MID  2e-12
ISPL_IP3_0|I_Q1|B 0 SPL_IP3_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_Q2|B SPL_IP3_0|QB1 SPL_IP3_0|I_Q2|MID  2e-12
ISPL_IP3_0|I_Q2|B 0 SPL_IP3_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP3_0|1|1 SPL_IP3_0|D1 SPL_IP3_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|1|P SPL_IP3_0|1|MID_SERIES 0  2e-13
RSPL_IP3_0|1|B SPL_IP3_0|D1 SPL_IP3_0|1|MID_SHUNT  2.7439617672
LSPL_IP3_0|1|RB SPL_IP3_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|2|1 SPL_IP3_0|D2 SPL_IP3_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|2|P SPL_IP3_0|2|MID_SERIES 0  2e-13
RSPL_IP3_0|2|B SPL_IP3_0|D2 SPL_IP3_0|2|MID_SHUNT  2.7439617672
LSPL_IP3_0|2|RB SPL_IP3_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|A|1 SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|A|P SPL_IP3_0|A|MID_SERIES 0  2e-13
RSPL_IP3_0|A|B SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SHUNT  2.7439617672
LSPL_IP3_0|A|RB SPL_IP3_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|B|1 SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|B|P SPL_IP3_0|B|MID_SERIES 0  2e-13
RSPL_IP3_0|B|B SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SHUNT  2.7439617672
LSPL_IP3_0|B|RB SPL_IP3_0|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|1 IP0_0_RX _PG0_01|P|A1  2.067833848e-12
L_PG0_01|P|2 _PG0_01|P|A1 _PG0_01|P|A2  4.135667696e-12
L_PG0_01|P|3 _PG0_01|P|A3 _PG0_01|P|A4  8.271335392e-12
L_PG0_01|P|T T04 _PG0_01|P|T1  2.067833848e-12
L_PG0_01|P|4 _PG0_01|P|T1 _PG0_01|P|T2  4.135667696e-12
L_PG0_01|P|5 _PG0_01|P|A4 _PG0_01|P|Q1  4.135667696e-12
L_PG0_01|P|6 _PG0_01|P|Q1 P0_1  2.067833848e-12
L_PG0_01|G|1 IG0_0_TO0 _PG0_01|G|A1  2.067833848e-12
L_PG0_01|G|2 _PG0_01|G|A1 _PG0_01|G|A2  4.135667696e-12
L_PG0_01|G|3 _PG0_01|G|A3 _PG0_01|G|A4  8.271335392e-12
L_PG0_01|G|T T04 _PG0_01|G|T1  2.067833848e-12
L_PG0_01|G|4 _PG0_01|G|T1 _PG0_01|G|T2  4.135667696e-12
L_PG0_01|G|5 _PG0_01|G|A4 _PG0_01|G|Q1  4.135667696e-12
L_PG0_01|G|6 _PG0_01|G|Q1 G0_1  2.067833848e-12
L_PG1_01|_SPL_G1|1 IG1_0_RX _PG1_01|_SPL_G1|D1  2e-12
L_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|D2  4.135667696e-12
L_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG1_01|_SPL_G1|5 _PG1_01|_SPL_G1|QA1 _PG1_01|G1_COPY_1  2e-12
L_PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|QB1 _PG1_01|G1_COPY_2  2e-12
L_PG1_01|_PG|A1 IP1_0_TO1 _PG1_01|_PG|A1  2.067833848e-12
L_PG1_01|_PG|A2 _PG1_01|_PG|A1 _PG1_01|_PG|A2  4.135667696e-12
L_PG1_01|_PG|A3 _PG1_01|_PG|A3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|B1 _PG1_01|G1_COPY_1 _PG1_01|_PG|B1  2.067833848e-12
L_PG1_01|_PG|B2 _PG1_01|_PG|B1 _PG1_01|_PG|B2  4.135667696e-12
L_PG1_01|_PG|B3 _PG1_01|_PG|B3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|Q3 _PG1_01|_PG|Q3 _PG1_01|_PG|Q2  4.135667696e-12
L_PG1_01|_PG|Q2 _PG1_01|_PG|Q2 _PG1_01|_PG|Q1  4.135667696e-12
L_PG1_01|_PG|Q1 _PG1_01|_PG|Q1 _PG1_01|PG  2.067833848e-12
L_PG1_01|_GG|A1 IG0_0_TO1 _PG1_01|_GG|A1  2.067833848e-12
L_PG1_01|_GG|A2 _PG1_01|_GG|A1 _PG1_01|_GG|A2  4.135667696e-12
L_PG1_01|_GG|A3 _PG1_01|_GG|A3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|B1 _PG1_01|G1_COPY_2 _PG1_01|_GG|B1  2.067833848e-12
L_PG1_01|_GG|B2 _PG1_01|_GG|B1 _PG1_01|_GG|B2  4.135667696e-12
L_PG1_01|_GG|B3 _PG1_01|_GG|B3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|Q3 _PG1_01|_GG|Q3 _PG1_01|_GG|Q2  4.135667696e-12
L_PG1_01|_GG|Q2 _PG1_01|_GG|Q2 _PG1_01|_GG|Q1  4.135667696e-12
L_PG1_01|_GG|Q1 _PG1_01|_GG|Q1 _PG1_01|GG  2.067833848e-12
L_PG1_01|_DFF_PG|1 _PG1_01|PG _PG1_01|_DFF_PG|A1  2.067833848e-12
L_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|A2  4.135667696e-12
L_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|A4  8.271335392e-12
L_PG1_01|_DFF_PG|T T05 _PG1_01|_DFF_PG|T1  2.067833848e-12
L_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T2  4.135667696e-12
L_PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|Q1  4.135667696e-12
L_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|Q1 _PG1_01|PG_SYNC  2.067833848e-12
L_PG1_01|_DFF_GG|1 _PG1_01|GG _PG1_01|_DFF_GG|A1  2.067833848e-12
L_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|A2  4.135667696e-12
L_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|A4  8.271335392e-12
L_PG1_01|_DFF_GG|T T05 _PG1_01|_DFF_GG|T1  2.067833848e-12
L_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T2  4.135667696e-12
L_PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|Q1  4.135667696e-12
L_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|Q1 _PG1_01|GG_SYNC  2.067833848e-12
L_PG1_01|_AND_G|A1 _PG1_01|PG_SYNC _PG1_01|_AND_G|A1  2.067833848e-12
L_PG1_01|_AND_G|A2 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A2  4.135667696e-12
L_PG1_01|_AND_G|A3 _PG1_01|_AND_G|A3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|B1 _PG1_01|GG_SYNC _PG1_01|_AND_G|B1  2.067833848e-12
L_PG1_01|_AND_G|B2 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B2  4.135667696e-12
L_PG1_01|_AND_G|B3 _PG1_01|_AND_G|B3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q2  4.135667696e-12
L_PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q1  4.135667696e-12
L_PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1 G1_1  2.067833848e-12
L_PG2_01|P|1 IP2_0_TO2 _PG2_01|P|A1  2.067833848e-12
L_PG2_01|P|2 _PG2_01|P|A1 _PG2_01|P|A2  4.135667696e-12
L_PG2_01|P|3 _PG2_01|P|A3 _PG2_01|P|A4  8.271335392e-12
L_PG2_01|P|T T06 _PG2_01|P|T1  2.067833848e-12
L_PG2_01|P|4 _PG2_01|P|T1 _PG2_01|P|T2  4.135667696e-12
L_PG2_01|P|5 _PG2_01|P|A4 _PG2_01|P|Q1  4.135667696e-12
L_PG2_01|P|6 _PG2_01|P|Q1 P2_1  2.067833848e-12
L_PG2_01|G|1 IG2_0_TO2 _PG2_01|G|A1  2.067833848e-12
L_PG2_01|G|2 _PG2_01|G|A1 _PG2_01|G|A2  4.135667696e-12
L_PG2_01|G|3 _PG2_01|G|A3 _PG2_01|G|A4  8.271335392e-12
L_PG2_01|G|T T06 _PG2_01|G|T1  2.067833848e-12
L_PG2_01|G|4 _PG2_01|G|T1 _PG2_01|G|T2  4.135667696e-12
L_PG2_01|G|5 _PG2_01|G|A4 _PG2_01|G|Q1  4.135667696e-12
L_PG2_01|G|6 _PG2_01|G|Q1 G2_1  2.067833848e-12
L_PG3_01|_SPL_G1|1 IG3_0_RX _PG3_01|_SPL_G1|D1  2e-12
L_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|D2  4.135667696e-12
L_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_G1|5 _PG3_01|_SPL_G1|QA1 _PG3_01|G1_COPY_1  2e-12
L_PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|QB1 _PG3_01|G1_COPY_2  2e-12
L_PG3_01|_SPL_P1|1 IP3_0_TO1 _PG3_01|_SPL_P1|D1  2e-12
L_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|D2  4.135667696e-12
L_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_P1|5 _PG3_01|_SPL_P1|QA1 _PG3_01|P1_COPY_1  2e-12
L_PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|QB1 _PG3_01|P1_COPY_2  2e-12
L_PG3_01|_PG|A1 _PG3_01|P1_COPY_1 _PG3_01|_PG|A1  2.067833848e-12
L_PG3_01|_PG|A2 _PG3_01|_PG|A1 _PG3_01|_PG|A2  4.135667696e-12
L_PG3_01|_PG|A3 _PG3_01|_PG|A3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|B1 _PG3_01|G1_COPY_1 _PG3_01|_PG|B1  2.067833848e-12
L_PG3_01|_PG|B2 _PG3_01|_PG|B1 _PG3_01|_PG|B2  4.135667696e-12
L_PG3_01|_PG|B3 _PG3_01|_PG|B3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|Q3 _PG3_01|_PG|Q3 _PG3_01|_PG|Q2  4.135667696e-12
L_PG3_01|_PG|Q2 _PG3_01|_PG|Q2 _PG3_01|_PG|Q1  4.135667696e-12
L_PG3_01|_PG|Q1 _PG3_01|_PG|Q1 _PG3_01|PG  2.067833848e-12
L_PG3_01|_GG|A1 IG2_0_TO3 _PG3_01|_GG|A1  2.067833848e-12
L_PG3_01|_GG|A2 _PG3_01|_GG|A1 _PG3_01|_GG|A2  4.135667696e-12
L_PG3_01|_GG|A3 _PG3_01|_GG|A3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|B1 _PG3_01|G1_COPY_2 _PG3_01|_GG|B1  2.067833848e-12
L_PG3_01|_GG|B2 _PG3_01|_GG|B1 _PG3_01|_GG|B2  4.135667696e-12
L_PG3_01|_GG|B3 _PG3_01|_GG|B3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|Q3 _PG3_01|_GG|Q3 _PG3_01|_GG|Q2  4.135667696e-12
L_PG3_01|_GG|Q2 _PG3_01|_GG|Q2 _PG3_01|_GG|Q1  4.135667696e-12
L_PG3_01|_GG|Q1 _PG3_01|_GG|Q1 _PG3_01|GG  2.067833848e-12
L_PG3_01|_DFF_P0|1 IP2_0_TO3 _PG3_01|_DFF_P0|A1  2.067833848e-12
L_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|A2  4.135667696e-12
L_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|A4  8.271335392e-12
L_PG3_01|_DFF_P0|T T07 _PG3_01|_DFF_P0|T1  2.067833848e-12
L_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T2  4.135667696e-12
L_PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|Q1  4.135667696e-12
L_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|Q1 _PG3_01|P0_SYNC  2.067833848e-12
L_PG3_01|_DFF_P1|1 _PG3_01|P1_COPY_2 _PG3_01|_DFF_P1|A1  2.067833848e-12
L_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|A2  4.135667696e-12
L_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|A4  8.271335392e-12
L_PG3_01|_DFF_P1|T T07 _PG3_01|_DFF_P1|T1  2.067833848e-12
L_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T2  4.135667696e-12
L_PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|Q1  4.135667696e-12
L_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|Q1 _PG3_01|P1_SYNC  2.067833848e-12
L_PG3_01|_DFF_PG|1 _PG3_01|PG _PG3_01|_DFF_PG|A1  2.067833848e-12
L_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|A2  4.135667696e-12
L_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|A4  8.271335392e-12
L_PG3_01|_DFF_PG|T T07 _PG3_01|_DFF_PG|T1  2.067833848e-12
L_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T2  4.135667696e-12
L_PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|Q1  4.135667696e-12
L_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|Q1 _PG3_01|PG_SYNC  2.067833848e-12
L_PG3_01|_DFF_GG|1 _PG3_01|GG _PG3_01|_DFF_GG|A1  2.067833848e-12
L_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|A2  4.135667696e-12
L_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|A4  8.271335392e-12
L_PG3_01|_DFF_GG|T T07 _PG3_01|_DFF_GG|T1  2.067833848e-12
L_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T2  4.135667696e-12
L_PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|Q1  4.135667696e-12
L_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|Q1 _PG3_01|GG_SYNC  2.067833848e-12
L_PG3_01|_AND_G|A1 _PG3_01|PG_SYNC _PG3_01|_AND_G|A1  2.067833848e-12
L_PG3_01|_AND_G|A2 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A2  4.135667696e-12
L_PG3_01|_AND_G|A3 _PG3_01|_AND_G|A3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|B1 _PG3_01|GG_SYNC _PG3_01|_AND_G|B1  2.067833848e-12
L_PG3_01|_AND_G|B2 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B2  4.135667696e-12
L_PG3_01|_AND_G|B3 _PG3_01|_AND_G|B3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q2  4.135667696e-12
L_PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q1  4.135667696e-12
L_PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1 G3_1  2.067833848e-12
L_PG3_01|_AND_P|A1 _PG3_01|P0_SYNC _PG3_01|_AND_P|A1  2.067833848e-12
L_PG3_01|_AND_P|A2 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A2  4.135667696e-12
L_PG3_01|_AND_P|A3 _PG3_01|_AND_P|A3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|B1 _PG3_01|P1_SYNC _PG3_01|_AND_P|B1  2.067833848e-12
L_PG3_01|_AND_P|B2 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B2  4.135667696e-12
L_PG3_01|_AND_P|B3 _PG3_01|_AND_P|B3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q2  4.135667696e-12
L_PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q1  4.135667696e-12
L_PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1 P3_1  2.067833848e-12
L_DFF_IP1_01|I_1|B _DFF_IP1_01|A1 _DFF_IP1_01|I_1|MID  2e-12
I_DFF_IP1_01|I_1|B 0 _DFF_IP1_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_3|B _DFF_IP1_01|A3 _DFF_IP1_01|I_3|MID  2e-12
I_DFF_IP1_01|I_3|B 0 _DFF_IP1_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_01|I_T|B _DFF_IP1_01|T1 _DFF_IP1_01|I_T|MID  2e-12
I_DFF_IP1_01|I_T|B 0 _DFF_IP1_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_6|B _DFF_IP1_01|Q1 _DFF_IP1_01|I_6|MID  2e-12
I_DFF_IP1_01|I_6|B 0 _DFF_IP1_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_01|1|1 _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|1|P _DFF_IP1_01|1|MID_SERIES 0  2e-13
R_DFF_IP1_01|1|B _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SHUNT  2.7439617672
L_DFF_IP1_01|1|RB _DFF_IP1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|23|1 _DFF_IP1_01|A2 _DFF_IP1_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|23|B _DFF_IP1_01|A2 _DFF_IP1_01|23|MID_SHUNT  3.84154647408
L_DFF_IP1_01|23|RB _DFF_IP1_01|23|MID_SHUNT _DFF_IP1_01|A3  2.1704737578552e-12
B_DFF_IP1_01|3|1 _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|3|P _DFF_IP1_01|3|MID_SERIES 0  2e-13
R_DFF_IP1_01|3|B _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SHUNT  2.7439617672
L_DFF_IP1_01|3|RB _DFF_IP1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|4|1 _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|4|P _DFF_IP1_01|4|MID_SERIES 0  2e-13
R_DFF_IP1_01|4|B _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SHUNT  2.7439617672
L_DFF_IP1_01|4|RB _DFF_IP1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|T|1 _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|T|P _DFF_IP1_01|T|MID_SERIES 0  2e-13
R_DFF_IP1_01|T|B _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SHUNT  2.7439617672
L_DFF_IP1_01|T|RB _DFF_IP1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|45|1 _DFF_IP1_01|T2 _DFF_IP1_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|45|B _DFF_IP1_01|T2 _DFF_IP1_01|45|MID_SHUNT  3.84154647408
L_DFF_IP1_01|45|RB _DFF_IP1_01|45|MID_SHUNT _DFF_IP1_01|A4  2.1704737578552e-12
B_DFF_IP1_01|6|1 _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|6|P _DFF_IP1_01|6|MID_SERIES 0  2e-13
R_DFF_IP1_01|6|B _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SHUNT  2.7439617672
L_DFF_IP1_01|6|RB _DFF_IP1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_01|I_1|B _DFF_IP2_01|A1 _DFF_IP2_01|I_1|MID  2e-12
I_DFF_IP2_01|I_1|B 0 _DFF_IP2_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_3|B _DFF_IP2_01|A3 _DFF_IP2_01|I_3|MID  2e-12
I_DFF_IP2_01|I_3|B 0 _DFF_IP2_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_01|I_T|B _DFF_IP2_01|T1 _DFF_IP2_01|I_T|MID  2e-12
I_DFF_IP2_01|I_T|B 0 _DFF_IP2_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_6|B _DFF_IP2_01|Q1 _DFF_IP2_01|I_6|MID  2e-12
I_DFF_IP2_01|I_6|B 0 _DFF_IP2_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_01|1|1 _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|1|P _DFF_IP2_01|1|MID_SERIES 0  2e-13
R_DFF_IP2_01|1|B _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SHUNT  2.7439617672
L_DFF_IP2_01|1|RB _DFF_IP2_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|23|1 _DFF_IP2_01|A2 _DFF_IP2_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|23|B _DFF_IP2_01|A2 _DFF_IP2_01|23|MID_SHUNT  3.84154647408
L_DFF_IP2_01|23|RB _DFF_IP2_01|23|MID_SHUNT _DFF_IP2_01|A3  2.1704737578552e-12
B_DFF_IP2_01|3|1 _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|3|P _DFF_IP2_01|3|MID_SERIES 0  2e-13
R_DFF_IP2_01|3|B _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SHUNT  2.7439617672
L_DFF_IP2_01|3|RB _DFF_IP2_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|4|1 _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|4|P _DFF_IP2_01|4|MID_SERIES 0  2e-13
R_DFF_IP2_01|4|B _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SHUNT  2.7439617672
L_DFF_IP2_01|4|RB _DFF_IP2_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|T|1 _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|T|P _DFF_IP2_01|T|MID_SERIES 0  2e-13
R_DFF_IP2_01|T|B _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SHUNT  2.7439617672
L_DFF_IP2_01|T|RB _DFF_IP2_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|45|1 _DFF_IP2_01|T2 _DFF_IP2_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|45|B _DFF_IP2_01|T2 _DFF_IP2_01|45|MID_SHUNT  3.84154647408
L_DFF_IP2_01|45|RB _DFF_IP2_01|45|MID_SHUNT _DFF_IP2_01|A4  2.1704737578552e-12
B_DFF_IP2_01|6|1 _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|6|P _DFF_IP2_01|6|MID_SERIES 0  2e-13
R_DFF_IP2_01|6|B _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SHUNT  2.7439617672
L_DFF_IP2_01|6|RB _DFF_IP2_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_01|I_1|B _DFF_IP3_01|A1 _DFF_IP3_01|I_1|MID  2e-12
I_DFF_IP3_01|I_1|B 0 _DFF_IP3_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_3|B _DFF_IP3_01|A3 _DFF_IP3_01|I_3|MID  2e-12
I_DFF_IP3_01|I_3|B 0 _DFF_IP3_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_01|I_T|B _DFF_IP3_01|T1 _DFF_IP3_01|I_T|MID  2e-12
I_DFF_IP3_01|I_T|B 0 _DFF_IP3_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_6|B _DFF_IP3_01|Q1 _DFF_IP3_01|I_6|MID  2e-12
I_DFF_IP3_01|I_6|B 0 _DFF_IP3_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_01|1|1 _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|1|P _DFF_IP3_01|1|MID_SERIES 0  2e-13
R_DFF_IP3_01|1|B _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SHUNT  2.7439617672
L_DFF_IP3_01|1|RB _DFF_IP3_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|23|1 _DFF_IP3_01|A2 _DFF_IP3_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|23|B _DFF_IP3_01|A2 _DFF_IP3_01|23|MID_SHUNT  3.84154647408
L_DFF_IP3_01|23|RB _DFF_IP3_01|23|MID_SHUNT _DFF_IP3_01|A3  2.1704737578552e-12
B_DFF_IP3_01|3|1 _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|3|P _DFF_IP3_01|3|MID_SERIES 0  2e-13
R_DFF_IP3_01|3|B _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SHUNT  2.7439617672
L_DFF_IP3_01|3|RB _DFF_IP3_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|4|1 _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|4|P _DFF_IP3_01|4|MID_SERIES 0  2e-13
R_DFF_IP3_01|4|B _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SHUNT  2.7439617672
L_DFF_IP3_01|4|RB _DFF_IP3_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|T|1 _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|T|P _DFF_IP3_01|T|MID_SERIES 0  2e-13
R_DFF_IP3_01|T|B _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SHUNT  2.7439617672
L_DFF_IP3_01|T|RB _DFF_IP3_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|45|1 _DFF_IP3_01|T2 _DFF_IP3_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|45|B _DFF_IP3_01|T2 _DFF_IP3_01|45|MID_SHUNT  3.84154647408
L_DFF_IP3_01|45|RB _DFF_IP3_01|45|MID_SHUNT _DFF_IP3_01|A4  2.1704737578552e-12
B_DFF_IP3_01|6|1 _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|6|P _DFF_IP3_01|6|MID_SERIES 0  2e-13
R_DFF_IP3_01|6|B _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SHUNT  2.7439617672
L_DFF_IP3_01|6|RB _DFF_IP3_01|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_P0_1|_TX|1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|2 JJMIT AREA=2.5
B_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|5 JJMIT AREA=2.5
I_PTL_P0_1|_TX|B1 0 _PTL_P0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_1|_TX|B2 0 _PTL_P0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|3  1.684e-12
L_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|6  3.596e-12
L_PTL_P0_1|_TX|1 P0_1 _PTL_P0_1|_TX|1  2.063e-12
L_PTL_P0_1|_TX|2 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|4  4.123e-12
L_PTL_P0_1|_TX|3 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|7  2.193e-12
R_PTL_P0_1|_TX|D _PTL_P0_1|_TX|7 _PTL_P0_1|A_PTL  1.36
L_PTL_P0_1|_TX|P1 _PTL_P0_1|_TX|2 0  5.254e-13
L_PTL_P0_1|_TX|P2 _PTL_P0_1|_TX|5 0  5.141e-13
R_PTL_P0_1|_TX|B1 _PTL_P0_1|_TX|1 _PTL_P0_1|_TX|101  2.7439617672
R_PTL_P0_1|_TX|B2 _PTL_P0_1|_TX|4 _PTL_P0_1|_TX|104  2.7439617672
L_PTL_P0_1|_TX|RB1 _PTL_P0_1|_TX|101 0  1.550338398468e-12
L_PTL_P0_1|_TX|RB2 _PTL_P0_1|_TX|104 0  1.550338398468e-12
B_PTL_P0_1|_RX|1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|5 JJMIT AREA=2.0
B_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|8 JJMIT AREA=2.5
I_PTL_P0_1|_RX|B1 0 _PTL_P0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|3  2.777e-12
I_PTL_P0_1|_RX|B2 0 _PTL_P0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|6  2.685e-12
I_PTL_P0_1|_RX|B3 0 _PTL_P0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|9  2.764e-12
L_PTL_P0_1|_RX|1 _PTL_P0_1|A_PTL _PTL_P0_1|_RX|1  1.346e-12
L_PTL_P0_1|_RX|2 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|4  6.348e-12
L_PTL_P0_1|_RX|3 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7  5.197e-12
L_PTL_P0_1|_RX|4 _PTL_P0_1|_RX|7 P0_1_RX  2.058e-12
L_PTL_P0_1|_RX|P1 _PTL_P0_1|_RX|2 0  4.795e-13
L_PTL_P0_1|_RX|P2 _PTL_P0_1|_RX|5 0  5.431e-13
L_PTL_P0_1|_RX|P3 _PTL_P0_1|_RX|8 0  5.339e-13
R_PTL_P0_1|_RX|B1 _PTL_P0_1|_RX|1 _PTL_P0_1|_RX|101  4.225701121488
R_PTL_P0_1|_RX|B2 _PTL_P0_1|_RX|4 _PTL_P0_1|_RX|104  3.429952209
R_PTL_P0_1|_RX|B3 _PTL_P0_1|_RX|7 _PTL_P0_1|_RX|107  2.7439617672
L_PTL_P0_1|_RX|RB1 _PTL_P0_1|_RX|101 0  2.38752113364072e-12
L_PTL_P0_1|_RX|RB2 _PTL_P0_1|_RX|104 0  1.937922998085e-12
L_PTL_P0_1|_RX|RB3 _PTL_P0_1|_RX|107 0  1.550338398468e-12
B_PTL_G0_1|_TX|1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|2 JJMIT AREA=2.5
B_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|5 JJMIT AREA=2.5
I_PTL_G0_1|_TX|B1 0 _PTL_G0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_1|_TX|B2 0 _PTL_G0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|3  1.684e-12
L_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|6  3.596e-12
L_PTL_G0_1|_TX|1 G0_1 _PTL_G0_1|_TX|1  2.063e-12
L_PTL_G0_1|_TX|2 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|4  4.123e-12
L_PTL_G0_1|_TX|3 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|7  2.193e-12
R_PTL_G0_1|_TX|D _PTL_G0_1|_TX|7 _PTL_G0_1|A_PTL  1.36
L_PTL_G0_1|_TX|P1 _PTL_G0_1|_TX|2 0  5.254e-13
L_PTL_G0_1|_TX|P2 _PTL_G0_1|_TX|5 0  5.141e-13
R_PTL_G0_1|_TX|B1 _PTL_G0_1|_TX|1 _PTL_G0_1|_TX|101  2.7439617672
R_PTL_G0_1|_TX|B2 _PTL_G0_1|_TX|4 _PTL_G0_1|_TX|104  2.7439617672
L_PTL_G0_1|_TX|RB1 _PTL_G0_1|_TX|101 0  1.550338398468e-12
L_PTL_G0_1|_TX|RB2 _PTL_G0_1|_TX|104 0  1.550338398468e-12
B_PTL_G0_1|_RX|1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|5 JJMIT AREA=2.0
B_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|8 JJMIT AREA=2.5
I_PTL_G0_1|_RX|B1 0 _PTL_G0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|3  2.777e-12
I_PTL_G0_1|_RX|B2 0 _PTL_G0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|6  2.685e-12
I_PTL_G0_1|_RX|B3 0 _PTL_G0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|9  2.764e-12
L_PTL_G0_1|_RX|1 _PTL_G0_1|A_PTL _PTL_G0_1|_RX|1  1.346e-12
L_PTL_G0_1|_RX|2 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|4  6.348e-12
L_PTL_G0_1|_RX|3 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7  5.197e-12
L_PTL_G0_1|_RX|4 _PTL_G0_1|_RX|7 G0_1_RX  2.058e-12
L_PTL_G0_1|_RX|P1 _PTL_G0_1|_RX|2 0  4.795e-13
L_PTL_G0_1|_RX|P2 _PTL_G0_1|_RX|5 0  5.431e-13
L_PTL_G0_1|_RX|P3 _PTL_G0_1|_RX|8 0  5.339e-13
R_PTL_G0_1|_RX|B1 _PTL_G0_1|_RX|1 _PTL_G0_1|_RX|101  4.225701121488
R_PTL_G0_1|_RX|B2 _PTL_G0_1|_RX|4 _PTL_G0_1|_RX|104  3.429952209
R_PTL_G0_1|_RX|B3 _PTL_G0_1|_RX|7 _PTL_G0_1|_RX|107  2.7439617672
L_PTL_G0_1|_RX|RB1 _PTL_G0_1|_RX|101 0  2.38752113364072e-12
L_PTL_G0_1|_RX|RB2 _PTL_G0_1|_RX|104 0  1.937922998085e-12
L_PTL_G0_1|_RX|RB3 _PTL_G0_1|_RX|107 0  1.550338398468e-12
B_PTL_G1_1|_TX|1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|2 JJMIT AREA=2.5
B_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|5 JJMIT AREA=2.5
I_PTL_G1_1|_TX|B1 0 _PTL_G1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_1|_TX|B2 0 _PTL_G1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|3  1.684e-12
L_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|6  3.596e-12
L_PTL_G1_1|_TX|1 G1_1 _PTL_G1_1|_TX|1  2.063e-12
L_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|4  4.123e-12
L_PTL_G1_1|_TX|3 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|7  2.193e-12
R_PTL_G1_1|_TX|D _PTL_G1_1|_TX|7 _PTL_G1_1|A_PTL  1.36
L_PTL_G1_1|_TX|P1 _PTL_G1_1|_TX|2 0  5.254e-13
L_PTL_G1_1|_TX|P2 _PTL_G1_1|_TX|5 0  5.141e-13
R_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|101  2.7439617672
R_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|104  2.7439617672
L_PTL_G1_1|_TX|RB1 _PTL_G1_1|_TX|101 0  1.550338398468e-12
L_PTL_G1_1|_TX|RB2 _PTL_G1_1|_TX|104 0  1.550338398468e-12
B_PTL_G1_1|_RX|1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|5 JJMIT AREA=2.0
B_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|8 JJMIT AREA=2.5
I_PTL_G1_1|_RX|B1 0 _PTL_G1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|3  2.777e-12
I_PTL_G1_1|_RX|B2 0 _PTL_G1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|6  2.685e-12
I_PTL_G1_1|_RX|B3 0 _PTL_G1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|9  2.764e-12
L_PTL_G1_1|_RX|1 _PTL_G1_1|A_PTL _PTL_G1_1|_RX|1  1.346e-12
L_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|4  6.348e-12
L_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7  5.197e-12
L_PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7 G1_1_RX  2.058e-12
L_PTL_G1_1|_RX|P1 _PTL_G1_1|_RX|2 0  4.795e-13
L_PTL_G1_1|_RX|P2 _PTL_G1_1|_RX|5 0  5.431e-13
L_PTL_G1_1|_RX|P3 _PTL_G1_1|_RX|8 0  5.339e-13
R_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|101  4.225701121488
R_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|104  3.429952209
R_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|107  2.7439617672
L_PTL_G1_1|_RX|RB1 _PTL_G1_1|_RX|101 0  2.38752113364072e-12
L_PTL_G1_1|_RX|RB2 _PTL_G1_1|_RX|104 0  1.937922998085e-12
L_PTL_G1_1|_RX|RB3 _PTL_G1_1|_RX|107 0  1.550338398468e-12
B_PTL_P2_1|_TX|1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|2 JJMIT AREA=2.5
B_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|5 JJMIT AREA=2.5
I_PTL_P2_1|_TX|B1 0 _PTL_P2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P2_1|_TX|B2 0 _PTL_P2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|3  1.684e-12
L_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|6  3.596e-12
L_PTL_P2_1|_TX|1 P2_1 _PTL_P2_1|_TX|1  2.063e-12
L_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|4  4.123e-12
L_PTL_P2_1|_TX|3 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|7  2.193e-12
R_PTL_P2_1|_TX|D _PTL_P2_1|_TX|7 _PTL_P2_1|A_PTL  1.36
L_PTL_P2_1|_TX|P1 _PTL_P2_1|_TX|2 0  5.254e-13
L_PTL_P2_1|_TX|P2 _PTL_P2_1|_TX|5 0  5.141e-13
R_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|101  2.7439617672
R_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|104  2.7439617672
L_PTL_P2_1|_TX|RB1 _PTL_P2_1|_TX|101 0  1.550338398468e-12
L_PTL_P2_1|_TX|RB2 _PTL_P2_1|_TX|104 0  1.550338398468e-12
B_PTL_P2_1|_RX|1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|5 JJMIT AREA=2.0
B_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|8 JJMIT AREA=2.5
I_PTL_P2_1|_RX|B1 0 _PTL_P2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|3  2.777e-12
I_PTL_P2_1|_RX|B2 0 _PTL_P2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|6  2.685e-12
I_PTL_P2_1|_RX|B3 0 _PTL_P2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|9  2.764e-12
L_PTL_P2_1|_RX|1 _PTL_P2_1|A_PTL _PTL_P2_1|_RX|1  1.346e-12
L_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|4  6.348e-12
L_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7  5.197e-12
L_PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7 P2_1_RX  2.058e-12
L_PTL_P2_1|_RX|P1 _PTL_P2_1|_RX|2 0  4.795e-13
L_PTL_P2_1|_RX|P2 _PTL_P2_1|_RX|5 0  5.431e-13
L_PTL_P2_1|_RX|P3 _PTL_P2_1|_RX|8 0  5.339e-13
R_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|101  4.225701121488
R_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|104  3.429952209
R_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|107  2.7439617672
L_PTL_P2_1|_RX|RB1 _PTL_P2_1|_RX|101 0  2.38752113364072e-12
L_PTL_P2_1|_RX|RB2 _PTL_P2_1|_RX|104 0  1.937922998085e-12
L_PTL_P2_1|_RX|RB3 _PTL_P2_1|_RX|107 0  1.550338398468e-12
B_PTL_G2_1|_TX|1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|2 JJMIT AREA=2.5
B_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|5 JJMIT AREA=2.5
I_PTL_G2_1|_TX|B1 0 _PTL_G2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_1|_TX|B2 0 _PTL_G2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|3  1.684e-12
L_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|6  3.596e-12
L_PTL_G2_1|_TX|1 G2_1 _PTL_G2_1|_TX|1  2.063e-12
L_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|4  4.123e-12
L_PTL_G2_1|_TX|3 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|7  2.193e-12
R_PTL_G2_1|_TX|D _PTL_G2_1|_TX|7 _PTL_G2_1|A_PTL  1.36
L_PTL_G2_1|_TX|P1 _PTL_G2_1|_TX|2 0  5.254e-13
L_PTL_G2_1|_TX|P2 _PTL_G2_1|_TX|5 0  5.141e-13
R_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|101  2.7439617672
R_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|104  2.7439617672
L_PTL_G2_1|_TX|RB1 _PTL_G2_1|_TX|101 0  1.550338398468e-12
L_PTL_G2_1|_TX|RB2 _PTL_G2_1|_TX|104 0  1.550338398468e-12
B_PTL_G2_1|_RX|1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|5 JJMIT AREA=2.0
B_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|8 JJMIT AREA=2.5
I_PTL_G2_1|_RX|B1 0 _PTL_G2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|3  2.777e-12
I_PTL_G2_1|_RX|B2 0 _PTL_G2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|6  2.685e-12
I_PTL_G2_1|_RX|B3 0 _PTL_G2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|9  2.764e-12
L_PTL_G2_1|_RX|1 _PTL_G2_1|A_PTL _PTL_G2_1|_RX|1  1.346e-12
L_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|4  6.348e-12
L_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7  5.197e-12
L_PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7 G2_1_RX  2.058e-12
L_PTL_G2_1|_RX|P1 _PTL_G2_1|_RX|2 0  4.795e-13
L_PTL_G2_1|_RX|P2 _PTL_G2_1|_RX|5 0  5.431e-13
L_PTL_G2_1|_RX|P3 _PTL_G2_1|_RX|8 0  5.339e-13
R_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|101  4.225701121488
R_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|104  3.429952209
R_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|107  2.7439617672
L_PTL_G2_1|_RX|RB1 _PTL_G2_1|_RX|101 0  2.38752113364072e-12
L_PTL_G2_1|_RX|RB2 _PTL_G2_1|_RX|104 0  1.937922998085e-12
L_PTL_G2_1|_RX|RB3 _PTL_G2_1|_RX|107 0  1.550338398468e-12
B_PTL_P3_1|_TX|1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|2 JJMIT AREA=2.5
B_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|5 JJMIT AREA=2.5
I_PTL_P3_1|_TX|B1 0 _PTL_P3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P3_1|_TX|B2 0 _PTL_P3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|3  1.684e-12
L_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|6  3.596e-12
L_PTL_P3_1|_TX|1 P3_1 _PTL_P3_1|_TX|1  2.063e-12
L_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|4  4.123e-12
L_PTL_P3_1|_TX|3 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|7  2.193e-12
R_PTL_P3_1|_TX|D _PTL_P3_1|_TX|7 _PTL_P3_1|A_PTL  1.36
L_PTL_P3_1|_TX|P1 _PTL_P3_1|_TX|2 0  5.254e-13
L_PTL_P3_1|_TX|P2 _PTL_P3_1|_TX|5 0  5.141e-13
R_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|101  2.7439617672
R_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|104  2.7439617672
L_PTL_P3_1|_TX|RB1 _PTL_P3_1|_TX|101 0  1.550338398468e-12
L_PTL_P3_1|_TX|RB2 _PTL_P3_1|_TX|104 0  1.550338398468e-12
B_PTL_P3_1|_RX|1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|5 JJMIT AREA=2.0
B_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|8 JJMIT AREA=2.5
I_PTL_P3_1|_RX|B1 0 _PTL_P3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|3  2.777e-12
I_PTL_P3_1|_RX|B2 0 _PTL_P3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|6  2.685e-12
I_PTL_P3_1|_RX|B3 0 _PTL_P3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|9  2.764e-12
L_PTL_P3_1|_RX|1 _PTL_P3_1|A_PTL _PTL_P3_1|_RX|1  1.346e-12
L_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|4  6.348e-12
L_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7  5.197e-12
L_PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7 P3_1_RX  2.058e-12
L_PTL_P3_1|_RX|P1 _PTL_P3_1|_RX|2 0  4.795e-13
L_PTL_P3_1|_RX|P2 _PTL_P3_1|_RX|5 0  5.431e-13
L_PTL_P3_1|_RX|P3 _PTL_P3_1|_RX|8 0  5.339e-13
R_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|101  4.225701121488
R_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|104  3.429952209
R_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|107  2.7439617672
L_PTL_P3_1|_RX|RB1 _PTL_P3_1|_RX|101 0  2.38752113364072e-12
L_PTL_P3_1|_RX|RB2 _PTL_P3_1|_RX|104 0  1.937922998085e-12
L_PTL_P3_1|_RX|RB3 _PTL_P3_1|_RX|107 0  1.550338398468e-12
B_PTL_G3_1|_TX|1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|2 JJMIT AREA=2.5
B_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|5 JJMIT AREA=2.5
I_PTL_G3_1|_TX|B1 0 _PTL_G3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_1|_TX|B2 0 _PTL_G3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|3  1.684e-12
L_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|6  3.596e-12
L_PTL_G3_1|_TX|1 G3_1 _PTL_G3_1|_TX|1  2.063e-12
L_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|4  4.123e-12
L_PTL_G3_1|_TX|3 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|7  2.193e-12
R_PTL_G3_1|_TX|D _PTL_G3_1|_TX|7 _PTL_G3_1|A_PTL  1.36
L_PTL_G3_1|_TX|P1 _PTL_G3_1|_TX|2 0  5.254e-13
L_PTL_G3_1|_TX|P2 _PTL_G3_1|_TX|5 0  5.141e-13
R_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|101  2.7439617672
R_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|104  2.7439617672
L_PTL_G3_1|_TX|RB1 _PTL_G3_1|_TX|101 0  1.550338398468e-12
L_PTL_G3_1|_TX|RB2 _PTL_G3_1|_TX|104 0  1.550338398468e-12
B_PTL_G3_1|_RX|1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|5 JJMIT AREA=2.0
B_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|8 JJMIT AREA=2.5
I_PTL_G3_1|_RX|B1 0 _PTL_G3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|3  2.777e-12
I_PTL_G3_1|_RX|B2 0 _PTL_G3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|6  2.685e-12
I_PTL_G3_1|_RX|B3 0 _PTL_G3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|9  2.764e-12
L_PTL_G3_1|_RX|1 _PTL_G3_1|A_PTL _PTL_G3_1|_RX|1  1.346e-12
L_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|4  6.348e-12
L_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7  5.197e-12
L_PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7 G3_1_RX  2.058e-12
L_PTL_G3_1|_RX|P1 _PTL_G3_1|_RX|2 0  4.795e-13
L_PTL_G3_1|_RX|P2 _PTL_G3_1|_RX|5 0  5.431e-13
L_PTL_G3_1|_RX|P3 _PTL_G3_1|_RX|8 0  5.339e-13
R_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|101  4.225701121488
R_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|104  3.429952209
R_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|107  2.7439617672
L_PTL_G3_1|_RX|RB1 _PTL_G3_1|_RX|101 0  2.38752113364072e-12
L_PTL_G3_1|_RX|RB2 _PTL_G3_1|_RX|104 0  1.937922998085e-12
L_PTL_G3_1|_RX|RB3 _PTL_G3_1|_RX|107 0  1.550338398468e-12
B_PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_1|_TX|B1 0 _PTL_IP1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_1|_TX|B2 0 _PTL_IP1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|3  1.684e-12
L_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|6  3.596e-12
L_PTL_IP1_1|_TX|1 IP1_1_OUT _PTL_IP1_1|_TX|1  2.063e-12
L_PTL_IP1_1|_TX|2 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|4  4.123e-12
L_PTL_IP1_1|_TX|3 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|7  2.193e-12
R_PTL_IP1_1|_TX|D _PTL_IP1_1|_TX|7 _PTL_IP1_1|A_PTL  1.36
L_PTL_IP1_1|_TX|P1 _PTL_IP1_1|_TX|2 0  5.254e-13
L_PTL_IP1_1|_TX|P2 _PTL_IP1_1|_TX|5 0  5.141e-13
R_PTL_IP1_1|_TX|B1 _PTL_IP1_1|_TX|1 _PTL_IP1_1|_TX|101  2.7439617672
R_PTL_IP1_1|_TX|B2 _PTL_IP1_1|_TX|4 _PTL_IP1_1|_TX|104  2.7439617672
L_PTL_IP1_1|_TX|RB1 _PTL_IP1_1|_TX|101 0  1.550338398468e-12
L_PTL_IP1_1|_TX|RB2 _PTL_IP1_1|_TX|104 0  1.550338398468e-12
B_PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_1|_RX|B1 0 _PTL_IP1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|3  2.777e-12
I_PTL_IP1_1|_RX|B2 0 _PTL_IP1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|6  2.685e-12
I_PTL_IP1_1|_RX|B3 0 _PTL_IP1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|9  2.764e-12
L_PTL_IP1_1|_RX|1 _PTL_IP1_1|A_PTL _PTL_IP1_1|_RX|1  1.346e-12
L_PTL_IP1_1|_RX|2 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|4  6.348e-12
L_PTL_IP1_1|_RX|3 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7  5.197e-12
L_PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|7 IP1_1_OUT_RX  2.058e-12
L_PTL_IP1_1|_RX|P1 _PTL_IP1_1|_RX|2 0  4.795e-13
L_PTL_IP1_1|_RX|P2 _PTL_IP1_1|_RX|5 0  5.431e-13
L_PTL_IP1_1|_RX|P3 _PTL_IP1_1|_RX|8 0  5.339e-13
R_PTL_IP1_1|_RX|B1 _PTL_IP1_1|_RX|1 _PTL_IP1_1|_RX|101  4.225701121488
R_PTL_IP1_1|_RX|B2 _PTL_IP1_1|_RX|4 _PTL_IP1_1|_RX|104  3.429952209
R_PTL_IP1_1|_RX|B3 _PTL_IP1_1|_RX|7 _PTL_IP1_1|_RX|107  2.7439617672
L_PTL_IP1_1|_RX|RB1 _PTL_IP1_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_1|_RX|RB2 _PTL_IP1_1|_RX|104 0  1.937922998085e-12
L_PTL_IP1_1|_RX|RB3 _PTL_IP1_1|_RX|107 0  1.550338398468e-12
B_PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_1|_TX|B1 0 _PTL_IP2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_1|_TX|B2 0 _PTL_IP2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|3  1.684e-12
L_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|6  3.596e-12
L_PTL_IP2_1|_TX|1 IP2_1_OUT _PTL_IP2_1|_TX|1  2.063e-12
L_PTL_IP2_1|_TX|2 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|4  4.123e-12
L_PTL_IP2_1|_TX|3 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|7  2.193e-12
R_PTL_IP2_1|_TX|D _PTL_IP2_1|_TX|7 _PTL_IP2_1|A_PTL  1.36
L_PTL_IP2_1|_TX|P1 _PTL_IP2_1|_TX|2 0  5.254e-13
L_PTL_IP2_1|_TX|P2 _PTL_IP2_1|_TX|5 0  5.141e-13
R_PTL_IP2_1|_TX|B1 _PTL_IP2_1|_TX|1 _PTL_IP2_1|_TX|101  2.7439617672
R_PTL_IP2_1|_TX|B2 _PTL_IP2_1|_TX|4 _PTL_IP2_1|_TX|104  2.7439617672
L_PTL_IP2_1|_TX|RB1 _PTL_IP2_1|_TX|101 0  1.550338398468e-12
L_PTL_IP2_1|_TX|RB2 _PTL_IP2_1|_TX|104 0  1.550338398468e-12
B_PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_1|_RX|B1 0 _PTL_IP2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|3  2.777e-12
I_PTL_IP2_1|_RX|B2 0 _PTL_IP2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|6  2.685e-12
I_PTL_IP2_1|_RX|B3 0 _PTL_IP2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|9  2.764e-12
L_PTL_IP2_1|_RX|1 _PTL_IP2_1|A_PTL _PTL_IP2_1|_RX|1  1.346e-12
L_PTL_IP2_1|_RX|2 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|4  6.348e-12
L_PTL_IP2_1|_RX|3 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7  5.197e-12
L_PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|7 IP2_1_OUT_RX  2.058e-12
L_PTL_IP2_1|_RX|P1 _PTL_IP2_1|_RX|2 0  4.795e-13
L_PTL_IP2_1|_RX|P2 _PTL_IP2_1|_RX|5 0  5.431e-13
L_PTL_IP2_1|_RX|P3 _PTL_IP2_1|_RX|8 0  5.339e-13
R_PTL_IP2_1|_RX|B1 _PTL_IP2_1|_RX|1 _PTL_IP2_1|_RX|101  4.225701121488
R_PTL_IP2_1|_RX|B2 _PTL_IP2_1|_RX|4 _PTL_IP2_1|_RX|104  3.429952209
R_PTL_IP2_1|_RX|B3 _PTL_IP2_1|_RX|7 _PTL_IP2_1|_RX|107  2.7439617672
L_PTL_IP2_1|_RX|RB1 _PTL_IP2_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_1|_RX|RB2 _PTL_IP2_1|_RX|104 0  1.937922998085e-12
L_PTL_IP2_1|_RX|RB3 _PTL_IP2_1|_RX|107 0  1.550338398468e-12
B_PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_1|_TX|B1 0 _PTL_IP3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_1|_TX|B2 0 _PTL_IP3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|3  1.684e-12
L_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|6  3.596e-12
L_PTL_IP3_1|_TX|1 IP3_1_OUT _PTL_IP3_1|_TX|1  2.063e-12
L_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|4  4.123e-12
L_PTL_IP3_1|_TX|3 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|7  2.193e-12
R_PTL_IP3_1|_TX|D _PTL_IP3_1|_TX|7 _PTL_IP3_1|A_PTL  1.36
L_PTL_IP3_1|_TX|P1 _PTL_IP3_1|_TX|2 0  5.254e-13
L_PTL_IP3_1|_TX|P2 _PTL_IP3_1|_TX|5 0  5.141e-13
R_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|101  2.7439617672
R_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|104  2.7439617672
L_PTL_IP3_1|_TX|RB1 _PTL_IP3_1|_TX|101 0  1.550338398468e-12
L_PTL_IP3_1|_TX|RB2 _PTL_IP3_1|_TX|104 0  1.550338398468e-12
B_PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_1|_RX|B1 0 _PTL_IP3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|3  2.777e-12
I_PTL_IP3_1|_RX|B2 0 _PTL_IP3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|6  2.685e-12
I_PTL_IP3_1|_RX|B3 0 _PTL_IP3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|9  2.764e-12
L_PTL_IP3_1|_RX|1 _PTL_IP3_1|A_PTL _PTL_IP3_1|_RX|1  1.346e-12
L_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|4  6.348e-12
L_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7  5.197e-12
L_PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7 IP3_1_OUT_RX  2.058e-12
L_PTL_IP3_1|_RX|P1 _PTL_IP3_1|_RX|2 0  4.795e-13
L_PTL_IP3_1|_RX|P2 _PTL_IP3_1|_RX|5 0  5.431e-13
L_PTL_IP3_1|_RX|P3 _PTL_IP3_1|_RX|8 0  5.339e-13
R_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|101  4.225701121488
R_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|104  3.429952209
R_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|107  2.7439617672
L_PTL_IP3_1|_RX|RB1 _PTL_IP3_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_1|_RX|RB2 _PTL_IP3_1|_RX|104 0  1.937922998085e-12
L_PTL_IP3_1|_RX|RB3 _PTL_IP3_1|_RX|107 0  1.550338398468e-12
LSPL_G1_1|SPL1|1 G1_1_RX SPL_G1_1|SPL1|D1  2e-12
LSPL_G1_1|SPL1|2 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|D2  4.135667696e-12
LSPL_G1_1|SPL1|3 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|JCT  9.84682784761905e-13
LSPL_G1_1|SPL1|4 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QA1  9.84682784761905e-13
LSPL_G1_1|SPL1|5 SPL_G1_1|SPL1|QA1 G1_1_TO1  2e-12
LSPL_G1_1|SPL1|6 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QB1  9.84682784761905e-13
LSPL_G1_1|SPL1|7 SPL_G1_1|SPL1|QB1 SPL_G1_1|QTMP  2e-12
LSPL_G1_1|SPL2|1 SPL_G1_1|QTMP SPL_G1_1|SPL2|D1  2e-12
LSPL_G1_1|SPL2|2 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|D2  4.135667696e-12
LSPL_G1_1|SPL2|3 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|JCT  9.84682784761905e-13
LSPL_G1_1|SPL2|4 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QA1  9.84682784761905e-13
LSPL_G1_1|SPL2|5 SPL_G1_1|SPL2|QA1 G1_1_TO2  2e-12
LSPL_G1_1|SPL2|6 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QB1  9.84682784761905e-13
LSPL_G1_1|SPL2|7 SPL_G1_1|SPL2|QB1 G1_1_TO3  2e-12
L_PG0_12|P|1 P0_1_RX _PG0_12|P|A1  2.067833848e-12
L_PG0_12|P|2 _PG0_12|P|A1 _PG0_12|P|A2  4.135667696e-12
L_PG0_12|P|3 _PG0_12|P|A3 _PG0_12|P|A4  8.271335392e-12
L_PG0_12|P|T T08 _PG0_12|P|T1  2.067833848e-12
L_PG0_12|P|4 _PG0_12|P|T1 _PG0_12|P|T2  4.135667696e-12
L_PG0_12|P|5 _PG0_12|P|A4 _PG0_12|P|Q1  4.135667696e-12
L_PG0_12|P|6 _PG0_12|P|Q1 P0_2  2.067833848e-12
L_PG0_12|G|1 G0_1_RX _PG0_12|G|A1  2.067833848e-12
L_PG0_12|G|2 _PG0_12|G|A1 _PG0_12|G|A2  4.135667696e-12
L_PG0_12|G|3 _PG0_12|G|A3 _PG0_12|G|A4  8.271335392e-12
L_PG0_12|G|T T08 _PG0_12|G|T1  2.067833848e-12
L_PG0_12|G|4 _PG0_12|G|T1 _PG0_12|G|T2  4.135667696e-12
L_PG0_12|G|5 _PG0_12|G|A4 _PG0_12|G|Q1  4.135667696e-12
L_PG0_12|G|6 _PG0_12|G|Q1 G0_2  2.067833848e-12
L_PG1_12|I_1|B _PG1_12|A1 _PG1_12|I_1|MID  2e-12
I_PG1_12|I_1|B 0 _PG1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_3|B _PG1_12|A3 _PG1_12|I_3|MID  2e-12
I_PG1_12|I_3|B 0 _PG1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_12|I_T|B _PG1_12|T1 _PG1_12|I_T|MID  2e-12
I_PG1_12|I_T|B 0 _PG1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_6|B _PG1_12|Q1 _PG1_12|I_6|MID  2e-12
I_PG1_12|I_6|B 0 _PG1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_12|1|1 _PG1_12|A1 _PG1_12|1|MID_SERIES JJMIT AREA=2.5
L_PG1_12|1|P _PG1_12|1|MID_SERIES 0  2e-13
R_PG1_12|1|B _PG1_12|A1 _PG1_12|1|MID_SHUNT  2.7439617672
L_PG1_12|1|RB _PG1_12|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|23|1 _PG1_12|A2 _PG1_12|A3 JJMIT AREA=1.7857142857142858
R_PG1_12|23|B _PG1_12|A2 _PG1_12|23|MID_SHUNT  3.84154647408
L_PG1_12|23|RB _PG1_12|23|MID_SHUNT _PG1_12|A3  2.1704737578552e-12
B_PG1_12|3|1 _PG1_12|A3 _PG1_12|3|MID_SERIES JJMIT AREA=2.5
L_PG1_12|3|P _PG1_12|3|MID_SERIES 0  2e-13
R_PG1_12|3|B _PG1_12|A3 _PG1_12|3|MID_SHUNT  2.7439617672
L_PG1_12|3|RB _PG1_12|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|4|1 _PG1_12|A4 _PG1_12|4|MID_SERIES JJMIT AREA=2.5
L_PG1_12|4|P _PG1_12|4|MID_SERIES 0  2e-13
R_PG1_12|4|B _PG1_12|A4 _PG1_12|4|MID_SHUNT  2.7439617672
L_PG1_12|4|RB _PG1_12|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|T|1 _PG1_12|T1 _PG1_12|T|MID_SERIES JJMIT AREA=2.5
L_PG1_12|T|P _PG1_12|T|MID_SERIES 0  2e-13
R_PG1_12|T|B _PG1_12|T1 _PG1_12|T|MID_SHUNT  2.7439617672
L_PG1_12|T|RB _PG1_12|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|45|1 _PG1_12|T2 _PG1_12|A4 JJMIT AREA=1.7857142857142858
R_PG1_12|45|B _PG1_12|T2 _PG1_12|45|MID_SHUNT  3.84154647408
L_PG1_12|45|RB _PG1_12|45|MID_SHUNT _PG1_12|A4  2.1704737578552e-12
B_PG1_12|6|1 _PG1_12|Q1 _PG1_12|6|MID_SERIES JJMIT AREA=2.5
L_PG1_12|6|P _PG1_12|6|MID_SERIES 0  2e-13
R_PG1_12|6|B _PG1_12|Q1 _PG1_12|6|MID_SHUNT  2.7439617672
L_PG1_12|6|RB _PG1_12|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|1 G2_1_RX _PG2_12|_SPL_G1|D1  2e-12
L_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|D2  4.135667696e-12
L_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG2_12|_SPL_G1|5 _PG2_12|_SPL_G1|QA1 _PG2_12|G1_COPY_1  2e-12
L_PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|QB1 _PG2_12|G1_COPY_2  2e-12
L_PG2_12|_PG|A1 P2_1_RX _PG2_12|_PG|A1  2.067833848e-12
L_PG2_12|_PG|A2 _PG2_12|_PG|A1 _PG2_12|_PG|A2  4.135667696e-12
L_PG2_12|_PG|A3 _PG2_12|_PG|A3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|B1 _PG2_12|G1_COPY_1 _PG2_12|_PG|B1  2.067833848e-12
L_PG2_12|_PG|B2 _PG2_12|_PG|B1 _PG2_12|_PG|B2  4.135667696e-12
L_PG2_12|_PG|B3 _PG2_12|_PG|B3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|Q3 _PG2_12|_PG|Q3 _PG2_12|_PG|Q2  4.135667696e-12
L_PG2_12|_PG|Q2 _PG2_12|_PG|Q2 _PG2_12|_PG|Q1  4.135667696e-12
L_PG2_12|_PG|Q1 _PG2_12|_PG|Q1 _PG2_12|PG  2.067833848e-12
L_PG2_12|_GG|A1 G1_1_TO2 _PG2_12|_GG|A1  2.067833848e-12
L_PG2_12|_GG|A2 _PG2_12|_GG|A1 _PG2_12|_GG|A2  4.135667696e-12
L_PG2_12|_GG|A3 _PG2_12|_GG|A3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|B1 _PG2_12|G1_COPY_2 _PG2_12|_GG|B1  2.067833848e-12
L_PG2_12|_GG|B2 _PG2_12|_GG|B1 _PG2_12|_GG|B2  4.135667696e-12
L_PG2_12|_GG|B3 _PG2_12|_GG|B3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|Q3 _PG2_12|_GG|Q3 _PG2_12|_GG|Q2  4.135667696e-12
L_PG2_12|_GG|Q2 _PG2_12|_GG|Q2 _PG2_12|_GG|Q1  4.135667696e-12
L_PG2_12|_GG|Q1 _PG2_12|_GG|Q1 _PG2_12|GG  2.067833848e-12
L_PG2_12|_DFF_PG|1 _PG2_12|PG _PG2_12|_DFF_PG|A1  2.067833848e-12
L_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|A2  4.135667696e-12
L_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|A4  8.271335392e-12
L_PG2_12|_DFF_PG|T T10 _PG2_12|_DFF_PG|T1  2.067833848e-12
L_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T2  4.135667696e-12
L_PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|Q1  4.135667696e-12
L_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|Q1 _PG2_12|PG_SYNC  2.067833848e-12
L_PG2_12|_DFF_GG|1 _PG2_12|GG _PG2_12|_DFF_GG|A1  2.067833848e-12
L_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|A2  4.135667696e-12
L_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|A4  8.271335392e-12
L_PG2_12|_DFF_GG|T T10 _PG2_12|_DFF_GG|T1  2.067833848e-12
L_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T2  4.135667696e-12
L_PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|Q1  4.135667696e-12
L_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|Q1 _PG2_12|GG_SYNC  2.067833848e-12
L_PG2_12|_AND_G|A1 _PG2_12|PG_SYNC _PG2_12|_AND_G|A1  2.067833848e-12
L_PG2_12|_AND_G|A2 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A2  4.135667696e-12
L_PG2_12|_AND_G|A3 _PG2_12|_AND_G|A3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|B1 _PG2_12|GG_SYNC _PG2_12|_AND_G|B1  2.067833848e-12
L_PG2_12|_AND_G|B2 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B2  4.135667696e-12
L_PG2_12|_AND_G|B3 _PG2_12|_AND_G|B3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q2  4.135667696e-12
L_PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q1  4.135667696e-12
L_PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1 G2_2  2.067833848e-12
L_PG3_12|_SPL_G1|1 G3_1_RX _PG3_12|_SPL_G1|D1  2e-12
L_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|D2  4.135667696e-12
L_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_12|_SPL_G1|5 _PG3_12|_SPL_G1|QA1 _PG3_12|G1_COPY_1  2e-12
L_PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|QB1 _PG3_12|G1_COPY_2  2e-12
L_PG3_12|_PG|A1 P3_1_RX _PG3_12|_PG|A1  2.067833848e-12
L_PG3_12|_PG|A2 _PG3_12|_PG|A1 _PG3_12|_PG|A2  4.135667696e-12
L_PG3_12|_PG|A3 _PG3_12|_PG|A3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|B1 _PG3_12|G1_COPY_1 _PG3_12|_PG|B1  2.067833848e-12
L_PG3_12|_PG|B2 _PG3_12|_PG|B1 _PG3_12|_PG|B2  4.135667696e-12
L_PG3_12|_PG|B3 _PG3_12|_PG|B3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|Q3 _PG3_12|_PG|Q3 _PG3_12|_PG|Q2  4.135667696e-12
L_PG3_12|_PG|Q2 _PG3_12|_PG|Q2 _PG3_12|_PG|Q1  4.135667696e-12
L_PG3_12|_PG|Q1 _PG3_12|_PG|Q1 _PG3_12|PG  2.067833848e-12
L_PG3_12|_GG|A1 G1_1_TO3 _PG3_12|_GG|A1  2.067833848e-12
L_PG3_12|_GG|A2 _PG3_12|_GG|A1 _PG3_12|_GG|A2  4.135667696e-12
L_PG3_12|_GG|A3 _PG3_12|_GG|A3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|B1 _PG3_12|G1_COPY_2 _PG3_12|_GG|B1  2.067833848e-12
L_PG3_12|_GG|B2 _PG3_12|_GG|B1 _PG3_12|_GG|B2  4.135667696e-12
L_PG3_12|_GG|B3 _PG3_12|_GG|B3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|Q3 _PG3_12|_GG|Q3 _PG3_12|_GG|Q2  4.135667696e-12
L_PG3_12|_GG|Q2 _PG3_12|_GG|Q2 _PG3_12|_GG|Q1  4.135667696e-12
L_PG3_12|_GG|Q1 _PG3_12|_GG|Q1 _PG3_12|GG  2.067833848e-12
L_PG3_12|_DFF_PG|1 _PG3_12|PG _PG3_12|_DFF_PG|A1  2.067833848e-12
L_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|A2  4.135667696e-12
L_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|A4  8.271335392e-12
L_PG3_12|_DFF_PG|T T11 _PG3_12|_DFF_PG|T1  2.067833848e-12
L_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T2  4.135667696e-12
L_PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|Q1  4.135667696e-12
L_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|Q1 _PG3_12|PG_SYNC  2.067833848e-12
L_PG3_12|_DFF_GG|1 _PG3_12|GG _PG3_12|_DFF_GG|A1  2.067833848e-12
L_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|A2  4.135667696e-12
L_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|A4  8.271335392e-12
L_PG3_12|_DFF_GG|T T11 _PG3_12|_DFF_GG|T1  2.067833848e-12
L_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T2  4.135667696e-12
L_PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|Q1  4.135667696e-12
L_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|Q1 _PG3_12|GG_SYNC  2.067833848e-12
L_PG3_12|_AND_G|A1 _PG3_12|PG_SYNC _PG3_12|_AND_G|A1  2.067833848e-12
L_PG3_12|_AND_G|A2 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A2  4.135667696e-12
L_PG3_12|_AND_G|A3 _PG3_12|_AND_G|A3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|B1 _PG3_12|GG_SYNC _PG3_12|_AND_G|B1  2.067833848e-12
L_PG3_12|_AND_G|B2 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B2  4.135667696e-12
L_PG3_12|_AND_G|B3 _PG3_12|_AND_G|B3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q2  4.135667696e-12
L_PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q1  4.135667696e-12
L_PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1 G3_2  2.067833848e-12
L_DFF_IP1_12|I_1|B _DFF_IP1_12|A1 _DFF_IP1_12|I_1|MID  2e-12
I_DFF_IP1_12|I_1|B 0 _DFF_IP1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_3|B _DFF_IP1_12|A3 _DFF_IP1_12|I_3|MID  2e-12
I_DFF_IP1_12|I_3|B 0 _DFF_IP1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_12|I_T|B _DFF_IP1_12|T1 _DFF_IP1_12|I_T|MID  2e-12
I_DFF_IP1_12|I_T|B 0 _DFF_IP1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_6|B _DFF_IP1_12|Q1 _DFF_IP1_12|I_6|MID  2e-12
I_DFF_IP1_12|I_6|B 0 _DFF_IP1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_12|1|1 _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|1|P _DFF_IP1_12|1|MID_SERIES 0  2e-13
R_DFF_IP1_12|1|B _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SHUNT  2.7439617672
L_DFF_IP1_12|1|RB _DFF_IP1_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|23|1 _DFF_IP1_12|A2 _DFF_IP1_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|23|B _DFF_IP1_12|A2 _DFF_IP1_12|23|MID_SHUNT  3.84154647408
L_DFF_IP1_12|23|RB _DFF_IP1_12|23|MID_SHUNT _DFF_IP1_12|A3  2.1704737578552e-12
B_DFF_IP1_12|3|1 _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|3|P _DFF_IP1_12|3|MID_SERIES 0  2e-13
R_DFF_IP1_12|3|B _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SHUNT  2.7439617672
L_DFF_IP1_12|3|RB _DFF_IP1_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|4|1 _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|4|P _DFF_IP1_12|4|MID_SERIES 0  2e-13
R_DFF_IP1_12|4|B _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SHUNT  2.7439617672
L_DFF_IP1_12|4|RB _DFF_IP1_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|T|1 _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|T|P _DFF_IP1_12|T|MID_SERIES 0  2e-13
R_DFF_IP1_12|T|B _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SHUNT  2.7439617672
L_DFF_IP1_12|T|RB _DFF_IP1_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|45|1 _DFF_IP1_12|T2 _DFF_IP1_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|45|B _DFF_IP1_12|T2 _DFF_IP1_12|45|MID_SHUNT  3.84154647408
L_DFF_IP1_12|45|RB _DFF_IP1_12|45|MID_SHUNT _DFF_IP1_12|A4  2.1704737578552e-12
B_DFF_IP1_12|6|1 _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|6|P _DFF_IP1_12|6|MID_SERIES 0  2e-13
R_DFF_IP1_12|6|B _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SHUNT  2.7439617672
L_DFF_IP1_12|6|RB _DFF_IP1_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_12|I_1|B _DFF_IP2_12|A1 _DFF_IP2_12|I_1|MID  2e-12
I_DFF_IP2_12|I_1|B 0 _DFF_IP2_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_3|B _DFF_IP2_12|A3 _DFF_IP2_12|I_3|MID  2e-12
I_DFF_IP2_12|I_3|B 0 _DFF_IP2_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_12|I_T|B _DFF_IP2_12|T1 _DFF_IP2_12|I_T|MID  2e-12
I_DFF_IP2_12|I_T|B 0 _DFF_IP2_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_6|B _DFF_IP2_12|Q1 _DFF_IP2_12|I_6|MID  2e-12
I_DFF_IP2_12|I_6|B 0 _DFF_IP2_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_12|1|1 _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|1|P _DFF_IP2_12|1|MID_SERIES 0  2e-13
R_DFF_IP2_12|1|B _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SHUNT  2.7439617672
L_DFF_IP2_12|1|RB _DFF_IP2_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|23|1 _DFF_IP2_12|A2 _DFF_IP2_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|23|B _DFF_IP2_12|A2 _DFF_IP2_12|23|MID_SHUNT  3.84154647408
L_DFF_IP2_12|23|RB _DFF_IP2_12|23|MID_SHUNT _DFF_IP2_12|A3  2.1704737578552e-12
B_DFF_IP2_12|3|1 _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|3|P _DFF_IP2_12|3|MID_SERIES 0  2e-13
R_DFF_IP2_12|3|B _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SHUNT  2.7439617672
L_DFF_IP2_12|3|RB _DFF_IP2_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|4|1 _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|4|P _DFF_IP2_12|4|MID_SERIES 0  2e-13
R_DFF_IP2_12|4|B _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SHUNT  2.7439617672
L_DFF_IP2_12|4|RB _DFF_IP2_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|T|1 _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|T|P _DFF_IP2_12|T|MID_SERIES 0  2e-13
R_DFF_IP2_12|T|B _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SHUNT  2.7439617672
L_DFF_IP2_12|T|RB _DFF_IP2_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|45|1 _DFF_IP2_12|T2 _DFF_IP2_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|45|B _DFF_IP2_12|T2 _DFF_IP2_12|45|MID_SHUNT  3.84154647408
L_DFF_IP2_12|45|RB _DFF_IP2_12|45|MID_SHUNT _DFF_IP2_12|A4  2.1704737578552e-12
B_DFF_IP2_12|6|1 _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|6|P _DFF_IP2_12|6|MID_SERIES 0  2e-13
R_DFF_IP2_12|6|B _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SHUNT  2.7439617672
L_DFF_IP2_12|6|RB _DFF_IP2_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_12|I_1|B _DFF_IP3_12|A1 _DFF_IP3_12|I_1|MID  2e-12
I_DFF_IP3_12|I_1|B 0 _DFF_IP3_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_3|B _DFF_IP3_12|A3 _DFF_IP3_12|I_3|MID  2e-12
I_DFF_IP3_12|I_3|B 0 _DFF_IP3_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_12|I_T|B _DFF_IP3_12|T1 _DFF_IP3_12|I_T|MID  2e-12
I_DFF_IP3_12|I_T|B 0 _DFF_IP3_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_6|B _DFF_IP3_12|Q1 _DFF_IP3_12|I_6|MID  2e-12
I_DFF_IP3_12|I_6|B 0 _DFF_IP3_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_12|1|1 _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|1|P _DFF_IP3_12|1|MID_SERIES 0  2e-13
R_DFF_IP3_12|1|B _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SHUNT  2.7439617672
L_DFF_IP3_12|1|RB _DFF_IP3_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|23|1 _DFF_IP3_12|A2 _DFF_IP3_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|23|B _DFF_IP3_12|A2 _DFF_IP3_12|23|MID_SHUNT  3.84154647408
L_DFF_IP3_12|23|RB _DFF_IP3_12|23|MID_SHUNT _DFF_IP3_12|A3  2.1704737578552e-12
B_DFF_IP3_12|3|1 _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|3|P _DFF_IP3_12|3|MID_SERIES 0  2e-13
R_DFF_IP3_12|3|B _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SHUNT  2.7439617672
L_DFF_IP3_12|3|RB _DFF_IP3_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|4|1 _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|4|P _DFF_IP3_12|4|MID_SERIES 0  2e-13
R_DFF_IP3_12|4|B _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SHUNT  2.7439617672
L_DFF_IP3_12|4|RB _DFF_IP3_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|T|1 _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|T|P _DFF_IP3_12|T|MID_SERIES 0  2e-13
R_DFF_IP3_12|T|B _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SHUNT  2.7439617672
L_DFF_IP3_12|T|RB _DFF_IP3_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|45|1 _DFF_IP3_12|T2 _DFF_IP3_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|45|B _DFF_IP3_12|T2 _DFF_IP3_12|45|MID_SHUNT  3.84154647408
L_DFF_IP3_12|45|RB _DFF_IP3_12|45|MID_SHUNT _DFF_IP3_12|A4  2.1704737578552e-12
B_DFF_IP3_12|6|1 _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|6|P _DFF_IP3_12|6|MID_SERIES 0  2e-13
R_DFF_IP3_12|6|B _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SHUNT  2.7439617672
L_DFF_IP3_12|6|RB _DFF_IP3_12|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_P0_2|_TX|1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|2 JJMIT AREA=2.5
B_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|5 JJMIT AREA=2.5
I_PTL_P0_2|_TX|B1 0 _PTL_P0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P0_2|_TX|B2 0 _PTL_P0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|3  1.684e-12
L_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|6  3.596e-12
L_PTL_P0_2|_TX|1 P0_2 _PTL_P0_2|_TX|1  2.063e-12
L_PTL_P0_2|_TX|2 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|4  4.123e-12
L_PTL_P0_2|_TX|3 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|7  2.193e-12
R_PTL_P0_2|_TX|D _PTL_P0_2|_TX|7 _PTL_P0_2|A_PTL  1.36
L_PTL_P0_2|_TX|P1 _PTL_P0_2|_TX|2 0  5.254e-13
L_PTL_P0_2|_TX|P2 _PTL_P0_2|_TX|5 0  5.141e-13
R_PTL_P0_2|_TX|B1 _PTL_P0_2|_TX|1 _PTL_P0_2|_TX|101  2.7439617672
R_PTL_P0_2|_TX|B2 _PTL_P0_2|_TX|4 _PTL_P0_2|_TX|104  2.7439617672
L_PTL_P0_2|_TX|RB1 _PTL_P0_2|_TX|101 0  1.550338398468e-12
L_PTL_P0_2|_TX|RB2 _PTL_P0_2|_TX|104 0  1.550338398468e-12
B_PTL_P0_2|_RX|1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|5 JJMIT AREA=2.0
B_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|8 JJMIT AREA=2.5
I_PTL_P0_2|_RX|B1 0 _PTL_P0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|3  2.777e-12
I_PTL_P0_2|_RX|B2 0 _PTL_P0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|6  2.685e-12
I_PTL_P0_2|_RX|B3 0 _PTL_P0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|9  2.764e-12
L_PTL_P0_2|_RX|1 _PTL_P0_2|A_PTL _PTL_P0_2|_RX|1  1.346e-12
L_PTL_P0_2|_RX|2 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|4  6.348e-12
L_PTL_P0_2|_RX|3 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7  5.197e-12
L_PTL_P0_2|_RX|4 _PTL_P0_2|_RX|7 _PTL_P0_2|A_PTL_RX  2.058e-12
L_PTL_P0_2|_RX|P1 _PTL_P0_2|_RX|2 0  4.795e-13
L_PTL_P0_2|_RX|P2 _PTL_P0_2|_RX|5 0  5.431e-13
L_PTL_P0_2|_RX|P3 _PTL_P0_2|_RX|8 0  5.339e-13
R_PTL_P0_2|_RX|B1 _PTL_P0_2|_RX|1 _PTL_P0_2|_RX|101  4.225701121488
R_PTL_P0_2|_RX|B2 _PTL_P0_2|_RX|4 _PTL_P0_2|_RX|104  3.429952209
R_PTL_P0_2|_RX|B3 _PTL_P0_2|_RX|7 _PTL_P0_2|_RX|107  2.7439617672
L_PTL_P0_2|_RX|RB1 _PTL_P0_2|_RX|101 0  2.38752113364072e-12
L_PTL_P0_2|_RX|RB2 _PTL_P0_2|_RX|104 0  1.937922998085e-12
L_PTL_P0_2|_RX|RB3 _PTL_P0_2|_RX|107 0  1.550338398468e-12
B_PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|2 JJMIT AREA=2.5
B_PTL_P0_2|_JTL|2 _PTL_P0_2|_JTL|6 _PTL_P0_2|_JTL|7 JJMIT AREA=2.5
I_PTL_P0_2|_JTL|B1 0 _PTL_P0_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_P0_2|_JTL|1 _PTL_P0_2|A_PTL_RX _PTL_P0_2|_JTL|1  2.067833848e-12
L_PTL_P0_2|_JTL|2 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|4  2.067833848e-12
L_PTL_P0_2|_JTL|3 _PTL_P0_2|_JTL|4 _PTL_P0_2|_JTL|6  2.067833848e-12
L_PTL_P0_2|_JTL|4 _PTL_P0_2|_JTL|6 P0_2_RX  2.067833848e-12
L_PTL_P0_2|_JTL|P1 _PTL_P0_2|_JTL|2 0  2e-13
L_PTL_P0_2|_JTL|P2 _PTL_P0_2|_JTL|7 0  2e-13
L_PTL_P0_2|_JTL|B1 _PTL_P0_2|_JTL|5 _PTL_P0_2|_JTL|4  2e-12
R_PTL_P0_2|_JTL|B1 _PTL_P0_2|_JTL|1 _PTL_P0_2|_JTL|3  2.7439617672
R_PTL_P0_2|_JTL|B2 _PTL_P0_2|_JTL|6 _PTL_P0_2|_JTL|8  2.7439617672
L_PTL_P0_2|_JTL|RB1 _PTL_P0_2|_JTL|3 0  1.750338398468e-12
L_PTL_P0_2|_JTL|RB2 _PTL_P0_2|_JTL|8 0  1.750338398468e-12
B_PTL_G0_2|_TX|1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|2 JJMIT AREA=2.5
B_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|5 JJMIT AREA=2.5
I_PTL_G0_2|_TX|B1 0 _PTL_G0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G0_2|_TX|B2 0 _PTL_G0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|3  1.684e-12
L_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|6  3.596e-12
L_PTL_G0_2|_TX|1 G0_2 _PTL_G0_2|_TX|1  2.063e-12
L_PTL_G0_2|_TX|2 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|4  4.123e-12
L_PTL_G0_2|_TX|3 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|7  2.193e-12
R_PTL_G0_2|_TX|D _PTL_G0_2|_TX|7 _PTL_G0_2|A_PTL  1.36
L_PTL_G0_2|_TX|P1 _PTL_G0_2|_TX|2 0  5.254e-13
L_PTL_G0_2|_TX|P2 _PTL_G0_2|_TX|5 0  5.141e-13
R_PTL_G0_2|_TX|B1 _PTL_G0_2|_TX|1 _PTL_G0_2|_TX|101  2.7439617672
R_PTL_G0_2|_TX|B2 _PTL_G0_2|_TX|4 _PTL_G0_2|_TX|104  2.7439617672
L_PTL_G0_2|_TX|RB1 _PTL_G0_2|_TX|101 0  1.550338398468e-12
L_PTL_G0_2|_TX|RB2 _PTL_G0_2|_TX|104 0  1.550338398468e-12
B_PTL_G0_2|_RX|1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|5 JJMIT AREA=2.0
B_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|8 JJMIT AREA=2.5
I_PTL_G0_2|_RX|B1 0 _PTL_G0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|3  2.777e-12
I_PTL_G0_2|_RX|B2 0 _PTL_G0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|6  2.685e-12
I_PTL_G0_2|_RX|B3 0 _PTL_G0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|9  2.764e-12
L_PTL_G0_2|_RX|1 _PTL_G0_2|A_PTL _PTL_G0_2|_RX|1  1.346e-12
L_PTL_G0_2|_RX|2 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|4  6.348e-12
L_PTL_G0_2|_RX|3 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7  5.197e-12
L_PTL_G0_2|_RX|4 _PTL_G0_2|_RX|7 _PTL_G0_2|A_PTL_RX  2.058e-12
L_PTL_G0_2|_RX|P1 _PTL_G0_2|_RX|2 0  4.795e-13
L_PTL_G0_2|_RX|P2 _PTL_G0_2|_RX|5 0  5.431e-13
L_PTL_G0_2|_RX|P3 _PTL_G0_2|_RX|8 0  5.339e-13
R_PTL_G0_2|_RX|B1 _PTL_G0_2|_RX|1 _PTL_G0_2|_RX|101  4.225701121488
R_PTL_G0_2|_RX|B2 _PTL_G0_2|_RX|4 _PTL_G0_2|_RX|104  3.429952209
R_PTL_G0_2|_RX|B3 _PTL_G0_2|_RX|7 _PTL_G0_2|_RX|107  2.7439617672
L_PTL_G0_2|_RX|RB1 _PTL_G0_2|_RX|101 0  2.38752113364072e-12
L_PTL_G0_2|_RX|RB2 _PTL_G0_2|_RX|104 0  1.937922998085e-12
L_PTL_G0_2|_RX|RB3 _PTL_G0_2|_RX|107 0  1.550338398468e-12
B_PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G0_2|_JTL|2 _PTL_G0_2|_JTL|6 _PTL_G0_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G0_2|_JTL|B1 0 _PTL_G0_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G0_2|_JTL|1 _PTL_G0_2|A_PTL_RX _PTL_G0_2|_JTL|1  2.067833848e-12
L_PTL_G0_2|_JTL|2 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|4  2.067833848e-12
L_PTL_G0_2|_JTL|3 _PTL_G0_2|_JTL|4 _PTL_G0_2|_JTL|6  2.067833848e-12
L_PTL_G0_2|_JTL|4 _PTL_G0_2|_JTL|6 G0_2_RX  2.067833848e-12
L_PTL_G0_2|_JTL|P1 _PTL_G0_2|_JTL|2 0  2e-13
L_PTL_G0_2|_JTL|P2 _PTL_G0_2|_JTL|7 0  2e-13
L_PTL_G0_2|_JTL|B1 _PTL_G0_2|_JTL|5 _PTL_G0_2|_JTL|4  2e-12
R_PTL_G0_2|_JTL|B1 _PTL_G0_2|_JTL|1 _PTL_G0_2|_JTL|3  2.7439617672
R_PTL_G0_2|_JTL|B2 _PTL_G0_2|_JTL|6 _PTL_G0_2|_JTL|8  2.7439617672
L_PTL_G0_2|_JTL|RB1 _PTL_G0_2|_JTL|3 0  1.750338398468e-12
L_PTL_G0_2|_JTL|RB2 _PTL_G0_2|_JTL|8 0  1.750338398468e-12
B_PTL_G1_2|_TX|1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|2 JJMIT AREA=2.5
B_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|5 JJMIT AREA=2.5
I_PTL_G1_2|_TX|B1 0 _PTL_G1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_2|_TX|B2 0 _PTL_G1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|3  1.684e-12
L_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|6  3.596e-12
L_PTL_G1_2|_TX|1 G1_2 _PTL_G1_2|_TX|1  2.063e-12
L_PTL_G1_2|_TX|2 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|4  4.123e-12
L_PTL_G1_2|_TX|3 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|7  2.193e-12
R_PTL_G1_2|_TX|D _PTL_G1_2|_TX|7 _PTL_G1_2|A_PTL  1.36
L_PTL_G1_2|_TX|P1 _PTL_G1_2|_TX|2 0  5.254e-13
L_PTL_G1_2|_TX|P2 _PTL_G1_2|_TX|5 0  5.141e-13
R_PTL_G1_2|_TX|B1 _PTL_G1_2|_TX|1 _PTL_G1_2|_TX|101  2.7439617672
R_PTL_G1_2|_TX|B2 _PTL_G1_2|_TX|4 _PTL_G1_2|_TX|104  2.7439617672
L_PTL_G1_2|_TX|RB1 _PTL_G1_2|_TX|101 0  1.550338398468e-12
L_PTL_G1_2|_TX|RB2 _PTL_G1_2|_TX|104 0  1.550338398468e-12
B_PTL_G1_2|_RX|1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|5 JJMIT AREA=2.0
B_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|8 JJMIT AREA=2.5
I_PTL_G1_2|_RX|B1 0 _PTL_G1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|3  2.777e-12
I_PTL_G1_2|_RX|B2 0 _PTL_G1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|6  2.685e-12
I_PTL_G1_2|_RX|B3 0 _PTL_G1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|9  2.764e-12
L_PTL_G1_2|_RX|1 _PTL_G1_2|A_PTL _PTL_G1_2|_RX|1  1.346e-12
L_PTL_G1_2|_RX|2 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|4  6.348e-12
L_PTL_G1_2|_RX|3 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7  5.197e-12
L_PTL_G1_2|_RX|4 _PTL_G1_2|_RX|7 _PTL_G1_2|A_PTL_RX  2.058e-12
L_PTL_G1_2|_RX|P1 _PTL_G1_2|_RX|2 0  4.795e-13
L_PTL_G1_2|_RX|P2 _PTL_G1_2|_RX|5 0  5.431e-13
L_PTL_G1_2|_RX|P3 _PTL_G1_2|_RX|8 0  5.339e-13
R_PTL_G1_2|_RX|B1 _PTL_G1_2|_RX|1 _PTL_G1_2|_RX|101  4.225701121488
R_PTL_G1_2|_RX|B2 _PTL_G1_2|_RX|4 _PTL_G1_2|_RX|104  3.429952209
R_PTL_G1_2|_RX|B3 _PTL_G1_2|_RX|7 _PTL_G1_2|_RX|107  2.7439617672
L_PTL_G1_2|_RX|RB1 _PTL_G1_2|_RX|101 0  2.38752113364072e-12
L_PTL_G1_2|_RX|RB2 _PTL_G1_2|_RX|104 0  1.937922998085e-12
L_PTL_G1_2|_RX|RB3 _PTL_G1_2|_RX|107 0  1.550338398468e-12
B_PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G1_2|_JTL|2 _PTL_G1_2|_JTL|6 _PTL_G1_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G1_2|_JTL|B1 0 _PTL_G1_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G1_2|_JTL|1 _PTL_G1_2|A_PTL_RX _PTL_G1_2|_JTL|1  2.067833848e-12
L_PTL_G1_2|_JTL|2 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|4  2.067833848e-12
L_PTL_G1_2|_JTL|3 _PTL_G1_2|_JTL|4 _PTL_G1_2|_JTL|6  2.067833848e-12
L_PTL_G1_2|_JTL|4 _PTL_G1_2|_JTL|6 G1_2_RX  2.067833848e-12
L_PTL_G1_2|_JTL|P1 _PTL_G1_2|_JTL|2 0  2e-13
L_PTL_G1_2|_JTL|P2 _PTL_G1_2|_JTL|7 0  2e-13
L_PTL_G1_2|_JTL|B1 _PTL_G1_2|_JTL|5 _PTL_G1_2|_JTL|4  2e-12
R_PTL_G1_2|_JTL|B1 _PTL_G1_2|_JTL|1 _PTL_G1_2|_JTL|3  2.7439617672
R_PTL_G1_2|_JTL|B2 _PTL_G1_2|_JTL|6 _PTL_G1_2|_JTL|8  2.7439617672
L_PTL_G1_2|_JTL|RB1 _PTL_G1_2|_JTL|3 0  1.750338398468e-12
L_PTL_G1_2|_JTL|RB2 _PTL_G1_2|_JTL|8 0  1.750338398468e-12
B_PTL_G2_2|_TX|1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|2 JJMIT AREA=2.5
B_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|5 JJMIT AREA=2.5
I_PTL_G2_2|_TX|B1 0 _PTL_G2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_2|_TX|B2 0 _PTL_G2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|3  1.684e-12
L_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|6  3.596e-12
L_PTL_G2_2|_TX|1 G2_2 _PTL_G2_2|_TX|1  2.063e-12
L_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|4  4.123e-12
L_PTL_G2_2|_TX|3 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|7  2.193e-12
R_PTL_G2_2|_TX|D _PTL_G2_2|_TX|7 _PTL_G2_2|A_PTL  1.36
L_PTL_G2_2|_TX|P1 _PTL_G2_2|_TX|2 0  5.254e-13
L_PTL_G2_2|_TX|P2 _PTL_G2_2|_TX|5 0  5.141e-13
R_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|101  2.7439617672
R_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|104  2.7439617672
L_PTL_G2_2|_TX|RB1 _PTL_G2_2|_TX|101 0  1.550338398468e-12
L_PTL_G2_2|_TX|RB2 _PTL_G2_2|_TX|104 0  1.550338398468e-12
B_PTL_G2_2|_RX|1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|5 JJMIT AREA=2.0
B_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|8 JJMIT AREA=2.5
I_PTL_G2_2|_RX|B1 0 _PTL_G2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|3  2.777e-12
I_PTL_G2_2|_RX|B2 0 _PTL_G2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|6  2.685e-12
I_PTL_G2_2|_RX|B3 0 _PTL_G2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|9  2.764e-12
L_PTL_G2_2|_RX|1 _PTL_G2_2|A_PTL _PTL_G2_2|_RX|1  1.346e-12
L_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|4  6.348e-12
L_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7  5.197e-12
L_PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7 _PTL_G2_2|A_PTL_RX  2.058e-12
L_PTL_G2_2|_RX|P1 _PTL_G2_2|_RX|2 0  4.795e-13
L_PTL_G2_2|_RX|P2 _PTL_G2_2|_RX|5 0  5.431e-13
L_PTL_G2_2|_RX|P3 _PTL_G2_2|_RX|8 0  5.339e-13
R_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|101  4.225701121488
R_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|104  3.429952209
R_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|107  2.7439617672
L_PTL_G2_2|_RX|RB1 _PTL_G2_2|_RX|101 0  2.38752113364072e-12
L_PTL_G2_2|_RX|RB2 _PTL_G2_2|_RX|104 0  1.937922998085e-12
L_PTL_G2_2|_RX|RB3 _PTL_G2_2|_RX|107 0  1.550338398468e-12
B_PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G2_2|_JTL|2 _PTL_G2_2|_JTL|6 _PTL_G2_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G2_2|_JTL|B1 0 _PTL_G2_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G2_2|_JTL|1 _PTL_G2_2|A_PTL_RX _PTL_G2_2|_JTL|1  2.067833848e-12
L_PTL_G2_2|_JTL|2 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|4  2.067833848e-12
L_PTL_G2_2|_JTL|3 _PTL_G2_2|_JTL|4 _PTL_G2_2|_JTL|6  2.067833848e-12
L_PTL_G2_2|_JTL|4 _PTL_G2_2|_JTL|6 G2_2_RX  2.067833848e-12
L_PTL_G2_2|_JTL|P1 _PTL_G2_2|_JTL|2 0  2e-13
L_PTL_G2_2|_JTL|P2 _PTL_G2_2|_JTL|7 0  2e-13
L_PTL_G2_2|_JTL|B1 _PTL_G2_2|_JTL|5 _PTL_G2_2|_JTL|4  2e-12
R_PTL_G2_2|_JTL|B1 _PTL_G2_2|_JTL|1 _PTL_G2_2|_JTL|3  2.7439617672
R_PTL_G2_2|_JTL|B2 _PTL_G2_2|_JTL|6 _PTL_G2_2|_JTL|8  2.7439617672
L_PTL_G2_2|_JTL|RB1 _PTL_G2_2|_JTL|3 0  1.750338398468e-12
L_PTL_G2_2|_JTL|RB2 _PTL_G2_2|_JTL|8 0  1.750338398468e-12
B_PTL_G3_2|_TX|1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|2 JJMIT AREA=2.5
B_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|5 JJMIT AREA=2.5
I_PTL_G3_2|_TX|B1 0 _PTL_G3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_2|_TX|B2 0 _PTL_G3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|3  1.684e-12
L_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|6  3.596e-12
L_PTL_G3_2|_TX|1 G3_2 _PTL_G3_2|_TX|1  2.063e-12
L_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|4  4.123e-12
L_PTL_G3_2|_TX|3 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|7  2.193e-12
R_PTL_G3_2|_TX|D _PTL_G3_2|_TX|7 _PTL_G3_2|A_PTL  1.36
L_PTL_G3_2|_TX|P1 _PTL_G3_2|_TX|2 0  5.254e-13
L_PTL_G3_2|_TX|P2 _PTL_G3_2|_TX|5 0  5.141e-13
R_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|101  2.7439617672
R_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|104  2.7439617672
L_PTL_G3_2|_TX|RB1 _PTL_G3_2|_TX|101 0  1.550338398468e-12
L_PTL_G3_2|_TX|RB2 _PTL_G3_2|_TX|104 0  1.550338398468e-12
B_PTL_G3_2|_RX|1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|5 JJMIT AREA=2.0
B_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|8 JJMIT AREA=2.5
I_PTL_G3_2|_RX|B1 0 _PTL_G3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|3  2.777e-12
I_PTL_G3_2|_RX|B2 0 _PTL_G3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|6  2.685e-12
I_PTL_G3_2|_RX|B3 0 _PTL_G3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|9  2.764e-12
L_PTL_G3_2|_RX|1 _PTL_G3_2|A_PTL _PTL_G3_2|_RX|1  1.346e-12
L_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|4  6.348e-12
L_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7  5.197e-12
L_PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7 _PTL_G3_2|A_PTL_RX  2.058e-12
L_PTL_G3_2|_RX|P1 _PTL_G3_2|_RX|2 0  4.795e-13
L_PTL_G3_2|_RX|P2 _PTL_G3_2|_RX|5 0  5.431e-13
L_PTL_G3_2|_RX|P3 _PTL_G3_2|_RX|8 0  5.339e-13
R_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|101  4.225701121488
R_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|104  3.429952209
R_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|107  2.7439617672
L_PTL_G3_2|_RX|RB1 _PTL_G3_2|_RX|101 0  2.38752113364072e-12
L_PTL_G3_2|_RX|RB2 _PTL_G3_2|_RX|104 0  1.937922998085e-12
L_PTL_G3_2|_RX|RB3 _PTL_G3_2|_RX|107 0  1.550338398468e-12
B_PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|2 JJMIT AREA=2.5
B_PTL_G3_2|_JTL|2 _PTL_G3_2|_JTL|6 _PTL_G3_2|_JTL|7 JJMIT AREA=2.5
I_PTL_G3_2|_JTL|B1 0 _PTL_G3_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_G3_2|_JTL|1 _PTL_G3_2|A_PTL_RX _PTL_G3_2|_JTL|1  2.067833848e-12
L_PTL_G3_2|_JTL|2 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|4  2.067833848e-12
L_PTL_G3_2|_JTL|3 _PTL_G3_2|_JTL|4 _PTL_G3_2|_JTL|6  2.067833848e-12
L_PTL_G3_2|_JTL|4 _PTL_G3_2|_JTL|6 G3_2_RX  2.067833848e-12
L_PTL_G3_2|_JTL|P1 _PTL_G3_2|_JTL|2 0  2e-13
L_PTL_G3_2|_JTL|P2 _PTL_G3_2|_JTL|7 0  2e-13
L_PTL_G3_2|_JTL|B1 _PTL_G3_2|_JTL|5 _PTL_G3_2|_JTL|4  2e-12
R_PTL_G3_2|_JTL|B1 _PTL_G3_2|_JTL|1 _PTL_G3_2|_JTL|3  2.7439617672
R_PTL_G3_2|_JTL|B2 _PTL_G3_2|_JTL|6 _PTL_G3_2|_JTL|8  2.7439617672
L_PTL_G3_2|_JTL|RB1 _PTL_G3_2|_JTL|3 0  1.750338398468e-12
L_PTL_G3_2|_JTL|RB2 _PTL_G3_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_2|_TX|B1 0 _PTL_IP1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_2|_TX|B2 0 _PTL_IP1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|3  1.684e-12
L_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|6  3.596e-12
L_PTL_IP1_2|_TX|1 IP1_2_OUT _PTL_IP1_2|_TX|1  2.063e-12
L_PTL_IP1_2|_TX|2 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|4  4.123e-12
L_PTL_IP1_2|_TX|3 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|7  2.193e-12
R_PTL_IP1_2|_TX|D _PTL_IP1_2|_TX|7 _PTL_IP1_2|A_PTL  1.36
L_PTL_IP1_2|_TX|P1 _PTL_IP1_2|_TX|2 0  5.254e-13
L_PTL_IP1_2|_TX|P2 _PTL_IP1_2|_TX|5 0  5.141e-13
R_PTL_IP1_2|_TX|B1 _PTL_IP1_2|_TX|1 _PTL_IP1_2|_TX|101  2.7439617672
R_PTL_IP1_2|_TX|B2 _PTL_IP1_2|_TX|4 _PTL_IP1_2|_TX|104  2.7439617672
L_PTL_IP1_2|_TX|RB1 _PTL_IP1_2|_TX|101 0  1.550338398468e-12
L_PTL_IP1_2|_TX|RB2 _PTL_IP1_2|_TX|104 0  1.550338398468e-12
B_PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_2|_RX|B1 0 _PTL_IP1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|3  2.777e-12
I_PTL_IP1_2|_RX|B2 0 _PTL_IP1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|6  2.685e-12
I_PTL_IP1_2|_RX|B3 0 _PTL_IP1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|9  2.764e-12
L_PTL_IP1_2|_RX|1 _PTL_IP1_2|A_PTL _PTL_IP1_2|_RX|1  1.346e-12
L_PTL_IP1_2|_RX|2 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|4  6.348e-12
L_PTL_IP1_2|_RX|3 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7  5.197e-12
L_PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|7 _PTL_IP1_2|A_PTL_RX  2.058e-12
L_PTL_IP1_2|_RX|P1 _PTL_IP1_2|_RX|2 0  4.795e-13
L_PTL_IP1_2|_RX|P2 _PTL_IP1_2|_RX|5 0  5.431e-13
L_PTL_IP1_2|_RX|P3 _PTL_IP1_2|_RX|8 0  5.339e-13
R_PTL_IP1_2|_RX|B1 _PTL_IP1_2|_RX|1 _PTL_IP1_2|_RX|101  4.225701121488
R_PTL_IP1_2|_RX|B2 _PTL_IP1_2|_RX|4 _PTL_IP1_2|_RX|104  3.429952209
R_PTL_IP1_2|_RX|B3 _PTL_IP1_2|_RX|7 _PTL_IP1_2|_RX|107  2.7439617672
L_PTL_IP1_2|_RX|RB1 _PTL_IP1_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_2|_RX|RB2 _PTL_IP1_2|_RX|104 0  1.937922998085e-12
L_PTL_IP1_2|_RX|RB3 _PTL_IP1_2|_RX|107 0  1.550338398468e-12
B_PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP1_2|_JTL|2 _PTL_IP1_2|_JTL|6 _PTL_IP1_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP1_2|_JTL|B1 0 _PTL_IP1_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP1_2|_JTL|1 _PTL_IP1_2|A_PTL_RX _PTL_IP1_2|_JTL|1  2.067833848e-12
L_PTL_IP1_2|_JTL|2 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|4  2.067833848e-12
L_PTL_IP1_2|_JTL|3 _PTL_IP1_2|_JTL|4 _PTL_IP1_2|_JTL|6  2.067833848e-12
L_PTL_IP1_2|_JTL|4 _PTL_IP1_2|_JTL|6 IP1_2_OUT_RX  2.067833848e-12
L_PTL_IP1_2|_JTL|P1 _PTL_IP1_2|_JTL|2 0  2e-13
L_PTL_IP1_2|_JTL|P2 _PTL_IP1_2|_JTL|7 0  2e-13
L_PTL_IP1_2|_JTL|B1 _PTL_IP1_2|_JTL|5 _PTL_IP1_2|_JTL|4  2e-12
R_PTL_IP1_2|_JTL|B1 _PTL_IP1_2|_JTL|1 _PTL_IP1_2|_JTL|3  2.7439617672
R_PTL_IP1_2|_JTL|B2 _PTL_IP1_2|_JTL|6 _PTL_IP1_2|_JTL|8  2.7439617672
L_PTL_IP1_2|_JTL|RB1 _PTL_IP1_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP1_2|_JTL|RB2 _PTL_IP1_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_2|_TX|B1 0 _PTL_IP2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_2|_TX|B2 0 _PTL_IP2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|3  1.684e-12
L_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|6  3.596e-12
L_PTL_IP2_2|_TX|1 IP2_2_OUT _PTL_IP2_2|_TX|1  2.063e-12
L_PTL_IP2_2|_TX|2 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|4  4.123e-12
L_PTL_IP2_2|_TX|3 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|7  2.193e-12
R_PTL_IP2_2|_TX|D _PTL_IP2_2|_TX|7 _PTL_IP2_2|A_PTL  1.36
L_PTL_IP2_2|_TX|P1 _PTL_IP2_2|_TX|2 0  5.254e-13
L_PTL_IP2_2|_TX|P2 _PTL_IP2_2|_TX|5 0  5.141e-13
R_PTL_IP2_2|_TX|B1 _PTL_IP2_2|_TX|1 _PTL_IP2_2|_TX|101  2.7439617672
R_PTL_IP2_2|_TX|B2 _PTL_IP2_2|_TX|4 _PTL_IP2_2|_TX|104  2.7439617672
L_PTL_IP2_2|_TX|RB1 _PTL_IP2_2|_TX|101 0  1.550338398468e-12
L_PTL_IP2_2|_TX|RB2 _PTL_IP2_2|_TX|104 0  1.550338398468e-12
B_PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_2|_RX|B1 0 _PTL_IP2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|3  2.777e-12
I_PTL_IP2_2|_RX|B2 0 _PTL_IP2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|6  2.685e-12
I_PTL_IP2_2|_RX|B3 0 _PTL_IP2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|9  2.764e-12
L_PTL_IP2_2|_RX|1 _PTL_IP2_2|A_PTL _PTL_IP2_2|_RX|1  1.346e-12
L_PTL_IP2_2|_RX|2 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|4  6.348e-12
L_PTL_IP2_2|_RX|3 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7  5.197e-12
L_PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|7 _PTL_IP2_2|A_PTL_RX  2.058e-12
L_PTL_IP2_2|_RX|P1 _PTL_IP2_2|_RX|2 0  4.795e-13
L_PTL_IP2_2|_RX|P2 _PTL_IP2_2|_RX|5 0  5.431e-13
L_PTL_IP2_2|_RX|P3 _PTL_IP2_2|_RX|8 0  5.339e-13
R_PTL_IP2_2|_RX|B1 _PTL_IP2_2|_RX|1 _PTL_IP2_2|_RX|101  4.225701121488
R_PTL_IP2_2|_RX|B2 _PTL_IP2_2|_RX|4 _PTL_IP2_2|_RX|104  3.429952209
R_PTL_IP2_2|_RX|B3 _PTL_IP2_2|_RX|7 _PTL_IP2_2|_RX|107  2.7439617672
L_PTL_IP2_2|_RX|RB1 _PTL_IP2_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_2|_RX|RB2 _PTL_IP2_2|_RX|104 0  1.937922998085e-12
L_PTL_IP2_2|_RX|RB3 _PTL_IP2_2|_RX|107 0  1.550338398468e-12
B_PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP2_2|_JTL|2 _PTL_IP2_2|_JTL|6 _PTL_IP2_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP2_2|_JTL|B1 0 _PTL_IP2_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP2_2|_JTL|1 _PTL_IP2_2|A_PTL_RX _PTL_IP2_2|_JTL|1  2.067833848e-12
L_PTL_IP2_2|_JTL|2 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|4  2.067833848e-12
L_PTL_IP2_2|_JTL|3 _PTL_IP2_2|_JTL|4 _PTL_IP2_2|_JTL|6  2.067833848e-12
L_PTL_IP2_2|_JTL|4 _PTL_IP2_2|_JTL|6 IP2_2_OUT_RX  2.067833848e-12
L_PTL_IP2_2|_JTL|P1 _PTL_IP2_2|_JTL|2 0  2e-13
L_PTL_IP2_2|_JTL|P2 _PTL_IP2_2|_JTL|7 0  2e-13
L_PTL_IP2_2|_JTL|B1 _PTL_IP2_2|_JTL|5 _PTL_IP2_2|_JTL|4  2e-12
R_PTL_IP2_2|_JTL|B1 _PTL_IP2_2|_JTL|1 _PTL_IP2_2|_JTL|3  2.7439617672
R_PTL_IP2_2|_JTL|B2 _PTL_IP2_2|_JTL|6 _PTL_IP2_2|_JTL|8  2.7439617672
L_PTL_IP2_2|_JTL|RB1 _PTL_IP2_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP2_2|_JTL|RB2 _PTL_IP2_2|_JTL|8 0  1.750338398468e-12
B_PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_2|_TX|B1 0 _PTL_IP3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_2|_TX|B2 0 _PTL_IP3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|3  1.684e-12
L_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|6  3.596e-12
L_PTL_IP3_2|_TX|1 IP3_2_OUT _PTL_IP3_2|_TX|1  2.063e-12
L_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|4  4.123e-12
L_PTL_IP3_2|_TX|3 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|7  2.193e-12
R_PTL_IP3_2|_TX|D _PTL_IP3_2|_TX|7 _PTL_IP3_2|A_PTL  1.36
L_PTL_IP3_2|_TX|P1 _PTL_IP3_2|_TX|2 0  5.254e-13
L_PTL_IP3_2|_TX|P2 _PTL_IP3_2|_TX|5 0  5.141e-13
R_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|101  2.7439617672
R_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|104  2.7439617672
L_PTL_IP3_2|_TX|RB1 _PTL_IP3_2|_TX|101 0  1.550338398468e-12
L_PTL_IP3_2|_TX|RB2 _PTL_IP3_2|_TX|104 0  1.550338398468e-12
B_PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_2|_RX|B1 0 _PTL_IP3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|3  2.777e-12
I_PTL_IP3_2|_RX|B2 0 _PTL_IP3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|6  2.685e-12
I_PTL_IP3_2|_RX|B3 0 _PTL_IP3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|9  2.764e-12
L_PTL_IP3_2|_RX|1 _PTL_IP3_2|A_PTL _PTL_IP3_2|_RX|1  1.346e-12
L_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|4  6.348e-12
L_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7  5.197e-12
L_PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7 _PTL_IP3_2|A_PTL_RX  2.058e-12
L_PTL_IP3_2|_RX|P1 _PTL_IP3_2|_RX|2 0  4.795e-13
L_PTL_IP3_2|_RX|P2 _PTL_IP3_2|_RX|5 0  5.431e-13
L_PTL_IP3_2|_RX|P3 _PTL_IP3_2|_RX|8 0  5.339e-13
R_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|101  4.225701121488
R_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|104  3.429952209
R_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|107  2.7439617672
L_PTL_IP3_2|_RX|RB1 _PTL_IP3_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_2|_RX|RB2 _PTL_IP3_2|_RX|104 0  1.937922998085e-12
L_PTL_IP3_2|_RX|RB3 _PTL_IP3_2|_RX|107 0  1.550338398468e-12
B_PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|2 JJMIT AREA=2.5
B_PTL_IP3_2|_JTL|2 _PTL_IP3_2|_JTL|6 _PTL_IP3_2|_JTL|7 JJMIT AREA=2.5
I_PTL_IP3_2|_JTL|B1 0 _PTL_IP3_2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_IP3_2|_JTL|1 _PTL_IP3_2|A_PTL_RX _PTL_IP3_2|_JTL|1  2.067833848e-12
L_PTL_IP3_2|_JTL|2 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|4  2.067833848e-12
L_PTL_IP3_2|_JTL|3 _PTL_IP3_2|_JTL|4 _PTL_IP3_2|_JTL|6  2.067833848e-12
L_PTL_IP3_2|_JTL|4 _PTL_IP3_2|_JTL|6 IP3_2_OUT_RX  2.067833848e-12
L_PTL_IP3_2|_JTL|P1 _PTL_IP3_2|_JTL|2 0  2e-13
L_PTL_IP3_2|_JTL|P2 _PTL_IP3_2|_JTL|7 0  2e-13
L_PTL_IP3_2|_JTL|B1 _PTL_IP3_2|_JTL|5 _PTL_IP3_2|_JTL|4  2e-12
R_PTL_IP3_2|_JTL|B1 _PTL_IP3_2|_JTL|1 _PTL_IP3_2|_JTL|3  2.7439617672
R_PTL_IP3_2|_JTL|B2 _PTL_IP3_2|_JTL|6 _PTL_IP3_2|_JTL|8  2.7439617672
L_PTL_IP3_2|_JTL|RB1 _PTL_IP3_2|_JTL|3 0  1.750338398468e-12
L_PTL_IP3_2|_JTL|RB2 _PTL_IP3_2|_JTL|8 0  1.750338398468e-12
L_S0|I_1|B _S0|A1 _S0|I_1|MID  2e-12
I_S0|I_1|B 0 _S0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_3|B _S0|A3 _S0|I_3|MID  2e-12
I_S0|I_3|B 0 _S0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0|I_T|B _S0|T1 _S0|I_T|MID  2e-12
I_S0|I_T|B 0 _S0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_6|B _S0|Q1 _S0|I_6|MID  2e-12
I_S0|I_6|B 0 _S0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0|1|1 _S0|A1 _S0|1|MID_SERIES JJMIT AREA=2.5
L_S0|1|P _S0|1|MID_SERIES 0  2e-13
R_S0|1|B _S0|A1 _S0|1|MID_SHUNT  2.7439617672
L_S0|1|RB _S0|1|MID_SHUNT 0  1.550338398468e-12
B_S0|23|1 _S0|A2 _S0|A3 JJMIT AREA=1.7857142857142858
R_S0|23|B _S0|A2 _S0|23|MID_SHUNT  3.84154647408
L_S0|23|RB _S0|23|MID_SHUNT _S0|A3  2.1704737578552e-12
B_S0|3|1 _S0|A3 _S0|3|MID_SERIES JJMIT AREA=2.5
L_S0|3|P _S0|3|MID_SERIES 0  2e-13
R_S0|3|B _S0|A3 _S0|3|MID_SHUNT  2.7439617672
L_S0|3|RB _S0|3|MID_SHUNT 0  1.550338398468e-12
B_S0|4|1 _S0|A4 _S0|4|MID_SERIES JJMIT AREA=2.5
L_S0|4|P _S0|4|MID_SERIES 0  2e-13
R_S0|4|B _S0|A4 _S0|4|MID_SHUNT  2.7439617672
L_S0|4|RB _S0|4|MID_SHUNT 0  1.550338398468e-12
B_S0|T|1 _S0|T1 _S0|T|MID_SERIES JJMIT AREA=2.5
L_S0|T|P _S0|T|MID_SERIES 0  2e-13
R_S0|T|B _S0|T1 _S0|T|MID_SHUNT  2.7439617672
L_S0|T|RB _S0|T|MID_SHUNT 0  1.550338398468e-12
B_S0|45|1 _S0|T2 _S0|A4 JJMIT AREA=1.7857142857142858
R_S0|45|B _S0|T2 _S0|45|MID_SHUNT  3.84154647408
L_S0|45|RB _S0|45|MID_SHUNT _S0|A4  2.1704737578552e-12
B_S0|6|1 _S0|Q1 _S0|6|MID_SERIES JJMIT AREA=2.5
L_S0|6|P _S0|6|MID_SERIES 0  2e-13
R_S0|6|B _S0|Q1 _S0|6|MID_SHUNT  2.7439617672
L_S0|6|RB _S0|6|MID_SHUNT 0  1.550338398468e-12
L_S1|I_A1|B _S1|A1 _S1|I_A1|MID  2e-12
I_S1|I_A1|B 0 _S1|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_A3|B _S1|A3 _S1|I_A3|MID  2e-12
I_S1|I_A3|B 0 _S1|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B1|B _S1|B1 _S1|I_B1|MID  2e-12
I_S1|I_B1|B 0 _S1|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B3|B _S1|B3 _S1|I_B3|MID  2e-12
I_S1|I_B3|B 0 _S1|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_Q1|B _S1|Q1 _S1|I_Q1|MID  2e-12
I_S1|I_Q1|B 0 _S1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S1|A1|1 _S1|A1 _S1|A1|MID_SERIES JJMIT AREA=2.5
L_S1|A1|P _S1|A1|MID_SERIES 0  5e-13
R_S1|A1|B _S1|A1 _S1|A1|MID_SHUNT  2.7439617672
L_S1|A1|RB _S1|A1|MID_SHUNT 0  2.050338398468e-12
B_S1|A2|1 _S1|A2 _S1|A2|MID_SERIES JJMIT AREA=2.5
L_S1|A2|P _S1|A2|MID_SERIES 0  5e-13
R_S1|A2|B _S1|A2 _S1|A2|MID_SHUNT  2.7439617672
L_S1|A2|RB _S1|A2|MID_SHUNT 0  2.050338398468e-12
B_S1|A3|1 _S1|A2 _S1|A3|MID_SERIES JJMIT AREA=2.5
L_S1|A3|P _S1|A3|MID_SERIES _S1|A3  1.2e-12
R_S1|A3|B _S1|A2 _S1|A3|MID_SHUNT  2.7439617672
L_S1|A3|RB _S1|A3|MID_SHUNT _S1|A3  2.050338398468e-12
B_S1|B1|1 _S1|B1 _S1|B1|MID_SERIES JJMIT AREA=2.5
L_S1|B1|P _S1|B1|MID_SERIES 0  5e-13
R_S1|B1|B _S1|B1 _S1|B1|MID_SHUNT  2.7439617672
L_S1|B1|RB _S1|B1|MID_SHUNT 0  2.050338398468e-12
B_S1|B2|1 _S1|B2 _S1|B2|MID_SERIES JJMIT AREA=2.5
L_S1|B2|P _S1|B2|MID_SERIES 0  5e-13
R_S1|B2|B _S1|B2 _S1|B2|MID_SHUNT  2.7439617672
L_S1|B2|RB _S1|B2|MID_SHUNT 0  2.050338398468e-12
B_S1|B3|1 _S1|B2 _S1|B3|MID_SERIES JJMIT AREA=2.5
L_S1|B3|P _S1|B3|MID_SERIES _S1|B3  1.2e-12
R_S1|B3|B _S1|B2 _S1|B3|MID_SHUNT  2.7439617672
L_S1|B3|RB _S1|B3|MID_SHUNT _S1|B3  2.050338398468e-12
B_S1|T1|1 _S1|T1 _S1|T1|MID_SERIES JJMIT AREA=2.5
L_S1|T1|P _S1|T1|MID_SERIES 0  5e-13
R_S1|T1|B _S1|T1 _S1|T1|MID_SHUNT  2.7439617672
L_S1|T1|RB _S1|T1|MID_SHUNT 0  2.050338398468e-12
B_S1|T2|1 _S1|T2 _S1|ABTQ JJMIT AREA=2.0
R_S1|T2|B _S1|T2 _S1|T2|MID_SHUNT  3.429952209
L_S1|T2|RB _S1|T2|MID_SHUNT _S1|ABTQ  2.437922998085e-12
B_S1|AB|1 _S1|AB _S1|AB|MID_SERIES JJMIT AREA=1.5
L_S1|AB|P _S1|AB|MID_SERIES _S1|ABTQ  1.2e-12
R_S1|AB|B _S1|AB _S1|AB|MID_SHUNT  4.573269612
L_S1|AB|RB _S1|AB|MID_SHUNT _S1|ABTQ  3.08389733078e-12
B_S1|ABTQ|1 _S1|ABTQ _S1|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S1|ABTQ|P _S1|ABTQ|MID_SERIES 0  5e-13
R_S1|ABTQ|B _S1|ABTQ _S1|ABTQ|MID_SHUNT  3.6586156896
L_S1|ABTQ|RB _S1|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S1|Q1|1 _S1|Q1 _S1|Q1|MID_SERIES JJMIT AREA=2.5
L_S1|Q1|P _S1|Q1|MID_SERIES 0  5e-13
R_S1|Q1|B _S1|Q1 _S1|Q1|MID_SHUNT  2.7439617672
L_S1|Q1|RB _S1|Q1|MID_SHUNT 0  2.050338398468e-12
L_S2|I_A1|B _S2|A1 _S2|I_A1|MID  2e-12
I_S2|I_A1|B 0 _S2|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_A3|B _S2|A3 _S2|I_A3|MID  2e-12
I_S2|I_A3|B 0 _S2|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B1|B _S2|B1 _S2|I_B1|MID  2e-12
I_S2|I_B1|B 0 _S2|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B3|B _S2|B3 _S2|I_B3|MID  2e-12
I_S2|I_B3|B 0 _S2|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_Q1|B _S2|Q1 _S2|I_Q1|MID  2e-12
I_S2|I_Q1|B 0 _S2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S2|A1|1 _S2|A1 _S2|A1|MID_SERIES JJMIT AREA=2.5
L_S2|A1|P _S2|A1|MID_SERIES 0  5e-13
R_S2|A1|B _S2|A1 _S2|A1|MID_SHUNT  2.7439617672
L_S2|A1|RB _S2|A1|MID_SHUNT 0  2.050338398468e-12
B_S2|A2|1 _S2|A2 _S2|A2|MID_SERIES JJMIT AREA=2.5
L_S2|A2|P _S2|A2|MID_SERIES 0  5e-13
R_S2|A2|B _S2|A2 _S2|A2|MID_SHUNT  2.7439617672
L_S2|A2|RB _S2|A2|MID_SHUNT 0  2.050338398468e-12
B_S2|A3|1 _S2|A2 _S2|A3|MID_SERIES JJMIT AREA=2.5
L_S2|A3|P _S2|A3|MID_SERIES _S2|A3  1.2e-12
R_S2|A3|B _S2|A2 _S2|A3|MID_SHUNT  2.7439617672
L_S2|A3|RB _S2|A3|MID_SHUNT _S2|A3  2.050338398468e-12
B_S2|B1|1 _S2|B1 _S2|B1|MID_SERIES JJMIT AREA=2.5
L_S2|B1|P _S2|B1|MID_SERIES 0  5e-13
R_S2|B1|B _S2|B1 _S2|B1|MID_SHUNT  2.7439617672
L_S2|B1|RB _S2|B1|MID_SHUNT 0  2.050338398468e-12
B_S2|B2|1 _S2|B2 _S2|B2|MID_SERIES JJMIT AREA=2.5
L_S2|B2|P _S2|B2|MID_SERIES 0  5e-13
R_S2|B2|B _S2|B2 _S2|B2|MID_SHUNT  2.7439617672
L_S2|B2|RB _S2|B2|MID_SHUNT 0  2.050338398468e-12
B_S2|B3|1 _S2|B2 _S2|B3|MID_SERIES JJMIT AREA=2.5
L_S2|B3|P _S2|B3|MID_SERIES _S2|B3  1.2e-12
R_S2|B3|B _S2|B2 _S2|B3|MID_SHUNT  2.7439617672
L_S2|B3|RB _S2|B3|MID_SHUNT _S2|B3  2.050338398468e-12
B_S2|T1|1 _S2|T1 _S2|T1|MID_SERIES JJMIT AREA=2.5
L_S2|T1|P _S2|T1|MID_SERIES 0  5e-13
R_S2|T1|B _S2|T1 _S2|T1|MID_SHUNT  2.7439617672
L_S2|T1|RB _S2|T1|MID_SHUNT 0  2.050338398468e-12
B_S2|T2|1 _S2|T2 _S2|ABTQ JJMIT AREA=2.0
R_S2|T2|B _S2|T2 _S2|T2|MID_SHUNT  3.429952209
L_S2|T2|RB _S2|T2|MID_SHUNT _S2|ABTQ  2.437922998085e-12
B_S2|AB|1 _S2|AB _S2|AB|MID_SERIES JJMIT AREA=1.5
L_S2|AB|P _S2|AB|MID_SERIES _S2|ABTQ  1.2e-12
R_S2|AB|B _S2|AB _S2|AB|MID_SHUNT  4.573269612
L_S2|AB|RB _S2|AB|MID_SHUNT _S2|ABTQ  3.08389733078e-12
B_S2|ABTQ|1 _S2|ABTQ _S2|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S2|ABTQ|P _S2|ABTQ|MID_SERIES 0  5e-13
R_S2|ABTQ|B _S2|ABTQ _S2|ABTQ|MID_SHUNT  3.6586156896
L_S2|ABTQ|RB _S2|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S2|Q1|1 _S2|Q1 _S2|Q1|MID_SERIES JJMIT AREA=2.5
L_S2|Q1|P _S2|Q1|MID_SERIES 0  5e-13
R_S2|Q1|B _S2|Q1 _S2|Q1|MID_SHUNT  2.7439617672
L_S2|Q1|RB _S2|Q1|MID_SHUNT 0  2.050338398468e-12
L_S3|I_A1|B _S3|A1 _S3|I_A1|MID  2e-12
I_S3|I_A1|B 0 _S3|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_A3|B _S3|A3 _S3|I_A3|MID  2e-12
I_S3|I_A3|B 0 _S3|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B1|B _S3|B1 _S3|I_B1|MID  2e-12
I_S3|I_B1|B 0 _S3|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B3|B _S3|B3 _S3|I_B3|MID  2e-12
I_S3|I_B3|B 0 _S3|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_Q1|B _S3|Q1 _S3|I_Q1|MID  2e-12
I_S3|I_Q1|B 0 _S3|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S3|A1|1 _S3|A1 _S3|A1|MID_SERIES JJMIT AREA=2.5
L_S3|A1|P _S3|A1|MID_SERIES 0  5e-13
R_S3|A1|B _S3|A1 _S3|A1|MID_SHUNT  2.7439617672
L_S3|A1|RB _S3|A1|MID_SHUNT 0  2.050338398468e-12
B_S3|A2|1 _S3|A2 _S3|A2|MID_SERIES JJMIT AREA=2.5
L_S3|A2|P _S3|A2|MID_SERIES 0  5e-13
R_S3|A2|B _S3|A2 _S3|A2|MID_SHUNT  2.7439617672
L_S3|A2|RB _S3|A2|MID_SHUNT 0  2.050338398468e-12
B_S3|A3|1 _S3|A2 _S3|A3|MID_SERIES JJMIT AREA=2.5
L_S3|A3|P _S3|A3|MID_SERIES _S3|A3  1.2e-12
R_S3|A3|B _S3|A2 _S3|A3|MID_SHUNT  2.7439617672
L_S3|A3|RB _S3|A3|MID_SHUNT _S3|A3  2.050338398468e-12
B_S3|B1|1 _S3|B1 _S3|B1|MID_SERIES JJMIT AREA=2.5
L_S3|B1|P _S3|B1|MID_SERIES 0  5e-13
R_S3|B1|B _S3|B1 _S3|B1|MID_SHUNT  2.7439617672
L_S3|B1|RB _S3|B1|MID_SHUNT 0  2.050338398468e-12
B_S3|B2|1 _S3|B2 _S3|B2|MID_SERIES JJMIT AREA=2.5
L_S3|B2|P _S3|B2|MID_SERIES 0  5e-13
R_S3|B2|B _S3|B2 _S3|B2|MID_SHUNT  2.7439617672
L_S3|B2|RB _S3|B2|MID_SHUNT 0  2.050338398468e-12
B_S3|B3|1 _S3|B2 _S3|B3|MID_SERIES JJMIT AREA=2.5
L_S3|B3|P _S3|B3|MID_SERIES _S3|B3  1.2e-12
R_S3|B3|B _S3|B2 _S3|B3|MID_SHUNT  2.7439617672
L_S3|B3|RB _S3|B3|MID_SHUNT _S3|B3  2.050338398468e-12
B_S3|T1|1 _S3|T1 _S3|T1|MID_SERIES JJMIT AREA=2.5
L_S3|T1|P _S3|T1|MID_SERIES 0  5e-13
R_S3|T1|B _S3|T1 _S3|T1|MID_SHUNT  2.7439617672
L_S3|T1|RB _S3|T1|MID_SHUNT 0  2.050338398468e-12
B_S3|T2|1 _S3|T2 _S3|ABTQ JJMIT AREA=2.0
R_S3|T2|B _S3|T2 _S3|T2|MID_SHUNT  3.429952209
L_S3|T2|RB _S3|T2|MID_SHUNT _S3|ABTQ  2.437922998085e-12
B_S3|AB|1 _S3|AB _S3|AB|MID_SERIES JJMIT AREA=1.5
L_S3|AB|P _S3|AB|MID_SERIES _S3|ABTQ  1.2e-12
R_S3|AB|B _S3|AB _S3|AB|MID_SHUNT  4.573269612
L_S3|AB|RB _S3|AB|MID_SHUNT _S3|ABTQ  3.08389733078e-12
B_S3|ABTQ|1 _S3|ABTQ _S3|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S3|ABTQ|P _S3|ABTQ|MID_SERIES 0  5e-13
R_S3|ABTQ|B _S3|ABTQ _S3|ABTQ|MID_SHUNT  3.6586156896
L_S3|ABTQ|RB _S3|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S3|Q1|1 _S3|Q1 _S3|Q1|MID_SERIES JJMIT AREA=2.5
L_S3|Q1|P _S3|Q1|MID_SERIES 0  5e-13
R_S3|Q1|B _S3|Q1 _S3|Q1|MID_SHUNT  2.7439617672
L_S3|Q1|RB _S3|Q1|MID_SHUNT 0  2.050338398468e-12
L_S4|I_1|B _S4|A1 _S4|I_1|MID  2e-12
I_S4|I_1|B 0 _S4|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_3|B _S4|A3 _S4|I_3|MID  2e-12
I_S4|I_3|B 0 _S4|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S4|I_T|B _S4|T1 _S4|I_T|MID  2e-12
I_S4|I_T|B 0 _S4|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_6|B _S4|Q1 _S4|I_6|MID  2e-12
I_S4|I_6|B 0 _S4|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S4|1|1 _S4|A1 _S4|1|MID_SERIES JJMIT AREA=2.5
L_S4|1|P _S4|1|MID_SERIES 0  2e-13
R_S4|1|B _S4|A1 _S4|1|MID_SHUNT  2.7439617672
L_S4|1|RB _S4|1|MID_SHUNT 0  1.550338398468e-12
B_S4|23|1 _S4|A2 _S4|A3 JJMIT AREA=1.7857142857142858
R_S4|23|B _S4|A2 _S4|23|MID_SHUNT  3.84154647408
L_S4|23|RB _S4|23|MID_SHUNT _S4|A3  2.1704737578552e-12
B_S4|3|1 _S4|A3 _S4|3|MID_SERIES JJMIT AREA=2.5
L_S4|3|P _S4|3|MID_SERIES 0  2e-13
R_S4|3|B _S4|A3 _S4|3|MID_SHUNT  2.7439617672
L_S4|3|RB _S4|3|MID_SHUNT 0  1.550338398468e-12
B_S4|4|1 _S4|A4 _S4|4|MID_SERIES JJMIT AREA=2.5
L_S4|4|P _S4|4|MID_SERIES 0  2e-13
R_S4|4|B _S4|A4 _S4|4|MID_SHUNT  2.7439617672
L_S4|4|RB _S4|4|MID_SHUNT 0  1.550338398468e-12
B_S4|T|1 _S4|T1 _S4|T|MID_SERIES JJMIT AREA=2.5
L_S4|T|P _S4|T|MID_SERIES 0  2e-13
R_S4|T|B _S4|T1 _S4|T|MID_SHUNT  2.7439617672
L_S4|T|RB _S4|T|MID_SHUNT 0  1.550338398468e-12
B_S4|45|1 _S4|T2 _S4|A4 JJMIT AREA=1.7857142857142858
R_S4|45|B _S4|T2 _S4|45|MID_SHUNT  3.84154647408
L_S4|45|RB _S4|45|MID_SHUNT _S4|A4  2.1704737578552e-12
B_S4|6|1 _S4|Q1 _S4|6|MID_SERIES JJMIT AREA=2.5
L_S4|6|P _S4|6|MID_SERIES 0  2e-13
R_S4|6|B _S4|Q1 _S4|6|MID_SHUNT  2.7439617672
L_S4|6|RB _S4|6|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_A|I_D1|B I0|_SPL_A|D1 I0|_SPL_A|I_D1|MID  2e-12
II0|_SPL_A|I_D1|B 0 I0|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_D2|B I0|_SPL_A|D2 I0|_SPL_A|I_D2|MID  2e-12
II0|_SPL_A|I_D2|B 0 I0|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_A|I_Q1|B I0|_SPL_A|QA1 I0|_SPL_A|I_Q1|MID  2e-12
II0|_SPL_A|I_Q1|B 0 I0|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_Q2|B I0|_SPL_A|QB1 I0|_SPL_A|I_Q2|MID  2e-12
II0|_SPL_A|I_Q2|B 0 I0|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_A|1|1 I0|_SPL_A|D1 I0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|1|P I0|_SPL_A|1|MID_SERIES 0  2e-13
RI0|_SPL_A|1|B I0|_SPL_A|D1 I0|_SPL_A|1|MID_SHUNT  2.7439617672
LI0|_SPL_A|1|RB I0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|2|1 I0|_SPL_A|D2 I0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|2|P I0|_SPL_A|2|MID_SERIES 0  2e-13
RI0|_SPL_A|2|B I0|_SPL_A|D2 I0|_SPL_A|2|MID_SHUNT  2.7439617672
LI0|_SPL_A|2|RB I0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|A|1 I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|A|P I0|_SPL_A|A|MID_SERIES 0  2e-13
RI0|_SPL_A|A|B I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SHUNT  2.7439617672
LI0|_SPL_A|A|RB I0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|B|1 I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|B|P I0|_SPL_A|B|MID_SERIES 0  2e-13
RI0|_SPL_A|B|B I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SHUNT  2.7439617672
LI0|_SPL_A|B|RB I0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_B|I_D1|B I0|_SPL_B|D1 I0|_SPL_B|I_D1|MID  2e-12
II0|_SPL_B|I_D1|B 0 I0|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_D2|B I0|_SPL_B|D2 I0|_SPL_B|I_D2|MID  2e-12
II0|_SPL_B|I_D2|B 0 I0|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_B|I_Q1|B I0|_SPL_B|QA1 I0|_SPL_B|I_Q1|MID  2e-12
II0|_SPL_B|I_Q1|B 0 I0|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_Q2|B I0|_SPL_B|QB1 I0|_SPL_B|I_Q2|MID  2e-12
II0|_SPL_B|I_Q2|B 0 I0|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_B|1|1 I0|_SPL_B|D1 I0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|1|P I0|_SPL_B|1|MID_SERIES 0  2e-13
RI0|_SPL_B|1|B I0|_SPL_B|D1 I0|_SPL_B|1|MID_SHUNT  2.7439617672
LI0|_SPL_B|1|RB I0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|2|1 I0|_SPL_B|D2 I0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|2|P I0|_SPL_B|2|MID_SERIES 0  2e-13
RI0|_SPL_B|2|B I0|_SPL_B|D2 I0|_SPL_B|2|MID_SHUNT  2.7439617672
LI0|_SPL_B|2|RB I0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|A|1 I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|A|P I0|_SPL_B|A|MID_SERIES 0  2e-13
RI0|_SPL_B|A|B I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SHUNT  2.7439617672
LI0|_SPL_B|A|RB I0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|B|1 I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|B|P I0|_SPL_B|B|MID_SERIES 0  2e-13
RI0|_SPL_B|B|B I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SHUNT  2.7439617672
LI0|_SPL_B|B|RB I0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_A|I_1|B I0|_DFF_A|A1 I0|_DFF_A|I_1|MID  2e-12
II0|_DFF_A|I_1|B 0 I0|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_3|B I0|_DFF_A|A3 I0|_DFF_A|I_3|MID  2e-12
II0|_DFF_A|I_3|B 0 I0|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_A|I_T|B I0|_DFF_A|T1 I0|_DFF_A|I_T|MID  2e-12
II0|_DFF_A|I_T|B 0 I0|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_6|B I0|_DFF_A|Q1 I0|_DFF_A|I_6|MID  2e-12
II0|_DFF_A|I_6|B 0 I0|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_A|1|1 I0|_DFF_A|A1 I0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|1|P I0|_DFF_A|1|MID_SERIES 0  2e-13
RI0|_DFF_A|1|B I0|_DFF_A|A1 I0|_DFF_A|1|MID_SHUNT  2.7439617672
LI0|_DFF_A|1|RB I0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|23|1 I0|_DFF_A|A2 I0|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|23|B I0|_DFF_A|A2 I0|_DFF_A|23|MID_SHUNT  3.84154647408
LI0|_DFF_A|23|RB I0|_DFF_A|23|MID_SHUNT I0|_DFF_A|A3  2.1704737578552e-12
BI0|_DFF_A|3|1 I0|_DFF_A|A3 I0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|3|P I0|_DFF_A|3|MID_SERIES 0  2e-13
RI0|_DFF_A|3|B I0|_DFF_A|A3 I0|_DFF_A|3|MID_SHUNT  2.7439617672
LI0|_DFF_A|3|RB I0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|4|1 I0|_DFF_A|A4 I0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|4|P I0|_DFF_A|4|MID_SERIES 0  2e-13
RI0|_DFF_A|4|B I0|_DFF_A|A4 I0|_DFF_A|4|MID_SHUNT  2.7439617672
LI0|_DFF_A|4|RB I0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|T|1 I0|_DFF_A|T1 I0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|T|P I0|_DFF_A|T|MID_SERIES 0  2e-13
RI0|_DFF_A|T|B I0|_DFF_A|T1 I0|_DFF_A|T|MID_SHUNT  2.7439617672
LI0|_DFF_A|T|RB I0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|45|1 I0|_DFF_A|T2 I0|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|45|B I0|_DFF_A|T2 I0|_DFF_A|45|MID_SHUNT  3.84154647408
LI0|_DFF_A|45|RB I0|_DFF_A|45|MID_SHUNT I0|_DFF_A|A4  2.1704737578552e-12
BI0|_DFF_A|6|1 I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|6|P I0|_DFF_A|6|MID_SERIES 0  2e-13
RI0|_DFF_A|6|B I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SHUNT  2.7439617672
LI0|_DFF_A|6|RB I0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_B|I_1|B I0|_DFF_B|A1 I0|_DFF_B|I_1|MID  2e-12
II0|_DFF_B|I_1|B 0 I0|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_3|B I0|_DFF_B|A3 I0|_DFF_B|I_3|MID  2e-12
II0|_DFF_B|I_3|B 0 I0|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_B|I_T|B I0|_DFF_B|T1 I0|_DFF_B|I_T|MID  2e-12
II0|_DFF_B|I_T|B 0 I0|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_6|B I0|_DFF_B|Q1 I0|_DFF_B|I_6|MID  2e-12
II0|_DFF_B|I_6|B 0 I0|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_B|1|1 I0|_DFF_B|A1 I0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|1|P I0|_DFF_B|1|MID_SERIES 0  2e-13
RI0|_DFF_B|1|B I0|_DFF_B|A1 I0|_DFF_B|1|MID_SHUNT  2.7439617672
LI0|_DFF_B|1|RB I0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|23|1 I0|_DFF_B|A2 I0|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|23|B I0|_DFF_B|A2 I0|_DFF_B|23|MID_SHUNT  3.84154647408
LI0|_DFF_B|23|RB I0|_DFF_B|23|MID_SHUNT I0|_DFF_B|A3  2.1704737578552e-12
BI0|_DFF_B|3|1 I0|_DFF_B|A3 I0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|3|P I0|_DFF_B|3|MID_SERIES 0  2e-13
RI0|_DFF_B|3|B I0|_DFF_B|A3 I0|_DFF_B|3|MID_SHUNT  2.7439617672
LI0|_DFF_B|3|RB I0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|4|1 I0|_DFF_B|A4 I0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|4|P I0|_DFF_B|4|MID_SERIES 0  2e-13
RI0|_DFF_B|4|B I0|_DFF_B|A4 I0|_DFF_B|4|MID_SHUNT  2.7439617672
LI0|_DFF_B|4|RB I0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|T|1 I0|_DFF_B|T1 I0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|T|P I0|_DFF_B|T|MID_SERIES 0  2e-13
RI0|_DFF_B|T|B I0|_DFF_B|T1 I0|_DFF_B|T|MID_SHUNT  2.7439617672
LI0|_DFF_B|T|RB I0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|45|1 I0|_DFF_B|T2 I0|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|45|B I0|_DFF_B|T2 I0|_DFF_B|45|MID_SHUNT  3.84154647408
LI0|_DFF_B|45|RB I0|_DFF_B|45|MID_SHUNT I0|_DFF_B|A4  2.1704737578552e-12
BI0|_DFF_B|6|1 I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|6|P I0|_DFF_B|6|MID_SERIES 0  2e-13
RI0|_DFF_B|6|B I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SHUNT  2.7439617672
LI0|_DFF_B|6|RB I0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI0|_XOR|I_A1|B I0|_XOR|A1 I0|_XOR|I_A1|MID  2e-12
II0|_XOR|I_A1|B 0 I0|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_A3|B I0|_XOR|A3 I0|_XOR|I_A3|MID  2e-12
II0|_XOR|I_A3|B 0 I0|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B1|B I0|_XOR|B1 I0|_XOR|I_B1|MID  2e-12
II0|_XOR|I_B1|B 0 I0|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B3|B I0|_XOR|B3 I0|_XOR|I_B3|MID  2e-12
II0|_XOR|I_B3|B 0 I0|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_Q1|B I0|_XOR|Q1 I0|_XOR|I_Q1|MID  2e-12
II0|_XOR|I_Q1|B 0 I0|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_XOR|A1|1 I0|_XOR|A1 I0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A1|P I0|_XOR|A1|MID_SERIES 0  5e-13
RI0|_XOR|A1|B I0|_XOR|A1 I0|_XOR|A1|MID_SHUNT  2.7439617672
LI0|_XOR|A1|RB I0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A2|1 I0|_XOR|A2 I0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A2|P I0|_XOR|A2|MID_SERIES 0  5e-13
RI0|_XOR|A2|B I0|_XOR|A2 I0|_XOR|A2|MID_SHUNT  2.7439617672
LI0|_XOR|A2|RB I0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A3|1 I0|_XOR|A2 I0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A3|P I0|_XOR|A3|MID_SERIES I0|_XOR|A3  1.2e-12
RI0|_XOR|A3|B I0|_XOR|A2 I0|_XOR|A3|MID_SHUNT  2.7439617672
LI0|_XOR|A3|RB I0|_XOR|A3|MID_SHUNT I0|_XOR|A3  2.050338398468e-12
BI0|_XOR|B1|1 I0|_XOR|B1 I0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B1|P I0|_XOR|B1|MID_SERIES 0  5e-13
RI0|_XOR|B1|B I0|_XOR|B1 I0|_XOR|B1|MID_SHUNT  2.7439617672
LI0|_XOR|B1|RB I0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B2|1 I0|_XOR|B2 I0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B2|P I0|_XOR|B2|MID_SERIES 0  5e-13
RI0|_XOR|B2|B I0|_XOR|B2 I0|_XOR|B2|MID_SHUNT  2.7439617672
LI0|_XOR|B2|RB I0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B3|1 I0|_XOR|B2 I0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B3|P I0|_XOR|B3|MID_SERIES I0|_XOR|B3  1.2e-12
RI0|_XOR|B3|B I0|_XOR|B2 I0|_XOR|B3|MID_SHUNT  2.7439617672
LI0|_XOR|B3|RB I0|_XOR|B3|MID_SHUNT I0|_XOR|B3  2.050338398468e-12
BI0|_XOR|T1|1 I0|_XOR|T1 I0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|T1|P I0|_XOR|T1|MID_SERIES 0  5e-13
RI0|_XOR|T1|B I0|_XOR|T1 I0|_XOR|T1|MID_SHUNT  2.7439617672
LI0|_XOR|T1|RB I0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|T2|1 I0|_XOR|T2 I0|_XOR|ABTQ JJMIT AREA=2.0
RI0|_XOR|T2|B I0|_XOR|T2 I0|_XOR|T2|MID_SHUNT  3.429952209
LI0|_XOR|T2|RB I0|_XOR|T2|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|AB|1 I0|_XOR|AB I0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI0|_XOR|AB|P I0|_XOR|AB|MID_SERIES I0|_XOR|ABTQ  1.2e-12
RI0|_XOR|AB|B I0|_XOR|AB I0|_XOR|AB|MID_SHUNT  3.429952209
LI0|_XOR|AB|RB I0|_XOR|AB|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|ABTQ|1 I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|ABTQ|P I0|_XOR|ABTQ|MID_SERIES 0  5e-13
RI0|_XOR|ABTQ|B I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI0|_XOR|ABTQ|RB I0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|Q1|1 I0|_XOR|Q1 I0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|Q1|P I0|_XOR|Q1|MID_SERIES 0  5e-13
RI0|_XOR|Q1|B I0|_XOR|Q1 I0|_XOR|Q1|MID_SHUNT  2.7439617672
LI0|_XOR|Q1|RB I0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI0|_AND|I_A1|B I0|_AND|A1 I0|_AND|I_A1|MID  2e-12
II0|_AND|I_A1|B 0 I0|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_B1|B I0|_AND|B1 I0|_AND|I_B1|MID  2e-12
II0|_AND|I_B1|B 0 I0|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q3|B I0|_AND|Q3 I0|_AND|I_Q3|MID  2e-12
II0|_AND|I_Q3|B 0 I0|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0|_AND|I_Q2|B I0|_AND|Q2 I0|_AND|I_Q2|MID  2e-12
II0|_AND|I_Q2|B 0 I0|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q1|B I0|_AND|Q1 I0|_AND|I_Q1|MID  2e-12
II0|_AND|I_Q1|B 0 I0|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_AND|A1|1 I0|_AND|A1 I0|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A1|P I0|_AND|A1|MID_SERIES 0  2e-13
RI0|_AND|A1|B I0|_AND|A1 I0|_AND|A1|MID_SHUNT  2.7439617672
LI0|_AND|A1|RB I0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A2|1 I0|_AND|A2 I0|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A2|P I0|_AND|A2|MID_SERIES 0  2e-13
RI0|_AND|A2|B I0|_AND|A2 I0|_AND|A2|MID_SHUNT  2.7439617672
LI0|_AND|A2|RB I0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A12|1 I0|_AND|A2 I0|_AND|A3 JJMIT AREA=1.7857142857142858
RI0|_AND|A12|B I0|_AND|A2 I0|_AND|A12|MID_SHUNT  3.84154647408
LI0|_AND|A12|RB I0|_AND|A12|MID_SHUNT I0|_AND|A3  2.1704737578552e-12
BI0|_AND|B1|1 I0|_AND|B1 I0|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B1|P I0|_AND|B1|MID_SERIES 0  2e-13
RI0|_AND|B1|B I0|_AND|B1 I0|_AND|B1|MID_SHUNT  2.7439617672
LI0|_AND|B1|RB I0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B2|1 I0|_AND|B2 I0|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B2|P I0|_AND|B2|MID_SERIES 0  2e-13
RI0|_AND|B2|B I0|_AND|B2 I0|_AND|B2|MID_SHUNT  2.7439617672
LI0|_AND|B2|RB I0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B12|1 I0|_AND|B2 I0|_AND|B3 JJMIT AREA=1.7857142857142858
RI0|_AND|B12|B I0|_AND|B2 I0|_AND|B12|MID_SHUNT  3.84154647408
LI0|_AND|B12|RB I0|_AND|B12|MID_SHUNT I0|_AND|B3  2.1704737578552e-12
BI0|_AND|Q2|1 I0|_AND|Q2 I0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q2|P I0|_AND|Q2|MID_SERIES 0  2e-13
RI0|_AND|Q2|B I0|_AND|Q2 I0|_AND|Q2|MID_SHUNT  2.7439617672
LI0|_AND|Q2|RB I0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|Q1|1 I0|_AND|Q1 I0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q1|P I0|_AND|Q1|MID_SERIES 0  2e-13
RI0|_AND|Q1|B I0|_AND|Q1 I0|_AND|Q1|MID_SHUNT  2.7439617672
LI0|_AND|Q1|RB I0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_A|I_D1|B I1|_SPL_A|D1 I1|_SPL_A|I_D1|MID  2e-12
II1|_SPL_A|I_D1|B 0 I1|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_D2|B I1|_SPL_A|D2 I1|_SPL_A|I_D2|MID  2e-12
II1|_SPL_A|I_D2|B 0 I1|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_A|I_Q1|B I1|_SPL_A|QA1 I1|_SPL_A|I_Q1|MID  2e-12
II1|_SPL_A|I_Q1|B 0 I1|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_Q2|B I1|_SPL_A|QB1 I1|_SPL_A|I_Q2|MID  2e-12
II1|_SPL_A|I_Q2|B 0 I1|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_A|1|1 I1|_SPL_A|D1 I1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|1|P I1|_SPL_A|1|MID_SERIES 0  2e-13
RI1|_SPL_A|1|B I1|_SPL_A|D1 I1|_SPL_A|1|MID_SHUNT  2.7439617672
LI1|_SPL_A|1|RB I1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|2|1 I1|_SPL_A|D2 I1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|2|P I1|_SPL_A|2|MID_SERIES 0  2e-13
RI1|_SPL_A|2|B I1|_SPL_A|D2 I1|_SPL_A|2|MID_SHUNT  2.7439617672
LI1|_SPL_A|2|RB I1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|A|1 I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|A|P I1|_SPL_A|A|MID_SERIES 0  2e-13
RI1|_SPL_A|A|B I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SHUNT  2.7439617672
LI1|_SPL_A|A|RB I1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|B|1 I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|B|P I1|_SPL_A|B|MID_SERIES 0  2e-13
RI1|_SPL_A|B|B I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SHUNT  2.7439617672
LI1|_SPL_A|B|RB I1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_B|I_D1|B I1|_SPL_B|D1 I1|_SPL_B|I_D1|MID  2e-12
II1|_SPL_B|I_D1|B 0 I1|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_D2|B I1|_SPL_B|D2 I1|_SPL_B|I_D2|MID  2e-12
II1|_SPL_B|I_D2|B 0 I1|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_B|I_Q1|B I1|_SPL_B|QA1 I1|_SPL_B|I_Q1|MID  2e-12
II1|_SPL_B|I_Q1|B 0 I1|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_Q2|B I1|_SPL_B|QB1 I1|_SPL_B|I_Q2|MID  2e-12
II1|_SPL_B|I_Q2|B 0 I1|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_B|1|1 I1|_SPL_B|D1 I1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|1|P I1|_SPL_B|1|MID_SERIES 0  2e-13
RI1|_SPL_B|1|B I1|_SPL_B|D1 I1|_SPL_B|1|MID_SHUNT  2.7439617672
LI1|_SPL_B|1|RB I1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|2|1 I1|_SPL_B|D2 I1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|2|P I1|_SPL_B|2|MID_SERIES 0  2e-13
RI1|_SPL_B|2|B I1|_SPL_B|D2 I1|_SPL_B|2|MID_SHUNT  2.7439617672
LI1|_SPL_B|2|RB I1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|A|1 I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|A|P I1|_SPL_B|A|MID_SERIES 0  2e-13
RI1|_SPL_B|A|B I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SHUNT  2.7439617672
LI1|_SPL_B|A|RB I1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|B|1 I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|B|P I1|_SPL_B|B|MID_SERIES 0  2e-13
RI1|_SPL_B|B|B I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SHUNT  2.7439617672
LI1|_SPL_B|B|RB I1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_A|I_1|B I1|_DFF_A|A1 I1|_DFF_A|I_1|MID  2e-12
II1|_DFF_A|I_1|B 0 I1|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_3|B I1|_DFF_A|A3 I1|_DFF_A|I_3|MID  2e-12
II1|_DFF_A|I_3|B 0 I1|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_A|I_T|B I1|_DFF_A|T1 I1|_DFF_A|I_T|MID  2e-12
II1|_DFF_A|I_T|B 0 I1|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_6|B I1|_DFF_A|Q1 I1|_DFF_A|I_6|MID  2e-12
II1|_DFF_A|I_6|B 0 I1|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_A|1|1 I1|_DFF_A|A1 I1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|1|P I1|_DFF_A|1|MID_SERIES 0  2e-13
RI1|_DFF_A|1|B I1|_DFF_A|A1 I1|_DFF_A|1|MID_SHUNT  2.7439617672
LI1|_DFF_A|1|RB I1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|23|1 I1|_DFF_A|A2 I1|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|23|B I1|_DFF_A|A2 I1|_DFF_A|23|MID_SHUNT  3.84154647408
LI1|_DFF_A|23|RB I1|_DFF_A|23|MID_SHUNT I1|_DFF_A|A3  2.1704737578552e-12
BI1|_DFF_A|3|1 I1|_DFF_A|A3 I1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|3|P I1|_DFF_A|3|MID_SERIES 0  2e-13
RI1|_DFF_A|3|B I1|_DFF_A|A3 I1|_DFF_A|3|MID_SHUNT  2.7439617672
LI1|_DFF_A|3|RB I1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|4|1 I1|_DFF_A|A4 I1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|4|P I1|_DFF_A|4|MID_SERIES 0  2e-13
RI1|_DFF_A|4|B I1|_DFF_A|A4 I1|_DFF_A|4|MID_SHUNT  2.7439617672
LI1|_DFF_A|4|RB I1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|T|1 I1|_DFF_A|T1 I1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|T|P I1|_DFF_A|T|MID_SERIES 0  2e-13
RI1|_DFF_A|T|B I1|_DFF_A|T1 I1|_DFF_A|T|MID_SHUNT  2.7439617672
LI1|_DFF_A|T|RB I1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|45|1 I1|_DFF_A|T2 I1|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|45|B I1|_DFF_A|T2 I1|_DFF_A|45|MID_SHUNT  3.84154647408
LI1|_DFF_A|45|RB I1|_DFF_A|45|MID_SHUNT I1|_DFF_A|A4  2.1704737578552e-12
BI1|_DFF_A|6|1 I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|6|P I1|_DFF_A|6|MID_SERIES 0  2e-13
RI1|_DFF_A|6|B I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SHUNT  2.7439617672
LI1|_DFF_A|6|RB I1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_B|I_1|B I1|_DFF_B|A1 I1|_DFF_B|I_1|MID  2e-12
II1|_DFF_B|I_1|B 0 I1|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_3|B I1|_DFF_B|A3 I1|_DFF_B|I_3|MID  2e-12
II1|_DFF_B|I_3|B 0 I1|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_B|I_T|B I1|_DFF_B|T1 I1|_DFF_B|I_T|MID  2e-12
II1|_DFF_B|I_T|B 0 I1|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_6|B I1|_DFF_B|Q1 I1|_DFF_B|I_6|MID  2e-12
II1|_DFF_B|I_6|B 0 I1|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_B|1|1 I1|_DFF_B|A1 I1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|1|P I1|_DFF_B|1|MID_SERIES 0  2e-13
RI1|_DFF_B|1|B I1|_DFF_B|A1 I1|_DFF_B|1|MID_SHUNT  2.7439617672
LI1|_DFF_B|1|RB I1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|23|1 I1|_DFF_B|A2 I1|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|23|B I1|_DFF_B|A2 I1|_DFF_B|23|MID_SHUNT  3.84154647408
LI1|_DFF_B|23|RB I1|_DFF_B|23|MID_SHUNT I1|_DFF_B|A3  2.1704737578552e-12
BI1|_DFF_B|3|1 I1|_DFF_B|A3 I1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|3|P I1|_DFF_B|3|MID_SERIES 0  2e-13
RI1|_DFF_B|3|B I1|_DFF_B|A3 I1|_DFF_B|3|MID_SHUNT  2.7439617672
LI1|_DFF_B|3|RB I1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|4|1 I1|_DFF_B|A4 I1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|4|P I1|_DFF_B|4|MID_SERIES 0  2e-13
RI1|_DFF_B|4|B I1|_DFF_B|A4 I1|_DFF_B|4|MID_SHUNT  2.7439617672
LI1|_DFF_B|4|RB I1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|T|1 I1|_DFF_B|T1 I1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|T|P I1|_DFF_B|T|MID_SERIES 0  2e-13
RI1|_DFF_B|T|B I1|_DFF_B|T1 I1|_DFF_B|T|MID_SHUNT  2.7439617672
LI1|_DFF_B|T|RB I1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|45|1 I1|_DFF_B|T2 I1|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|45|B I1|_DFF_B|T2 I1|_DFF_B|45|MID_SHUNT  3.84154647408
LI1|_DFF_B|45|RB I1|_DFF_B|45|MID_SHUNT I1|_DFF_B|A4  2.1704737578552e-12
BI1|_DFF_B|6|1 I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|6|P I1|_DFF_B|6|MID_SERIES 0  2e-13
RI1|_DFF_B|6|B I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SHUNT  2.7439617672
LI1|_DFF_B|6|RB I1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI1|_XOR|I_A1|B I1|_XOR|A1 I1|_XOR|I_A1|MID  2e-12
II1|_XOR|I_A1|B 0 I1|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_A3|B I1|_XOR|A3 I1|_XOR|I_A3|MID  2e-12
II1|_XOR|I_A3|B 0 I1|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B1|B I1|_XOR|B1 I1|_XOR|I_B1|MID  2e-12
II1|_XOR|I_B1|B 0 I1|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B3|B I1|_XOR|B3 I1|_XOR|I_B3|MID  2e-12
II1|_XOR|I_B3|B 0 I1|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_Q1|B I1|_XOR|Q1 I1|_XOR|I_Q1|MID  2e-12
II1|_XOR|I_Q1|B 0 I1|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_XOR|A1|1 I1|_XOR|A1 I1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A1|P I1|_XOR|A1|MID_SERIES 0  5e-13
RI1|_XOR|A1|B I1|_XOR|A1 I1|_XOR|A1|MID_SHUNT  2.7439617672
LI1|_XOR|A1|RB I1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A2|1 I1|_XOR|A2 I1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A2|P I1|_XOR|A2|MID_SERIES 0  5e-13
RI1|_XOR|A2|B I1|_XOR|A2 I1|_XOR|A2|MID_SHUNT  2.7439617672
LI1|_XOR|A2|RB I1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A3|1 I1|_XOR|A2 I1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A3|P I1|_XOR|A3|MID_SERIES I1|_XOR|A3  1.2e-12
RI1|_XOR|A3|B I1|_XOR|A2 I1|_XOR|A3|MID_SHUNT  2.7439617672
LI1|_XOR|A3|RB I1|_XOR|A3|MID_SHUNT I1|_XOR|A3  2.050338398468e-12
BI1|_XOR|B1|1 I1|_XOR|B1 I1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B1|P I1|_XOR|B1|MID_SERIES 0  5e-13
RI1|_XOR|B1|B I1|_XOR|B1 I1|_XOR|B1|MID_SHUNT  2.7439617672
LI1|_XOR|B1|RB I1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B2|1 I1|_XOR|B2 I1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B2|P I1|_XOR|B2|MID_SERIES 0  5e-13
RI1|_XOR|B2|B I1|_XOR|B2 I1|_XOR|B2|MID_SHUNT  2.7439617672
LI1|_XOR|B2|RB I1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B3|1 I1|_XOR|B2 I1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B3|P I1|_XOR|B3|MID_SERIES I1|_XOR|B3  1.2e-12
RI1|_XOR|B3|B I1|_XOR|B2 I1|_XOR|B3|MID_SHUNT  2.7439617672
LI1|_XOR|B3|RB I1|_XOR|B3|MID_SHUNT I1|_XOR|B3  2.050338398468e-12
BI1|_XOR|T1|1 I1|_XOR|T1 I1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|T1|P I1|_XOR|T1|MID_SERIES 0  5e-13
RI1|_XOR|T1|B I1|_XOR|T1 I1|_XOR|T1|MID_SHUNT  2.7439617672
LI1|_XOR|T1|RB I1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|T2|1 I1|_XOR|T2 I1|_XOR|ABTQ JJMIT AREA=2.0
RI1|_XOR|T2|B I1|_XOR|T2 I1|_XOR|T2|MID_SHUNT  3.429952209
LI1|_XOR|T2|RB I1|_XOR|T2|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|AB|1 I1|_XOR|AB I1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI1|_XOR|AB|P I1|_XOR|AB|MID_SERIES I1|_XOR|ABTQ  1.2e-12
RI1|_XOR|AB|B I1|_XOR|AB I1|_XOR|AB|MID_SHUNT  3.429952209
LI1|_XOR|AB|RB I1|_XOR|AB|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|ABTQ|1 I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|ABTQ|P I1|_XOR|ABTQ|MID_SERIES 0  5e-13
RI1|_XOR|ABTQ|B I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI1|_XOR|ABTQ|RB I1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|Q1|1 I1|_XOR|Q1 I1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|Q1|P I1|_XOR|Q1|MID_SERIES 0  5e-13
RI1|_XOR|Q1|B I1|_XOR|Q1 I1|_XOR|Q1|MID_SHUNT  2.7439617672
LI1|_XOR|Q1|RB I1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI1|_AND|I_A1|B I1|_AND|A1 I1|_AND|I_A1|MID  2e-12
II1|_AND|I_A1|B 0 I1|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_B1|B I1|_AND|B1 I1|_AND|I_B1|MID  2e-12
II1|_AND|I_B1|B 0 I1|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q3|B I1|_AND|Q3 I1|_AND|I_Q3|MID  2e-12
II1|_AND|I_Q3|B 0 I1|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1|_AND|I_Q2|B I1|_AND|Q2 I1|_AND|I_Q2|MID  2e-12
II1|_AND|I_Q2|B 0 I1|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q1|B I1|_AND|Q1 I1|_AND|I_Q1|MID  2e-12
II1|_AND|I_Q1|B 0 I1|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_AND|A1|1 I1|_AND|A1 I1|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A1|P I1|_AND|A1|MID_SERIES 0  2e-13
RI1|_AND|A1|B I1|_AND|A1 I1|_AND|A1|MID_SHUNT  2.7439617672
LI1|_AND|A1|RB I1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A2|1 I1|_AND|A2 I1|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A2|P I1|_AND|A2|MID_SERIES 0  2e-13
RI1|_AND|A2|B I1|_AND|A2 I1|_AND|A2|MID_SHUNT  2.7439617672
LI1|_AND|A2|RB I1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A12|1 I1|_AND|A2 I1|_AND|A3 JJMIT AREA=1.7857142857142858
RI1|_AND|A12|B I1|_AND|A2 I1|_AND|A12|MID_SHUNT  3.84154647408
LI1|_AND|A12|RB I1|_AND|A12|MID_SHUNT I1|_AND|A3  2.1704737578552e-12
BI1|_AND|B1|1 I1|_AND|B1 I1|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B1|P I1|_AND|B1|MID_SERIES 0  2e-13
RI1|_AND|B1|B I1|_AND|B1 I1|_AND|B1|MID_SHUNT  2.7439617672
LI1|_AND|B1|RB I1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B2|1 I1|_AND|B2 I1|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B2|P I1|_AND|B2|MID_SERIES 0  2e-13
RI1|_AND|B2|B I1|_AND|B2 I1|_AND|B2|MID_SHUNT  2.7439617672
LI1|_AND|B2|RB I1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B12|1 I1|_AND|B2 I1|_AND|B3 JJMIT AREA=1.7857142857142858
RI1|_AND|B12|B I1|_AND|B2 I1|_AND|B12|MID_SHUNT  3.84154647408
LI1|_AND|B12|RB I1|_AND|B12|MID_SHUNT I1|_AND|B3  2.1704737578552e-12
BI1|_AND|Q2|1 I1|_AND|Q2 I1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q2|P I1|_AND|Q2|MID_SERIES 0  2e-13
RI1|_AND|Q2|B I1|_AND|Q2 I1|_AND|Q2|MID_SHUNT  2.7439617672
LI1|_AND|Q2|RB I1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|Q1|1 I1|_AND|Q1 I1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q1|P I1|_AND|Q1|MID_SERIES 0  2e-13
RI1|_AND|Q1|B I1|_AND|Q1 I1|_AND|Q1|MID_SHUNT  2.7439617672
LI1|_AND|Q1|RB I1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_A|I_D1|B I2|_SPL_A|D1 I2|_SPL_A|I_D1|MID  2e-12
II2|_SPL_A|I_D1|B 0 I2|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_D2|B I2|_SPL_A|D2 I2|_SPL_A|I_D2|MID  2e-12
II2|_SPL_A|I_D2|B 0 I2|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_A|I_Q1|B I2|_SPL_A|QA1 I2|_SPL_A|I_Q1|MID  2e-12
II2|_SPL_A|I_Q1|B 0 I2|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_Q2|B I2|_SPL_A|QB1 I2|_SPL_A|I_Q2|MID  2e-12
II2|_SPL_A|I_Q2|B 0 I2|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_A|1|1 I2|_SPL_A|D1 I2|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|1|P I2|_SPL_A|1|MID_SERIES 0  2e-13
RI2|_SPL_A|1|B I2|_SPL_A|D1 I2|_SPL_A|1|MID_SHUNT  2.7439617672
LI2|_SPL_A|1|RB I2|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|2|1 I2|_SPL_A|D2 I2|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|2|P I2|_SPL_A|2|MID_SERIES 0  2e-13
RI2|_SPL_A|2|B I2|_SPL_A|D2 I2|_SPL_A|2|MID_SHUNT  2.7439617672
LI2|_SPL_A|2|RB I2|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|A|1 I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|A|P I2|_SPL_A|A|MID_SERIES 0  2e-13
RI2|_SPL_A|A|B I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SHUNT  2.7439617672
LI2|_SPL_A|A|RB I2|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|B|1 I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|B|P I2|_SPL_A|B|MID_SERIES 0  2e-13
RI2|_SPL_A|B|B I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SHUNT  2.7439617672
LI2|_SPL_A|B|RB I2|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_B|I_D1|B I2|_SPL_B|D1 I2|_SPL_B|I_D1|MID  2e-12
II2|_SPL_B|I_D1|B 0 I2|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_D2|B I2|_SPL_B|D2 I2|_SPL_B|I_D2|MID  2e-12
II2|_SPL_B|I_D2|B 0 I2|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_B|I_Q1|B I2|_SPL_B|QA1 I2|_SPL_B|I_Q1|MID  2e-12
II2|_SPL_B|I_Q1|B 0 I2|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_Q2|B I2|_SPL_B|QB1 I2|_SPL_B|I_Q2|MID  2e-12
II2|_SPL_B|I_Q2|B 0 I2|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_B|1|1 I2|_SPL_B|D1 I2|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|1|P I2|_SPL_B|1|MID_SERIES 0  2e-13
RI2|_SPL_B|1|B I2|_SPL_B|D1 I2|_SPL_B|1|MID_SHUNT  2.7439617672
LI2|_SPL_B|1|RB I2|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|2|1 I2|_SPL_B|D2 I2|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|2|P I2|_SPL_B|2|MID_SERIES 0  2e-13
RI2|_SPL_B|2|B I2|_SPL_B|D2 I2|_SPL_B|2|MID_SHUNT  2.7439617672
LI2|_SPL_B|2|RB I2|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|A|1 I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|A|P I2|_SPL_B|A|MID_SERIES 0  2e-13
RI2|_SPL_B|A|B I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SHUNT  2.7439617672
LI2|_SPL_B|A|RB I2|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|B|1 I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|B|P I2|_SPL_B|B|MID_SERIES 0  2e-13
RI2|_SPL_B|B|B I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SHUNT  2.7439617672
LI2|_SPL_B|B|RB I2|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_A|I_1|B I2|_DFF_A|A1 I2|_DFF_A|I_1|MID  2e-12
II2|_DFF_A|I_1|B 0 I2|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_3|B I2|_DFF_A|A3 I2|_DFF_A|I_3|MID  2e-12
II2|_DFF_A|I_3|B 0 I2|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_A|I_T|B I2|_DFF_A|T1 I2|_DFF_A|I_T|MID  2e-12
II2|_DFF_A|I_T|B 0 I2|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_6|B I2|_DFF_A|Q1 I2|_DFF_A|I_6|MID  2e-12
II2|_DFF_A|I_6|B 0 I2|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_A|1|1 I2|_DFF_A|A1 I2|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|1|P I2|_DFF_A|1|MID_SERIES 0  2e-13
RI2|_DFF_A|1|B I2|_DFF_A|A1 I2|_DFF_A|1|MID_SHUNT  2.7439617672
LI2|_DFF_A|1|RB I2|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|23|1 I2|_DFF_A|A2 I2|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|23|B I2|_DFF_A|A2 I2|_DFF_A|23|MID_SHUNT  3.84154647408
LI2|_DFF_A|23|RB I2|_DFF_A|23|MID_SHUNT I2|_DFF_A|A3  2.1704737578552e-12
BI2|_DFF_A|3|1 I2|_DFF_A|A3 I2|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|3|P I2|_DFF_A|3|MID_SERIES 0  2e-13
RI2|_DFF_A|3|B I2|_DFF_A|A3 I2|_DFF_A|3|MID_SHUNT  2.7439617672
LI2|_DFF_A|3|RB I2|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|4|1 I2|_DFF_A|A4 I2|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|4|P I2|_DFF_A|4|MID_SERIES 0  2e-13
RI2|_DFF_A|4|B I2|_DFF_A|A4 I2|_DFF_A|4|MID_SHUNT  2.7439617672
LI2|_DFF_A|4|RB I2|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|T|1 I2|_DFF_A|T1 I2|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|T|P I2|_DFF_A|T|MID_SERIES 0  2e-13
RI2|_DFF_A|T|B I2|_DFF_A|T1 I2|_DFF_A|T|MID_SHUNT  2.7439617672
LI2|_DFF_A|T|RB I2|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|45|1 I2|_DFF_A|T2 I2|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|45|B I2|_DFF_A|T2 I2|_DFF_A|45|MID_SHUNT  3.84154647408
LI2|_DFF_A|45|RB I2|_DFF_A|45|MID_SHUNT I2|_DFF_A|A4  2.1704737578552e-12
BI2|_DFF_A|6|1 I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|6|P I2|_DFF_A|6|MID_SERIES 0  2e-13
RI2|_DFF_A|6|B I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SHUNT  2.7439617672
LI2|_DFF_A|6|RB I2|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_B|I_1|B I2|_DFF_B|A1 I2|_DFF_B|I_1|MID  2e-12
II2|_DFF_B|I_1|B 0 I2|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_3|B I2|_DFF_B|A3 I2|_DFF_B|I_3|MID  2e-12
II2|_DFF_B|I_3|B 0 I2|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_B|I_T|B I2|_DFF_B|T1 I2|_DFF_B|I_T|MID  2e-12
II2|_DFF_B|I_T|B 0 I2|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_6|B I2|_DFF_B|Q1 I2|_DFF_B|I_6|MID  2e-12
II2|_DFF_B|I_6|B 0 I2|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_B|1|1 I2|_DFF_B|A1 I2|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|1|P I2|_DFF_B|1|MID_SERIES 0  2e-13
RI2|_DFF_B|1|B I2|_DFF_B|A1 I2|_DFF_B|1|MID_SHUNT  2.7439617672
LI2|_DFF_B|1|RB I2|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|23|1 I2|_DFF_B|A2 I2|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|23|B I2|_DFF_B|A2 I2|_DFF_B|23|MID_SHUNT  3.84154647408
LI2|_DFF_B|23|RB I2|_DFF_B|23|MID_SHUNT I2|_DFF_B|A3  2.1704737578552e-12
BI2|_DFF_B|3|1 I2|_DFF_B|A3 I2|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|3|P I2|_DFF_B|3|MID_SERIES 0  2e-13
RI2|_DFF_B|3|B I2|_DFF_B|A3 I2|_DFF_B|3|MID_SHUNT  2.7439617672
LI2|_DFF_B|3|RB I2|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|4|1 I2|_DFF_B|A4 I2|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|4|P I2|_DFF_B|4|MID_SERIES 0  2e-13
RI2|_DFF_B|4|B I2|_DFF_B|A4 I2|_DFF_B|4|MID_SHUNT  2.7439617672
LI2|_DFF_B|4|RB I2|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|T|1 I2|_DFF_B|T1 I2|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|T|P I2|_DFF_B|T|MID_SERIES 0  2e-13
RI2|_DFF_B|T|B I2|_DFF_B|T1 I2|_DFF_B|T|MID_SHUNT  2.7439617672
LI2|_DFF_B|T|RB I2|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|45|1 I2|_DFF_B|T2 I2|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|45|B I2|_DFF_B|T2 I2|_DFF_B|45|MID_SHUNT  3.84154647408
LI2|_DFF_B|45|RB I2|_DFF_B|45|MID_SHUNT I2|_DFF_B|A4  2.1704737578552e-12
BI2|_DFF_B|6|1 I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|6|P I2|_DFF_B|6|MID_SERIES 0  2e-13
RI2|_DFF_B|6|B I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SHUNT  2.7439617672
LI2|_DFF_B|6|RB I2|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI2|_XOR|I_A1|B I2|_XOR|A1 I2|_XOR|I_A1|MID  2e-12
II2|_XOR|I_A1|B 0 I2|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_A3|B I2|_XOR|A3 I2|_XOR|I_A3|MID  2e-12
II2|_XOR|I_A3|B 0 I2|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B1|B I2|_XOR|B1 I2|_XOR|I_B1|MID  2e-12
II2|_XOR|I_B1|B 0 I2|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B3|B I2|_XOR|B3 I2|_XOR|I_B3|MID  2e-12
II2|_XOR|I_B3|B 0 I2|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_Q1|B I2|_XOR|Q1 I2|_XOR|I_Q1|MID  2e-12
II2|_XOR|I_Q1|B 0 I2|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_XOR|A1|1 I2|_XOR|A1 I2|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A1|P I2|_XOR|A1|MID_SERIES 0  5e-13
RI2|_XOR|A1|B I2|_XOR|A1 I2|_XOR|A1|MID_SHUNT  2.7439617672
LI2|_XOR|A1|RB I2|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A2|1 I2|_XOR|A2 I2|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A2|P I2|_XOR|A2|MID_SERIES 0  5e-13
RI2|_XOR|A2|B I2|_XOR|A2 I2|_XOR|A2|MID_SHUNT  2.7439617672
LI2|_XOR|A2|RB I2|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A3|1 I2|_XOR|A2 I2|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A3|P I2|_XOR|A3|MID_SERIES I2|_XOR|A3  1.2e-12
RI2|_XOR|A3|B I2|_XOR|A2 I2|_XOR|A3|MID_SHUNT  2.7439617672
LI2|_XOR|A3|RB I2|_XOR|A3|MID_SHUNT I2|_XOR|A3  2.050338398468e-12
BI2|_XOR|B1|1 I2|_XOR|B1 I2|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B1|P I2|_XOR|B1|MID_SERIES 0  5e-13
RI2|_XOR|B1|B I2|_XOR|B1 I2|_XOR|B1|MID_SHUNT  2.7439617672
LI2|_XOR|B1|RB I2|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B2|1 I2|_XOR|B2 I2|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B2|P I2|_XOR|B2|MID_SERIES 0  5e-13
RI2|_XOR|B2|B I2|_XOR|B2 I2|_XOR|B2|MID_SHUNT  2.7439617672
LI2|_XOR|B2|RB I2|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B3|1 I2|_XOR|B2 I2|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B3|P I2|_XOR|B3|MID_SERIES I2|_XOR|B3  1.2e-12
RI2|_XOR|B3|B I2|_XOR|B2 I2|_XOR|B3|MID_SHUNT  2.7439617672
LI2|_XOR|B3|RB I2|_XOR|B3|MID_SHUNT I2|_XOR|B3  2.050338398468e-12
BI2|_XOR|T1|1 I2|_XOR|T1 I2|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|T1|P I2|_XOR|T1|MID_SERIES 0  5e-13
RI2|_XOR|T1|B I2|_XOR|T1 I2|_XOR|T1|MID_SHUNT  2.7439617672
LI2|_XOR|T1|RB I2|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|T2|1 I2|_XOR|T2 I2|_XOR|ABTQ JJMIT AREA=2.0
RI2|_XOR|T2|B I2|_XOR|T2 I2|_XOR|T2|MID_SHUNT  3.429952209
LI2|_XOR|T2|RB I2|_XOR|T2|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|AB|1 I2|_XOR|AB I2|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI2|_XOR|AB|P I2|_XOR|AB|MID_SERIES I2|_XOR|ABTQ  1.2e-12
RI2|_XOR|AB|B I2|_XOR|AB I2|_XOR|AB|MID_SHUNT  3.429952209
LI2|_XOR|AB|RB I2|_XOR|AB|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|ABTQ|1 I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|ABTQ|P I2|_XOR|ABTQ|MID_SERIES 0  5e-13
RI2|_XOR|ABTQ|B I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI2|_XOR|ABTQ|RB I2|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|Q1|1 I2|_XOR|Q1 I2|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|Q1|P I2|_XOR|Q1|MID_SERIES 0  5e-13
RI2|_XOR|Q1|B I2|_XOR|Q1 I2|_XOR|Q1|MID_SHUNT  2.7439617672
LI2|_XOR|Q1|RB I2|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI2|_AND|I_A1|B I2|_AND|A1 I2|_AND|I_A1|MID  2e-12
II2|_AND|I_A1|B 0 I2|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_B1|B I2|_AND|B1 I2|_AND|I_B1|MID  2e-12
II2|_AND|I_B1|B 0 I2|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q3|B I2|_AND|Q3 I2|_AND|I_Q3|MID  2e-12
II2|_AND|I_Q3|B 0 I2|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2|_AND|I_Q2|B I2|_AND|Q2 I2|_AND|I_Q2|MID  2e-12
II2|_AND|I_Q2|B 0 I2|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q1|B I2|_AND|Q1 I2|_AND|I_Q1|MID  2e-12
II2|_AND|I_Q1|B 0 I2|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_AND|A1|1 I2|_AND|A1 I2|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A1|P I2|_AND|A1|MID_SERIES 0  2e-13
RI2|_AND|A1|B I2|_AND|A1 I2|_AND|A1|MID_SHUNT  2.7439617672
LI2|_AND|A1|RB I2|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A2|1 I2|_AND|A2 I2|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A2|P I2|_AND|A2|MID_SERIES 0  2e-13
RI2|_AND|A2|B I2|_AND|A2 I2|_AND|A2|MID_SHUNT  2.7439617672
LI2|_AND|A2|RB I2|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A12|1 I2|_AND|A2 I2|_AND|A3 JJMIT AREA=1.7857142857142858
RI2|_AND|A12|B I2|_AND|A2 I2|_AND|A12|MID_SHUNT  3.84154647408
LI2|_AND|A12|RB I2|_AND|A12|MID_SHUNT I2|_AND|A3  2.1704737578552e-12
BI2|_AND|B1|1 I2|_AND|B1 I2|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B1|P I2|_AND|B1|MID_SERIES 0  2e-13
RI2|_AND|B1|B I2|_AND|B1 I2|_AND|B1|MID_SHUNT  2.7439617672
LI2|_AND|B1|RB I2|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B2|1 I2|_AND|B2 I2|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B2|P I2|_AND|B2|MID_SERIES 0  2e-13
RI2|_AND|B2|B I2|_AND|B2 I2|_AND|B2|MID_SHUNT  2.7439617672
LI2|_AND|B2|RB I2|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B12|1 I2|_AND|B2 I2|_AND|B3 JJMIT AREA=1.7857142857142858
RI2|_AND|B12|B I2|_AND|B2 I2|_AND|B12|MID_SHUNT  3.84154647408
LI2|_AND|B12|RB I2|_AND|B12|MID_SHUNT I2|_AND|B3  2.1704737578552e-12
BI2|_AND|Q2|1 I2|_AND|Q2 I2|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q2|P I2|_AND|Q2|MID_SERIES 0  2e-13
RI2|_AND|Q2|B I2|_AND|Q2 I2|_AND|Q2|MID_SHUNT  2.7439617672
LI2|_AND|Q2|RB I2|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|Q1|1 I2|_AND|Q1 I2|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q1|P I2|_AND|Q1|MID_SERIES 0  2e-13
RI2|_AND|Q1|B I2|_AND|Q1 I2|_AND|Q1|MID_SHUNT  2.7439617672
LI2|_AND|Q1|RB I2|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_A|I_D1|B I3|_SPL_A|D1 I3|_SPL_A|I_D1|MID  2e-12
II3|_SPL_A|I_D1|B 0 I3|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_D2|B I3|_SPL_A|D2 I3|_SPL_A|I_D2|MID  2e-12
II3|_SPL_A|I_D2|B 0 I3|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_A|I_Q1|B I3|_SPL_A|QA1 I3|_SPL_A|I_Q1|MID  2e-12
II3|_SPL_A|I_Q1|B 0 I3|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_Q2|B I3|_SPL_A|QB1 I3|_SPL_A|I_Q2|MID  2e-12
II3|_SPL_A|I_Q2|B 0 I3|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_A|1|1 I3|_SPL_A|D1 I3|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|1|P I3|_SPL_A|1|MID_SERIES 0  2e-13
RI3|_SPL_A|1|B I3|_SPL_A|D1 I3|_SPL_A|1|MID_SHUNT  2.7439617672
LI3|_SPL_A|1|RB I3|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|2|1 I3|_SPL_A|D2 I3|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|2|P I3|_SPL_A|2|MID_SERIES 0  2e-13
RI3|_SPL_A|2|B I3|_SPL_A|D2 I3|_SPL_A|2|MID_SHUNT  2.7439617672
LI3|_SPL_A|2|RB I3|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|A|1 I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|A|P I3|_SPL_A|A|MID_SERIES 0  2e-13
RI3|_SPL_A|A|B I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SHUNT  2.7439617672
LI3|_SPL_A|A|RB I3|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|B|1 I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|B|P I3|_SPL_A|B|MID_SERIES 0  2e-13
RI3|_SPL_A|B|B I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SHUNT  2.7439617672
LI3|_SPL_A|B|RB I3|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_B|I_D1|B I3|_SPL_B|D1 I3|_SPL_B|I_D1|MID  2e-12
II3|_SPL_B|I_D1|B 0 I3|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_D2|B I3|_SPL_B|D2 I3|_SPL_B|I_D2|MID  2e-12
II3|_SPL_B|I_D2|B 0 I3|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_B|I_Q1|B I3|_SPL_B|QA1 I3|_SPL_B|I_Q1|MID  2e-12
II3|_SPL_B|I_Q1|B 0 I3|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_Q2|B I3|_SPL_B|QB1 I3|_SPL_B|I_Q2|MID  2e-12
II3|_SPL_B|I_Q2|B 0 I3|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_B|1|1 I3|_SPL_B|D1 I3|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|1|P I3|_SPL_B|1|MID_SERIES 0  2e-13
RI3|_SPL_B|1|B I3|_SPL_B|D1 I3|_SPL_B|1|MID_SHUNT  2.7439617672
LI3|_SPL_B|1|RB I3|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|2|1 I3|_SPL_B|D2 I3|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|2|P I3|_SPL_B|2|MID_SERIES 0  2e-13
RI3|_SPL_B|2|B I3|_SPL_B|D2 I3|_SPL_B|2|MID_SHUNT  2.7439617672
LI3|_SPL_B|2|RB I3|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|A|1 I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|A|P I3|_SPL_B|A|MID_SERIES 0  2e-13
RI3|_SPL_B|A|B I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SHUNT  2.7439617672
LI3|_SPL_B|A|RB I3|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|B|1 I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|B|P I3|_SPL_B|B|MID_SERIES 0  2e-13
RI3|_SPL_B|B|B I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SHUNT  2.7439617672
LI3|_SPL_B|B|RB I3|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_A|I_1|B I3|_DFF_A|A1 I3|_DFF_A|I_1|MID  2e-12
II3|_DFF_A|I_1|B 0 I3|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_3|B I3|_DFF_A|A3 I3|_DFF_A|I_3|MID  2e-12
II3|_DFF_A|I_3|B 0 I3|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_A|I_T|B I3|_DFF_A|T1 I3|_DFF_A|I_T|MID  2e-12
II3|_DFF_A|I_T|B 0 I3|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_6|B I3|_DFF_A|Q1 I3|_DFF_A|I_6|MID  2e-12
II3|_DFF_A|I_6|B 0 I3|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_A|1|1 I3|_DFF_A|A1 I3|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|1|P I3|_DFF_A|1|MID_SERIES 0  2e-13
RI3|_DFF_A|1|B I3|_DFF_A|A1 I3|_DFF_A|1|MID_SHUNT  2.7439617672
LI3|_DFF_A|1|RB I3|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|23|1 I3|_DFF_A|A2 I3|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|23|B I3|_DFF_A|A2 I3|_DFF_A|23|MID_SHUNT  3.84154647408
LI3|_DFF_A|23|RB I3|_DFF_A|23|MID_SHUNT I3|_DFF_A|A3  2.1704737578552e-12
BI3|_DFF_A|3|1 I3|_DFF_A|A3 I3|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|3|P I3|_DFF_A|3|MID_SERIES 0  2e-13
RI3|_DFF_A|3|B I3|_DFF_A|A3 I3|_DFF_A|3|MID_SHUNT  2.7439617672
LI3|_DFF_A|3|RB I3|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|4|1 I3|_DFF_A|A4 I3|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|4|P I3|_DFF_A|4|MID_SERIES 0  2e-13
RI3|_DFF_A|4|B I3|_DFF_A|A4 I3|_DFF_A|4|MID_SHUNT  2.7439617672
LI3|_DFF_A|4|RB I3|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|T|1 I3|_DFF_A|T1 I3|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|T|P I3|_DFF_A|T|MID_SERIES 0  2e-13
RI3|_DFF_A|T|B I3|_DFF_A|T1 I3|_DFF_A|T|MID_SHUNT  2.7439617672
LI3|_DFF_A|T|RB I3|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|45|1 I3|_DFF_A|T2 I3|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|45|B I3|_DFF_A|T2 I3|_DFF_A|45|MID_SHUNT  3.84154647408
LI3|_DFF_A|45|RB I3|_DFF_A|45|MID_SHUNT I3|_DFF_A|A4  2.1704737578552e-12
BI3|_DFF_A|6|1 I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|6|P I3|_DFF_A|6|MID_SERIES 0  2e-13
RI3|_DFF_A|6|B I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SHUNT  2.7439617672
LI3|_DFF_A|6|RB I3|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_B|I_1|B I3|_DFF_B|A1 I3|_DFF_B|I_1|MID  2e-12
II3|_DFF_B|I_1|B 0 I3|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_3|B I3|_DFF_B|A3 I3|_DFF_B|I_3|MID  2e-12
II3|_DFF_B|I_3|B 0 I3|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_B|I_T|B I3|_DFF_B|T1 I3|_DFF_B|I_T|MID  2e-12
II3|_DFF_B|I_T|B 0 I3|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_6|B I3|_DFF_B|Q1 I3|_DFF_B|I_6|MID  2e-12
II3|_DFF_B|I_6|B 0 I3|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_B|1|1 I3|_DFF_B|A1 I3|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|1|P I3|_DFF_B|1|MID_SERIES 0  2e-13
RI3|_DFF_B|1|B I3|_DFF_B|A1 I3|_DFF_B|1|MID_SHUNT  2.7439617672
LI3|_DFF_B|1|RB I3|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|23|1 I3|_DFF_B|A2 I3|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|23|B I3|_DFF_B|A2 I3|_DFF_B|23|MID_SHUNT  3.84154647408
LI3|_DFF_B|23|RB I3|_DFF_B|23|MID_SHUNT I3|_DFF_B|A3  2.1704737578552e-12
BI3|_DFF_B|3|1 I3|_DFF_B|A3 I3|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|3|P I3|_DFF_B|3|MID_SERIES 0  2e-13
RI3|_DFF_B|3|B I3|_DFF_B|A3 I3|_DFF_B|3|MID_SHUNT  2.7439617672
LI3|_DFF_B|3|RB I3|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|4|1 I3|_DFF_B|A4 I3|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|4|P I3|_DFF_B|4|MID_SERIES 0  2e-13
RI3|_DFF_B|4|B I3|_DFF_B|A4 I3|_DFF_B|4|MID_SHUNT  2.7439617672
LI3|_DFF_B|4|RB I3|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|T|1 I3|_DFF_B|T1 I3|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|T|P I3|_DFF_B|T|MID_SERIES 0  2e-13
RI3|_DFF_B|T|B I3|_DFF_B|T1 I3|_DFF_B|T|MID_SHUNT  2.7439617672
LI3|_DFF_B|T|RB I3|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|45|1 I3|_DFF_B|T2 I3|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|45|B I3|_DFF_B|T2 I3|_DFF_B|45|MID_SHUNT  3.84154647408
LI3|_DFF_B|45|RB I3|_DFF_B|45|MID_SHUNT I3|_DFF_B|A4  2.1704737578552e-12
BI3|_DFF_B|6|1 I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|6|P I3|_DFF_B|6|MID_SERIES 0  2e-13
RI3|_DFF_B|6|B I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SHUNT  2.7439617672
LI3|_DFF_B|6|RB I3|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI3|_XOR|I_A1|B I3|_XOR|A1 I3|_XOR|I_A1|MID  2e-12
II3|_XOR|I_A1|B 0 I3|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_A3|B I3|_XOR|A3 I3|_XOR|I_A3|MID  2e-12
II3|_XOR|I_A3|B 0 I3|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B1|B I3|_XOR|B1 I3|_XOR|I_B1|MID  2e-12
II3|_XOR|I_B1|B 0 I3|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B3|B I3|_XOR|B3 I3|_XOR|I_B3|MID  2e-12
II3|_XOR|I_B3|B 0 I3|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_Q1|B I3|_XOR|Q1 I3|_XOR|I_Q1|MID  2e-12
II3|_XOR|I_Q1|B 0 I3|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_XOR|A1|1 I3|_XOR|A1 I3|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A1|P I3|_XOR|A1|MID_SERIES 0  5e-13
RI3|_XOR|A1|B I3|_XOR|A1 I3|_XOR|A1|MID_SHUNT  2.7439617672
LI3|_XOR|A1|RB I3|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A2|1 I3|_XOR|A2 I3|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A2|P I3|_XOR|A2|MID_SERIES 0  5e-13
RI3|_XOR|A2|B I3|_XOR|A2 I3|_XOR|A2|MID_SHUNT  2.7439617672
LI3|_XOR|A2|RB I3|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A3|1 I3|_XOR|A2 I3|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A3|P I3|_XOR|A3|MID_SERIES I3|_XOR|A3  1.2e-12
RI3|_XOR|A3|B I3|_XOR|A2 I3|_XOR|A3|MID_SHUNT  2.7439617672
LI3|_XOR|A3|RB I3|_XOR|A3|MID_SHUNT I3|_XOR|A3  2.050338398468e-12
BI3|_XOR|B1|1 I3|_XOR|B1 I3|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B1|P I3|_XOR|B1|MID_SERIES 0  5e-13
RI3|_XOR|B1|B I3|_XOR|B1 I3|_XOR|B1|MID_SHUNT  2.7439617672
LI3|_XOR|B1|RB I3|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B2|1 I3|_XOR|B2 I3|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B2|P I3|_XOR|B2|MID_SERIES 0  5e-13
RI3|_XOR|B2|B I3|_XOR|B2 I3|_XOR|B2|MID_SHUNT  2.7439617672
LI3|_XOR|B2|RB I3|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B3|1 I3|_XOR|B2 I3|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B3|P I3|_XOR|B3|MID_SERIES I3|_XOR|B3  1.2e-12
RI3|_XOR|B3|B I3|_XOR|B2 I3|_XOR|B3|MID_SHUNT  2.7439617672
LI3|_XOR|B3|RB I3|_XOR|B3|MID_SHUNT I3|_XOR|B3  2.050338398468e-12
BI3|_XOR|T1|1 I3|_XOR|T1 I3|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|T1|P I3|_XOR|T1|MID_SERIES 0  5e-13
RI3|_XOR|T1|B I3|_XOR|T1 I3|_XOR|T1|MID_SHUNT  2.7439617672
LI3|_XOR|T1|RB I3|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|T2|1 I3|_XOR|T2 I3|_XOR|ABTQ JJMIT AREA=2.0
RI3|_XOR|T2|B I3|_XOR|T2 I3|_XOR|T2|MID_SHUNT  3.429952209
LI3|_XOR|T2|RB I3|_XOR|T2|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|AB|1 I3|_XOR|AB I3|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI3|_XOR|AB|P I3|_XOR|AB|MID_SERIES I3|_XOR|ABTQ  1.2e-12
RI3|_XOR|AB|B I3|_XOR|AB I3|_XOR|AB|MID_SHUNT  3.429952209
LI3|_XOR|AB|RB I3|_XOR|AB|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|ABTQ|1 I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|ABTQ|P I3|_XOR|ABTQ|MID_SERIES 0  5e-13
RI3|_XOR|ABTQ|B I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI3|_XOR|ABTQ|RB I3|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|Q1|1 I3|_XOR|Q1 I3|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|Q1|P I3|_XOR|Q1|MID_SERIES 0  5e-13
RI3|_XOR|Q1|B I3|_XOR|Q1 I3|_XOR|Q1|MID_SHUNT  2.7439617672
LI3|_XOR|Q1|RB I3|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI3|_AND|I_A1|B I3|_AND|A1 I3|_AND|I_A1|MID  2e-12
II3|_AND|I_A1|B 0 I3|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_B1|B I3|_AND|B1 I3|_AND|I_B1|MID  2e-12
II3|_AND|I_B1|B 0 I3|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q3|B I3|_AND|Q3 I3|_AND|I_Q3|MID  2e-12
II3|_AND|I_Q3|B 0 I3|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3|_AND|I_Q2|B I3|_AND|Q2 I3|_AND|I_Q2|MID  2e-12
II3|_AND|I_Q2|B 0 I3|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q1|B I3|_AND|Q1 I3|_AND|I_Q1|MID  2e-12
II3|_AND|I_Q1|B 0 I3|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_AND|A1|1 I3|_AND|A1 I3|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A1|P I3|_AND|A1|MID_SERIES 0  2e-13
RI3|_AND|A1|B I3|_AND|A1 I3|_AND|A1|MID_SHUNT  2.7439617672
LI3|_AND|A1|RB I3|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A2|1 I3|_AND|A2 I3|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A2|P I3|_AND|A2|MID_SERIES 0  2e-13
RI3|_AND|A2|B I3|_AND|A2 I3|_AND|A2|MID_SHUNT  2.7439617672
LI3|_AND|A2|RB I3|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A12|1 I3|_AND|A2 I3|_AND|A3 JJMIT AREA=1.7857142857142858
RI3|_AND|A12|B I3|_AND|A2 I3|_AND|A12|MID_SHUNT  3.84154647408
LI3|_AND|A12|RB I3|_AND|A12|MID_SHUNT I3|_AND|A3  2.1704737578552e-12
BI3|_AND|B1|1 I3|_AND|B1 I3|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B1|P I3|_AND|B1|MID_SERIES 0  2e-13
RI3|_AND|B1|B I3|_AND|B1 I3|_AND|B1|MID_SHUNT  2.7439617672
LI3|_AND|B1|RB I3|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B2|1 I3|_AND|B2 I3|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B2|P I3|_AND|B2|MID_SERIES 0  2e-13
RI3|_AND|B2|B I3|_AND|B2 I3|_AND|B2|MID_SHUNT  2.7439617672
LI3|_AND|B2|RB I3|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B12|1 I3|_AND|B2 I3|_AND|B3 JJMIT AREA=1.7857142857142858
RI3|_AND|B12|B I3|_AND|B2 I3|_AND|B12|MID_SHUNT  3.84154647408
LI3|_AND|B12|RB I3|_AND|B12|MID_SHUNT I3|_AND|B3  2.1704737578552e-12
BI3|_AND|Q2|1 I3|_AND|Q2 I3|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q2|P I3|_AND|Q2|MID_SERIES 0  2e-13
RI3|_AND|Q2|B I3|_AND|Q2 I3|_AND|Q2|MID_SHUNT  2.7439617672
LI3|_AND|Q2|RB I3|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|Q1|1 I3|_AND|Q1 I3|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q1|P I3|_AND|Q1|MID_SERIES 0  2e-13
RI3|_AND|Q1|B I3|_AND|Q1 I3|_AND|Q1|MID_SHUNT  2.7439617672
LI3|_AND|Q1|RB I3|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|I_D1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|I_D1|MID  2e-12
ISPL_IP2_0|SPL1|I_D1|B 0 SPL_IP2_0|SPL1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP2_0|SPL1|I_D2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|I_D2|MID  2e-12
ISPL_IP2_0|SPL1|I_D2|B 0 SPL_IP2_0|SPL1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP2_0|SPL1|I_Q1|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|I_Q1|MID  2e-12
ISPL_IP2_0|SPL1|I_Q1|B 0 SPL_IP2_0|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP2_0|SPL1|I_Q2|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|I_Q2|MID  2e-12
ISPL_IP2_0|SPL1|I_Q2|B 0 SPL_IP2_0|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP2_0|SPL1|1|1 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|1|P SPL_IP2_0|SPL1|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|1|RB SPL_IP2_0|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|2|1 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|2|P SPL_IP2_0|SPL1|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|2|RB SPL_IP2_0|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|A|1 SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|A|P SPL_IP2_0|SPL1|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|A|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|A|RB SPL_IP2_0|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|B|1 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|B|P SPL_IP2_0|SPL1|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|B|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|B|RB SPL_IP2_0|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL2|I_D1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|I_D1|MID  2e-12
ISPL_IP2_0|SPL2|I_D1|B 0 SPL_IP2_0|SPL2|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP2_0|SPL2|I_D2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|I_D2|MID  2e-12
ISPL_IP2_0|SPL2|I_D2|B 0 SPL_IP2_0|SPL2|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP2_0|SPL2|I_Q1|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|I_Q1|MID  2e-12
ISPL_IP2_0|SPL2|I_Q1|B 0 SPL_IP2_0|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP2_0|SPL2|I_Q2|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|I_Q2|MID  2e-12
ISPL_IP2_0|SPL2|I_Q2|B 0 SPL_IP2_0|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP2_0|SPL2|1|1 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|1|P SPL_IP2_0|SPL2|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|1|RB SPL_IP2_0|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|2|1 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|2|P SPL_IP2_0|SPL2|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|2|RB SPL_IP2_0|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|A|1 SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|A|P SPL_IP2_0|SPL2|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|A|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|A|RB SPL_IP2_0|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|B|1 SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|B|P SPL_IP2_0|SPL2|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|B|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|B|RB SPL_IP2_0|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|I_1|B _PG0_01|P|A1 _PG0_01|P|I_1|MID  2e-12
I_PG0_01|P|I_1|B 0 _PG0_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_3|B _PG0_01|P|A3 _PG0_01|P|I_3|MID  2e-12
I_PG0_01|P|I_3|B 0 _PG0_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|P|I_T|B _PG0_01|P|T1 _PG0_01|P|I_T|MID  2e-12
I_PG0_01|P|I_T|B 0 _PG0_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_6|B _PG0_01|P|Q1 _PG0_01|P|I_6|MID  2e-12
I_PG0_01|P|I_6|B 0 _PG0_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|P|1|1 _PG0_01|P|A1 _PG0_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|1|P _PG0_01|P|1|MID_SERIES 0  2e-13
R_PG0_01|P|1|B _PG0_01|P|A1 _PG0_01|P|1|MID_SHUNT  2.7439617672
L_PG0_01|P|1|RB _PG0_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|23|1 _PG0_01|P|A2 _PG0_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|P|23|B _PG0_01|P|A2 _PG0_01|P|23|MID_SHUNT  3.84154647408
L_PG0_01|P|23|RB _PG0_01|P|23|MID_SHUNT _PG0_01|P|A3  2.1704737578552e-12
B_PG0_01|P|3|1 _PG0_01|P|A3 _PG0_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|3|P _PG0_01|P|3|MID_SERIES 0  2e-13
R_PG0_01|P|3|B _PG0_01|P|A3 _PG0_01|P|3|MID_SHUNT  2.7439617672
L_PG0_01|P|3|RB _PG0_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|4|1 _PG0_01|P|A4 _PG0_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|4|P _PG0_01|P|4|MID_SERIES 0  2e-13
R_PG0_01|P|4|B _PG0_01|P|A4 _PG0_01|P|4|MID_SHUNT  2.7439617672
L_PG0_01|P|4|RB _PG0_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|T|1 _PG0_01|P|T1 _PG0_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|T|P _PG0_01|P|T|MID_SERIES 0  2e-13
R_PG0_01|P|T|B _PG0_01|P|T1 _PG0_01|P|T|MID_SHUNT  2.7439617672
L_PG0_01|P|T|RB _PG0_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|45|1 _PG0_01|P|T2 _PG0_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|P|45|B _PG0_01|P|T2 _PG0_01|P|45|MID_SHUNT  3.84154647408
L_PG0_01|P|45|RB _PG0_01|P|45|MID_SHUNT _PG0_01|P|A4  2.1704737578552e-12
B_PG0_01|P|6|1 _PG0_01|P|Q1 _PG0_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|6|P _PG0_01|P|6|MID_SERIES 0  2e-13
R_PG0_01|P|6|B _PG0_01|P|Q1 _PG0_01|P|6|MID_SHUNT  2.7439617672
L_PG0_01|P|6|RB _PG0_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|G|I_1|B _PG0_01|G|A1 _PG0_01|G|I_1|MID  2e-12
I_PG0_01|G|I_1|B 0 _PG0_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_3|B _PG0_01|G|A3 _PG0_01|G|I_3|MID  2e-12
I_PG0_01|G|I_3|B 0 _PG0_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|G|I_T|B _PG0_01|G|T1 _PG0_01|G|I_T|MID  2e-12
I_PG0_01|G|I_T|B 0 _PG0_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_6|B _PG0_01|G|Q1 _PG0_01|G|I_6|MID  2e-12
I_PG0_01|G|I_6|B 0 _PG0_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|G|1|1 _PG0_01|G|A1 _PG0_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|1|P _PG0_01|G|1|MID_SERIES 0  2e-13
R_PG0_01|G|1|B _PG0_01|G|A1 _PG0_01|G|1|MID_SHUNT  2.7439617672
L_PG0_01|G|1|RB _PG0_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|23|1 _PG0_01|G|A2 _PG0_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|G|23|B _PG0_01|G|A2 _PG0_01|G|23|MID_SHUNT  3.84154647408
L_PG0_01|G|23|RB _PG0_01|G|23|MID_SHUNT _PG0_01|G|A3  2.1704737578552e-12
B_PG0_01|G|3|1 _PG0_01|G|A3 _PG0_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|3|P _PG0_01|G|3|MID_SERIES 0  2e-13
R_PG0_01|G|3|B _PG0_01|G|A3 _PG0_01|G|3|MID_SHUNT  2.7439617672
L_PG0_01|G|3|RB _PG0_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|4|1 _PG0_01|G|A4 _PG0_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|4|P _PG0_01|G|4|MID_SERIES 0  2e-13
R_PG0_01|G|4|B _PG0_01|G|A4 _PG0_01|G|4|MID_SHUNT  2.7439617672
L_PG0_01|G|4|RB _PG0_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|T|1 _PG0_01|G|T1 _PG0_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|T|P _PG0_01|G|T|MID_SERIES 0  2e-13
R_PG0_01|G|T|B _PG0_01|G|T1 _PG0_01|G|T|MID_SHUNT  2.7439617672
L_PG0_01|G|T|RB _PG0_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|45|1 _PG0_01|G|T2 _PG0_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|G|45|B _PG0_01|G|T2 _PG0_01|G|45|MID_SHUNT  3.84154647408
L_PG0_01|G|45|RB _PG0_01|G|45|MID_SHUNT _PG0_01|G|A4  2.1704737578552e-12
B_PG0_01|G|6|1 _PG0_01|G|Q1 _PG0_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|6|P _PG0_01|G|6|MID_SERIES 0  2e-13
R_PG0_01|G|6|B _PG0_01|G|Q1 _PG0_01|G|6|MID_SHUNT  2.7439617672
L_PG0_01|G|6|RB _PG0_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_SPL_G1|I_D1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|I_D1|MID  2e-12
I_PG1_01|_SPL_G1|I_D1|B 0 _PG1_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_D2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|I_D2|MID  2e-12
I_PG1_01|_SPL_G1|I_D2|B 0 _PG1_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG1_01|_SPL_G1|I_Q1|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|I_Q1|MID  2e-12
I_PG1_01|_SPL_G1|I_Q1|B 0 _PG1_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_Q2|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|I_Q2|MID  2e-12
I_PG1_01|_SPL_G1|I_Q2|B 0 _PG1_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG1_01|_SPL_G1|1|1 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|1|P _PG1_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|1|RB _PG1_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|2|1 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|2|P _PG1_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|2|RB _PG1_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|A|1 _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|A|P _PG1_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|A|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|A|RB _PG1_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|B|1 _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|B|P _PG1_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|B|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|B|RB _PG1_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_PG|I_A1|B _PG1_01|_PG|A1 _PG1_01|_PG|I_A1|MID  2e-12
I_PG1_01|_PG|I_A1|B 0 _PG1_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_B1|B _PG1_01|_PG|B1 _PG1_01|_PG|I_B1|MID  2e-12
I_PG1_01|_PG|I_B1|B 0 _PG1_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q3|B _PG1_01|_PG|Q3 _PG1_01|_PG|I_Q3|MID  2e-12
I_PG1_01|_PG|I_Q3|B 0 _PG1_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_PG|I_Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|I_Q2|MID  2e-12
I_PG1_01|_PG|I_Q2|B 0 _PG1_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|I_Q1|MID  2e-12
I_PG1_01|_PG|I_Q1|B 0 _PG1_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_PG|A1|1 _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A1|P _PG1_01|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01|_PG|A1|B _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A1|RB _PG1_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A2|1 _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A2|P _PG1_01|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01|_PG|A2|B _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A2|RB _PG1_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A12|1 _PG1_01|_PG|A2 _PG1_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|A12|B _PG1_01|_PG|A2 _PG1_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|A12|RB _PG1_01|_PG|A12|MID_SHUNT _PG1_01|_PG|A3  2.1704737578552e-12
B_PG1_01|_PG|B1|1 _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B1|P _PG1_01|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01|_PG|B1|B _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B1|RB _PG1_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B2|1 _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B2|P _PG1_01|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01|_PG|B2|B _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B2|RB _PG1_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B12|1 _PG1_01|_PG|B2 _PG1_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|B12|B _PG1_01|_PG|B2 _PG1_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|B12|RB _PG1_01|_PG|B12|MID_SHUNT _PG1_01|_PG|B3  2.1704737578552e-12
B_PG1_01|_PG|Q2|1 _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q2|P _PG1_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q2|RB _PG1_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|Q1|1 _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q1|P _PG1_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q1|RB _PG1_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_GG|I_A1|B _PG1_01|_GG|A1 _PG1_01|_GG|I_A1|MID  2e-12
I_PG1_01|_GG|I_A1|B 0 _PG1_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_B1|B _PG1_01|_GG|B1 _PG1_01|_GG|I_B1|MID  2e-12
I_PG1_01|_GG|I_B1|B 0 _PG1_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q3|B _PG1_01|_GG|Q3 _PG1_01|_GG|I_Q3|MID  2e-12
I_PG1_01|_GG|I_Q3|B 0 _PG1_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_GG|I_Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|I_Q2|MID  2e-12
I_PG1_01|_GG|I_Q2|B 0 _PG1_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|I_Q1|MID  2e-12
I_PG1_01|_GG|I_Q1|B 0 _PG1_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_GG|A1|1 _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A1|P _PG1_01|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01|_GG|A1|B _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A1|RB _PG1_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A2|1 _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A2|P _PG1_01|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01|_GG|A2|B _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A2|RB _PG1_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A12|1 _PG1_01|_GG|A2 _PG1_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|A12|B _PG1_01|_GG|A2 _PG1_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|A12|RB _PG1_01|_GG|A12|MID_SHUNT _PG1_01|_GG|A3  2.1704737578552e-12
B_PG1_01|_GG|B1|1 _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B1|P _PG1_01|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01|_GG|B1|B _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B1|RB _PG1_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B2|1 _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B2|P _PG1_01|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01|_GG|B2|B _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B2|RB _PG1_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B12|1 _PG1_01|_GG|B2 _PG1_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|B12|B _PG1_01|_GG|B2 _PG1_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|B12|RB _PG1_01|_GG|B12|MID_SHUNT _PG1_01|_GG|B3  2.1704737578552e-12
B_PG1_01|_GG|Q2|1 _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q2|P _PG1_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q2|RB _PG1_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|Q1|1 _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q1|P _PG1_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q1|RB _PG1_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_PG|I_1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|I_1|MID  2e-12
I_PG1_01|_DFF_PG|I_1|B 0 _PG1_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|I_3|MID  2e-12
I_PG1_01|_DFF_PG|I_3|B 0 _PG1_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_PG|I_T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|I_T|MID  2e-12
I_PG1_01|_DFF_PG|I_T|B 0 _PG1_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|I_6|MID  2e-12
I_PG1_01|_DFF_PG|I_6|B 0 _PG1_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_PG|1|1 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|1|P _PG1_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|1|RB _PG1_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|23|1 _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|23|B _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|23|RB _PG1_01|_DFF_PG|23|MID_SHUNT _PG1_01|_DFF_PG|A3  2.1704737578552e-12
B_PG1_01|_DFF_PG|3|1 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|3|P _PG1_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|3|RB _PG1_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|4|1 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|4|P _PG1_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|4|B _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|4|RB _PG1_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|T|1 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|T|P _PG1_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|T|RB _PG1_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|45|1 _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|45|B _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|45|RB _PG1_01|_DFF_PG|45|MID_SHUNT _PG1_01|_DFF_PG|A4  2.1704737578552e-12
B_PG1_01|_DFF_PG|6|1 _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|6|P _PG1_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|6|RB _PG1_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_GG|I_1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|I_1|MID  2e-12
I_PG1_01|_DFF_GG|I_1|B 0 _PG1_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|I_3|MID  2e-12
I_PG1_01|_DFF_GG|I_3|B 0 _PG1_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_GG|I_T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|I_T|MID  2e-12
I_PG1_01|_DFF_GG|I_T|B 0 _PG1_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|I_6|MID  2e-12
I_PG1_01|_DFF_GG|I_6|B 0 _PG1_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_GG|1|1 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|1|P _PG1_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|1|RB _PG1_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|23|1 _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|23|B _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|23|RB _PG1_01|_DFF_GG|23|MID_SHUNT _PG1_01|_DFF_GG|A3  2.1704737578552e-12
B_PG1_01|_DFF_GG|3|1 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|3|P _PG1_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|3|RB _PG1_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|4|1 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|4|P _PG1_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|4|B _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|4|RB _PG1_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|T|1 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|T|P _PG1_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|T|RB _PG1_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|45|1 _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|45|B _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|45|RB _PG1_01|_DFF_GG|45|MID_SHUNT _PG1_01|_DFF_GG|A4  2.1704737578552e-12
B_PG1_01|_DFF_GG|6|1 _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|6|P _PG1_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|6|RB _PG1_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_G|I_A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|I_A1|MID  2e-12
I_PG1_01|_AND_G|I_A1|B 0 _PG1_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|I_B1|MID  2e-12
I_PG1_01|_AND_G|I_B1|B 0 _PG1_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q3|B _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|I_Q3|MID  2e-12
I_PG1_01|_AND_G|I_Q3|B 0 _PG1_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_G|I_Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|I_Q2|MID  2e-12
I_PG1_01|_AND_G|I_Q2|B 0 _PG1_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|I_Q1|MID  2e-12
I_PG1_01|_AND_G|I_Q1|B 0 _PG1_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_G|A1|1 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A1|P _PG1_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A1|RB _PG1_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A2|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A2|P _PG1_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A2|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A2|RB _PG1_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A12|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|A12|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|A12|RB _PG1_01|_AND_G|A12|MID_SHUNT _PG1_01|_AND_G|A3  2.1704737578552e-12
B_PG1_01|_AND_G|B1|1 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B1|P _PG1_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B1|RB _PG1_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B2|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B2|P _PG1_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B2|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B2|RB _PG1_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B12|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|B12|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|B12|RB _PG1_01|_AND_G|B12|MID_SHUNT _PG1_01|_AND_G|B3  2.1704737578552e-12
B_PG1_01|_AND_G|Q2|1 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q2|P _PG1_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q2|RB _PG1_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|Q1|1 _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q1|P _PG1_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q1|RB _PG1_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|P|I_1|B _PG2_01|P|A1 _PG2_01|P|I_1|MID  2e-12
I_PG2_01|P|I_1|B 0 _PG2_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_3|B _PG2_01|P|A3 _PG2_01|P|I_3|MID  2e-12
I_PG2_01|P|I_3|B 0 _PG2_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|P|I_T|B _PG2_01|P|T1 _PG2_01|P|I_T|MID  2e-12
I_PG2_01|P|I_T|B 0 _PG2_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_6|B _PG2_01|P|Q1 _PG2_01|P|I_6|MID  2e-12
I_PG2_01|P|I_6|B 0 _PG2_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|P|1|1 _PG2_01|P|A1 _PG2_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|1|P _PG2_01|P|1|MID_SERIES 0  2e-13
R_PG2_01|P|1|B _PG2_01|P|A1 _PG2_01|P|1|MID_SHUNT  2.7439617672
L_PG2_01|P|1|RB _PG2_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|23|1 _PG2_01|P|A2 _PG2_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|P|23|B _PG2_01|P|A2 _PG2_01|P|23|MID_SHUNT  3.84154647408
L_PG2_01|P|23|RB _PG2_01|P|23|MID_SHUNT _PG2_01|P|A3  2.1704737578552e-12
B_PG2_01|P|3|1 _PG2_01|P|A3 _PG2_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|3|P _PG2_01|P|3|MID_SERIES 0  2e-13
R_PG2_01|P|3|B _PG2_01|P|A3 _PG2_01|P|3|MID_SHUNT  2.7439617672
L_PG2_01|P|3|RB _PG2_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|4|1 _PG2_01|P|A4 _PG2_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|4|P _PG2_01|P|4|MID_SERIES 0  2e-13
R_PG2_01|P|4|B _PG2_01|P|A4 _PG2_01|P|4|MID_SHUNT  2.7439617672
L_PG2_01|P|4|RB _PG2_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|T|1 _PG2_01|P|T1 _PG2_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|T|P _PG2_01|P|T|MID_SERIES 0  2e-13
R_PG2_01|P|T|B _PG2_01|P|T1 _PG2_01|P|T|MID_SHUNT  2.7439617672
L_PG2_01|P|T|RB _PG2_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|45|1 _PG2_01|P|T2 _PG2_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|P|45|B _PG2_01|P|T2 _PG2_01|P|45|MID_SHUNT  3.84154647408
L_PG2_01|P|45|RB _PG2_01|P|45|MID_SHUNT _PG2_01|P|A4  2.1704737578552e-12
B_PG2_01|P|6|1 _PG2_01|P|Q1 _PG2_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|6|P _PG2_01|P|6|MID_SERIES 0  2e-13
R_PG2_01|P|6|B _PG2_01|P|Q1 _PG2_01|P|6|MID_SHUNT  2.7439617672
L_PG2_01|P|6|RB _PG2_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|G|I_1|B _PG2_01|G|A1 _PG2_01|G|I_1|MID  2e-12
I_PG2_01|G|I_1|B 0 _PG2_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_3|B _PG2_01|G|A3 _PG2_01|G|I_3|MID  2e-12
I_PG2_01|G|I_3|B 0 _PG2_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|G|I_T|B _PG2_01|G|T1 _PG2_01|G|I_T|MID  2e-12
I_PG2_01|G|I_T|B 0 _PG2_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_6|B _PG2_01|G|Q1 _PG2_01|G|I_6|MID  2e-12
I_PG2_01|G|I_6|B 0 _PG2_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|G|1|1 _PG2_01|G|A1 _PG2_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|1|P _PG2_01|G|1|MID_SERIES 0  2e-13
R_PG2_01|G|1|B _PG2_01|G|A1 _PG2_01|G|1|MID_SHUNT  2.7439617672
L_PG2_01|G|1|RB _PG2_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|23|1 _PG2_01|G|A2 _PG2_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|G|23|B _PG2_01|G|A2 _PG2_01|G|23|MID_SHUNT  3.84154647408
L_PG2_01|G|23|RB _PG2_01|G|23|MID_SHUNT _PG2_01|G|A3  2.1704737578552e-12
B_PG2_01|G|3|1 _PG2_01|G|A3 _PG2_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|3|P _PG2_01|G|3|MID_SERIES 0  2e-13
R_PG2_01|G|3|B _PG2_01|G|A3 _PG2_01|G|3|MID_SHUNT  2.7439617672
L_PG2_01|G|3|RB _PG2_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|4|1 _PG2_01|G|A4 _PG2_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|4|P _PG2_01|G|4|MID_SERIES 0  2e-13
R_PG2_01|G|4|B _PG2_01|G|A4 _PG2_01|G|4|MID_SHUNT  2.7439617672
L_PG2_01|G|4|RB _PG2_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|T|1 _PG2_01|G|T1 _PG2_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|T|P _PG2_01|G|T|MID_SERIES 0  2e-13
R_PG2_01|G|T|B _PG2_01|G|T1 _PG2_01|G|T|MID_SHUNT  2.7439617672
L_PG2_01|G|T|RB _PG2_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|45|1 _PG2_01|G|T2 _PG2_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|G|45|B _PG2_01|G|T2 _PG2_01|G|45|MID_SHUNT  3.84154647408
L_PG2_01|G|45|RB _PG2_01|G|45|MID_SHUNT _PG2_01|G|A4  2.1704737578552e-12
B_PG2_01|G|6|1 _PG2_01|G|Q1 _PG2_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|6|P _PG2_01|G|6|MID_SERIES 0  2e-13
R_PG2_01|G|6|B _PG2_01|G|Q1 _PG2_01|G|6|MID_SHUNT  2.7439617672
L_PG2_01|G|6|RB _PG2_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_G1|I_D1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|I_D1|MID  2e-12
I_PG3_01|_SPL_G1|I_D1|B 0 _PG3_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_D2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|I_D2|MID  2e-12
I_PG3_01|_SPL_G1|I_D2|B 0 _PG3_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_G1|I_Q1|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|I_Q1|MID  2e-12
I_PG3_01|_SPL_G1|I_Q1|B 0 _PG3_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_Q2|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|I_Q2|MID  2e-12
I_PG3_01|_SPL_G1|I_Q2|B 0 _PG3_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_G1|1|1 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|1|P _PG3_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|1|RB _PG3_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|2|1 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|2|P _PG3_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|2|RB _PG3_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|A|1 _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|A|P _PG3_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|A|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|A|RB _PG3_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|B|1 _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|B|P _PG3_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|B|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|B|RB _PG3_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_P1|I_D1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|I_D1|MID  2e-12
I_PG3_01|_SPL_P1|I_D1|B 0 _PG3_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_D2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|I_D2|MID  2e-12
I_PG3_01|_SPL_P1|I_D2|B 0 _PG3_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_P1|I_Q1|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|I_Q1|MID  2e-12
I_PG3_01|_SPL_P1|I_Q1|B 0 _PG3_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_Q2|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|I_Q2|MID  2e-12
I_PG3_01|_SPL_P1|I_Q2|B 0 _PG3_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_P1|1|1 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|1|P _PG3_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|1|RB _PG3_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|2|1 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|2|P _PG3_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|2|RB _PG3_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|A|1 _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|A|P _PG3_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|A|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|A|RB _PG3_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|B|1 _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|B|P _PG3_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|B|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|B|RB _PG3_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_PG|I_A1|B _PG3_01|_PG|A1 _PG3_01|_PG|I_A1|MID  2e-12
I_PG3_01|_PG|I_A1|B 0 _PG3_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_B1|B _PG3_01|_PG|B1 _PG3_01|_PG|I_B1|MID  2e-12
I_PG3_01|_PG|I_B1|B 0 _PG3_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q3|B _PG3_01|_PG|Q3 _PG3_01|_PG|I_Q3|MID  2e-12
I_PG3_01|_PG|I_Q3|B 0 _PG3_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_PG|I_Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|I_Q2|MID  2e-12
I_PG3_01|_PG|I_Q2|B 0 _PG3_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|I_Q1|MID  2e-12
I_PG3_01|_PG|I_Q1|B 0 _PG3_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_PG|A1|1 _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A1|P _PG3_01|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01|_PG|A1|B _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A1|RB _PG3_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A2|1 _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A2|P _PG3_01|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01|_PG|A2|B _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A2|RB _PG3_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A12|1 _PG3_01|_PG|A2 _PG3_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|A12|B _PG3_01|_PG|A2 _PG3_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|A12|RB _PG3_01|_PG|A12|MID_SHUNT _PG3_01|_PG|A3  2.1704737578552e-12
B_PG3_01|_PG|B1|1 _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B1|P _PG3_01|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01|_PG|B1|B _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B1|RB _PG3_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B2|1 _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B2|P _PG3_01|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01|_PG|B2|B _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B2|RB _PG3_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B12|1 _PG3_01|_PG|B2 _PG3_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|B12|B _PG3_01|_PG|B2 _PG3_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|B12|RB _PG3_01|_PG|B12|MID_SHUNT _PG3_01|_PG|B3  2.1704737578552e-12
B_PG3_01|_PG|Q2|1 _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q2|P _PG3_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q2|RB _PG3_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|Q1|1 _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q1|P _PG3_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q1|RB _PG3_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_GG|I_A1|B _PG3_01|_GG|A1 _PG3_01|_GG|I_A1|MID  2e-12
I_PG3_01|_GG|I_A1|B 0 _PG3_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_B1|B _PG3_01|_GG|B1 _PG3_01|_GG|I_B1|MID  2e-12
I_PG3_01|_GG|I_B1|B 0 _PG3_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q3|B _PG3_01|_GG|Q3 _PG3_01|_GG|I_Q3|MID  2e-12
I_PG3_01|_GG|I_Q3|B 0 _PG3_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_GG|I_Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|I_Q2|MID  2e-12
I_PG3_01|_GG|I_Q2|B 0 _PG3_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|I_Q1|MID  2e-12
I_PG3_01|_GG|I_Q1|B 0 _PG3_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_GG|A1|1 _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A1|P _PG3_01|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01|_GG|A1|B _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A1|RB _PG3_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A2|1 _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A2|P _PG3_01|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01|_GG|A2|B _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A2|RB _PG3_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A12|1 _PG3_01|_GG|A2 _PG3_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|A12|B _PG3_01|_GG|A2 _PG3_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|A12|RB _PG3_01|_GG|A12|MID_SHUNT _PG3_01|_GG|A3  2.1704737578552e-12
B_PG3_01|_GG|B1|1 _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B1|P _PG3_01|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01|_GG|B1|B _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B1|RB _PG3_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B2|1 _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B2|P _PG3_01|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01|_GG|B2|B _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B2|RB _PG3_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B12|1 _PG3_01|_GG|B2 _PG3_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|B12|B _PG3_01|_GG|B2 _PG3_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|B12|RB _PG3_01|_GG|B12|MID_SHUNT _PG3_01|_GG|B3  2.1704737578552e-12
B_PG3_01|_GG|Q2|1 _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q2|P _PG3_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q2|RB _PG3_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|Q1|1 _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q1|P _PG3_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q1|RB _PG3_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P0|I_1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|I_1|MID  2e-12
I_PG3_01|_DFF_P0|I_1|B 0 _PG3_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|I_3|MID  2e-12
I_PG3_01|_DFF_P0|I_3|B 0 _PG3_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P0|I_T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|I_T|MID  2e-12
I_PG3_01|_DFF_P0|I_T|B 0 _PG3_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|I_6|MID  2e-12
I_PG3_01|_DFF_P0|I_6|B 0 _PG3_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P0|1|1 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|1|P _PG3_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|1|RB _PG3_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|23|1 _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|23|B _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|23|RB _PG3_01|_DFF_P0|23|MID_SHUNT _PG3_01|_DFF_P0|A3  2.1704737578552e-12
B_PG3_01|_DFF_P0|3|1 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|3|P _PG3_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|3|RB _PG3_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|4|1 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|4|P _PG3_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|4|B _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|4|RB _PG3_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|T|1 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|T|P _PG3_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|T|RB _PG3_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|45|1 _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|45|B _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|45|RB _PG3_01|_DFF_P0|45|MID_SHUNT _PG3_01|_DFF_P0|A4  2.1704737578552e-12
B_PG3_01|_DFF_P0|6|1 _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|6|P _PG3_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|6|RB _PG3_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P1|I_1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|I_1|MID  2e-12
I_PG3_01|_DFF_P1|I_1|B 0 _PG3_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|I_3|MID  2e-12
I_PG3_01|_DFF_P1|I_3|B 0 _PG3_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P1|I_T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|I_T|MID  2e-12
I_PG3_01|_DFF_P1|I_T|B 0 _PG3_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|I_6|MID  2e-12
I_PG3_01|_DFF_P1|I_6|B 0 _PG3_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P1|1|1 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|1|P _PG3_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|1|RB _PG3_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|23|1 _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|23|B _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|23|RB _PG3_01|_DFF_P1|23|MID_SHUNT _PG3_01|_DFF_P1|A3  2.1704737578552e-12
B_PG3_01|_DFF_P1|3|1 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|3|P _PG3_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|3|RB _PG3_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|4|1 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|4|P _PG3_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|4|B _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|4|RB _PG3_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|T|1 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|T|P _PG3_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|T|RB _PG3_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|45|1 _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|45|B _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|45|RB _PG3_01|_DFF_P1|45|MID_SHUNT _PG3_01|_DFF_P1|A4  2.1704737578552e-12
B_PG3_01|_DFF_P1|6|1 _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|6|P _PG3_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|6|RB _PG3_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_PG|I_1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|I_1|MID  2e-12
I_PG3_01|_DFF_PG|I_1|B 0 _PG3_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|I_3|MID  2e-12
I_PG3_01|_DFF_PG|I_3|B 0 _PG3_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_PG|I_T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|I_T|MID  2e-12
I_PG3_01|_DFF_PG|I_T|B 0 _PG3_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|I_6|MID  2e-12
I_PG3_01|_DFF_PG|I_6|B 0 _PG3_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_PG|1|1 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|1|P _PG3_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|1|RB _PG3_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|23|1 _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|23|B _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|23|RB _PG3_01|_DFF_PG|23|MID_SHUNT _PG3_01|_DFF_PG|A3  2.1704737578552e-12
B_PG3_01|_DFF_PG|3|1 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|3|P _PG3_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|3|RB _PG3_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|4|1 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|4|P _PG3_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|4|B _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|4|RB _PG3_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|T|1 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|T|P _PG3_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|T|RB _PG3_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|45|1 _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|45|B _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|45|RB _PG3_01|_DFF_PG|45|MID_SHUNT _PG3_01|_DFF_PG|A4  2.1704737578552e-12
B_PG3_01|_DFF_PG|6|1 _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|6|P _PG3_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|6|RB _PG3_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_GG|I_1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|I_1|MID  2e-12
I_PG3_01|_DFF_GG|I_1|B 0 _PG3_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|I_3|MID  2e-12
I_PG3_01|_DFF_GG|I_3|B 0 _PG3_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_GG|I_T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|I_T|MID  2e-12
I_PG3_01|_DFF_GG|I_T|B 0 _PG3_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|I_6|MID  2e-12
I_PG3_01|_DFF_GG|I_6|B 0 _PG3_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_GG|1|1 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|1|P _PG3_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|1|RB _PG3_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|23|1 _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|23|B _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|23|RB _PG3_01|_DFF_GG|23|MID_SHUNT _PG3_01|_DFF_GG|A3  2.1704737578552e-12
B_PG3_01|_DFF_GG|3|1 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|3|P _PG3_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|3|RB _PG3_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|4|1 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|4|P _PG3_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|4|B _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|4|RB _PG3_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|T|1 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|T|P _PG3_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|T|RB _PG3_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|45|1 _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|45|B _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|45|RB _PG3_01|_DFF_GG|45|MID_SHUNT _PG3_01|_DFF_GG|A4  2.1704737578552e-12
B_PG3_01|_DFF_GG|6|1 _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|6|P _PG3_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|6|RB _PG3_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_G|I_A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|I_A1|MID  2e-12
I_PG3_01|_AND_G|I_A1|B 0 _PG3_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|I_B1|MID  2e-12
I_PG3_01|_AND_G|I_B1|B 0 _PG3_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q3|B _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|I_Q3|MID  2e-12
I_PG3_01|_AND_G|I_Q3|B 0 _PG3_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_G|I_Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|I_Q2|MID  2e-12
I_PG3_01|_AND_G|I_Q2|B 0 _PG3_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|I_Q1|MID  2e-12
I_PG3_01|_AND_G|I_Q1|B 0 _PG3_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_G|A1|1 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A1|P _PG3_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A1|RB _PG3_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A2|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A2|P _PG3_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A2|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A2|RB _PG3_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A12|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|A12|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|A12|RB _PG3_01|_AND_G|A12|MID_SHUNT _PG3_01|_AND_G|A3  2.1704737578552e-12
B_PG3_01|_AND_G|B1|1 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B1|P _PG3_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B1|RB _PG3_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B2|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B2|P _PG3_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B2|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B2|RB _PG3_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B12|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|B12|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|B12|RB _PG3_01|_AND_G|B12|MID_SHUNT _PG3_01|_AND_G|B3  2.1704737578552e-12
B_PG3_01|_AND_G|Q2|1 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q2|P _PG3_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q2|RB _PG3_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|Q1|1 _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q1|P _PG3_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q1|RB _PG3_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_P|I_A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|I_A1|MID  2e-12
I_PG3_01|_AND_P|I_A1|B 0 _PG3_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|I_B1|MID  2e-12
I_PG3_01|_AND_P|I_B1|B 0 _PG3_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q3|B _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|I_Q3|MID  2e-12
I_PG3_01|_AND_P|I_Q3|B 0 _PG3_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_P|I_Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|I_Q2|MID  2e-12
I_PG3_01|_AND_P|I_Q2|B 0 _PG3_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|I_Q1|MID  2e-12
I_PG3_01|_AND_P|I_Q1|B 0 _PG3_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_P|A1|1 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A1|P _PG3_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A1|RB _PG3_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A2|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A2|P _PG3_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A2|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A2|RB _PG3_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A12|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|A12|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|A12|RB _PG3_01|_AND_P|A12|MID_SHUNT _PG3_01|_AND_P|A3  2.1704737578552e-12
B_PG3_01|_AND_P|B1|1 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B1|P _PG3_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B1|RB _PG3_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B2|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B2|P _PG3_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B2|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B2|RB _PG3_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B12|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|B12|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|B12|RB _PG3_01|_AND_P|B12|MID_SHUNT _PG3_01|_AND_P|B3  2.1704737578552e-12
B_PG3_01|_AND_P|Q2|1 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q2|P _PG3_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q2|RB _PG3_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|Q1|1 _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q1|P _PG3_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q1|RB _PG3_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL1|I_D1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|I_D1|MID  2e-12
ISPL_G1_1|SPL1|I_D1|B 0 SPL_G1_1|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_D2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|I_D2|MID  2e-12
ISPL_G1_1|SPL1|I_D2|B 0 SPL_G1_1|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL1|I_Q1|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|I_Q1|MID  2e-12
ISPL_G1_1|SPL1|I_Q1|B 0 SPL_G1_1|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_Q2|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|I_Q2|MID  2e-12
ISPL_G1_1|SPL1|I_Q2|B 0 SPL_G1_1|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL1|1|1 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|1|P SPL_G1_1|SPL1|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|1|RB SPL_G1_1|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|2|1 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|2|P SPL_G1_1|SPL1|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|2|RB SPL_G1_1|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|A|1 SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|A|P SPL_G1_1|SPL1|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|A|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|A|RB SPL_G1_1|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|B|1 SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|B|P SPL_G1_1|SPL1|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|B|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|B|RB SPL_G1_1|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL2|I_D1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|I_D1|MID  2e-12
ISPL_G1_1|SPL2|I_D1|B 0 SPL_G1_1|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_D2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|I_D2|MID  2e-12
ISPL_G1_1|SPL2|I_D2|B 0 SPL_G1_1|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL2|I_Q1|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|I_Q1|MID  2e-12
ISPL_G1_1|SPL2|I_Q1|B 0 SPL_G1_1|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_Q2|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|I_Q2|MID  2e-12
ISPL_G1_1|SPL2|I_Q2|B 0 SPL_G1_1|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL2|1|1 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|1|P SPL_G1_1|SPL2|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|1|RB SPL_G1_1|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|2|1 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|2|P SPL_G1_1|SPL2|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|2|RB SPL_G1_1|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|A|1 SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|A|P SPL_G1_1|SPL2|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|A|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|A|RB SPL_G1_1|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|B|1 SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|B|P SPL_G1_1|SPL2|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|B|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|B|RB SPL_G1_1|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|P|I_1|B _PG0_12|P|A1 _PG0_12|P|I_1|MID  2e-12
I_PG0_12|P|I_1|B 0 _PG0_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_3|B _PG0_12|P|A3 _PG0_12|P|I_3|MID  2e-12
I_PG0_12|P|I_3|B 0 _PG0_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|P|I_T|B _PG0_12|P|T1 _PG0_12|P|I_T|MID  2e-12
I_PG0_12|P|I_T|B 0 _PG0_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_6|B _PG0_12|P|Q1 _PG0_12|P|I_6|MID  2e-12
I_PG0_12|P|I_6|B 0 _PG0_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|P|1|1 _PG0_12|P|A1 _PG0_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|1|P _PG0_12|P|1|MID_SERIES 0  2e-13
R_PG0_12|P|1|B _PG0_12|P|A1 _PG0_12|P|1|MID_SHUNT  2.7439617672
L_PG0_12|P|1|RB _PG0_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|23|1 _PG0_12|P|A2 _PG0_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|P|23|B _PG0_12|P|A2 _PG0_12|P|23|MID_SHUNT  3.84154647408
L_PG0_12|P|23|RB _PG0_12|P|23|MID_SHUNT _PG0_12|P|A3  2.1704737578552e-12
B_PG0_12|P|3|1 _PG0_12|P|A3 _PG0_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|3|P _PG0_12|P|3|MID_SERIES 0  2e-13
R_PG0_12|P|3|B _PG0_12|P|A3 _PG0_12|P|3|MID_SHUNT  2.7439617672
L_PG0_12|P|3|RB _PG0_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|4|1 _PG0_12|P|A4 _PG0_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|4|P _PG0_12|P|4|MID_SERIES 0  2e-13
R_PG0_12|P|4|B _PG0_12|P|A4 _PG0_12|P|4|MID_SHUNT  2.7439617672
L_PG0_12|P|4|RB _PG0_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|T|1 _PG0_12|P|T1 _PG0_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|T|P _PG0_12|P|T|MID_SERIES 0  2e-13
R_PG0_12|P|T|B _PG0_12|P|T1 _PG0_12|P|T|MID_SHUNT  2.7439617672
L_PG0_12|P|T|RB _PG0_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|45|1 _PG0_12|P|T2 _PG0_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|P|45|B _PG0_12|P|T2 _PG0_12|P|45|MID_SHUNT  3.84154647408
L_PG0_12|P|45|RB _PG0_12|P|45|MID_SHUNT _PG0_12|P|A4  2.1704737578552e-12
B_PG0_12|P|6|1 _PG0_12|P|Q1 _PG0_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|6|P _PG0_12|P|6|MID_SERIES 0  2e-13
R_PG0_12|P|6|B _PG0_12|P|Q1 _PG0_12|P|6|MID_SHUNT  2.7439617672
L_PG0_12|P|6|RB _PG0_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|G|I_1|B _PG0_12|G|A1 _PG0_12|G|I_1|MID  2e-12
I_PG0_12|G|I_1|B 0 _PG0_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_3|B _PG0_12|G|A3 _PG0_12|G|I_3|MID  2e-12
I_PG0_12|G|I_3|B 0 _PG0_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|G|I_T|B _PG0_12|G|T1 _PG0_12|G|I_T|MID  2e-12
I_PG0_12|G|I_T|B 0 _PG0_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_6|B _PG0_12|G|Q1 _PG0_12|G|I_6|MID  2e-12
I_PG0_12|G|I_6|B 0 _PG0_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|G|1|1 _PG0_12|G|A1 _PG0_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|1|P _PG0_12|G|1|MID_SERIES 0  2e-13
R_PG0_12|G|1|B _PG0_12|G|A1 _PG0_12|G|1|MID_SHUNT  2.7439617672
L_PG0_12|G|1|RB _PG0_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|23|1 _PG0_12|G|A2 _PG0_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|G|23|B _PG0_12|G|A2 _PG0_12|G|23|MID_SHUNT  3.84154647408
L_PG0_12|G|23|RB _PG0_12|G|23|MID_SHUNT _PG0_12|G|A3  2.1704737578552e-12
B_PG0_12|G|3|1 _PG0_12|G|A3 _PG0_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|3|P _PG0_12|G|3|MID_SERIES 0  2e-13
R_PG0_12|G|3|B _PG0_12|G|A3 _PG0_12|G|3|MID_SHUNT  2.7439617672
L_PG0_12|G|3|RB _PG0_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|4|1 _PG0_12|G|A4 _PG0_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|4|P _PG0_12|G|4|MID_SERIES 0  2e-13
R_PG0_12|G|4|B _PG0_12|G|A4 _PG0_12|G|4|MID_SHUNT  2.7439617672
L_PG0_12|G|4|RB _PG0_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|T|1 _PG0_12|G|T1 _PG0_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|T|P _PG0_12|G|T|MID_SERIES 0  2e-13
R_PG0_12|G|T|B _PG0_12|G|T1 _PG0_12|G|T|MID_SHUNT  2.7439617672
L_PG0_12|G|T|RB _PG0_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|45|1 _PG0_12|G|T2 _PG0_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|G|45|B _PG0_12|G|T2 _PG0_12|G|45|MID_SHUNT  3.84154647408
L_PG0_12|G|45|RB _PG0_12|G|45|MID_SHUNT _PG0_12|G|A4  2.1704737578552e-12
B_PG0_12|G|6|1 _PG0_12|G|Q1 _PG0_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|6|P _PG0_12|G|6|MID_SERIES 0  2e-13
R_PG0_12|G|6|B _PG0_12|G|Q1 _PG0_12|G|6|MID_SHUNT  2.7439617672
L_PG0_12|G|6|RB _PG0_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|I_D1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|I_D1|MID  2e-12
I_PG2_12|_SPL_G1|I_D1|B 0 _PG2_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_D2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|I_D2|MID  2e-12
I_PG2_12|_SPL_G1|I_D2|B 0 _PG2_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG2_12|_SPL_G1|I_Q1|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|I_Q1|MID  2e-12
I_PG2_12|_SPL_G1|I_Q1|B 0 _PG2_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_Q2|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|I_Q2|MID  2e-12
I_PG2_12|_SPL_G1|I_Q2|B 0 _PG2_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG2_12|_SPL_G1|1|1 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|1|P _PG2_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|1|RB _PG2_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|2|1 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|2|P _PG2_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|2|RB _PG2_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|A|1 _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|A|P _PG2_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|A|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|A|RB _PG2_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|B|1 _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|B|P _PG2_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|B|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|B|RB _PG2_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_PG|I_A1|B _PG2_12|_PG|A1 _PG2_12|_PG|I_A1|MID  2e-12
I_PG2_12|_PG|I_A1|B 0 _PG2_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_B1|B _PG2_12|_PG|B1 _PG2_12|_PG|I_B1|MID  2e-12
I_PG2_12|_PG|I_B1|B 0 _PG2_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q3|B _PG2_12|_PG|Q3 _PG2_12|_PG|I_Q3|MID  2e-12
I_PG2_12|_PG|I_Q3|B 0 _PG2_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_PG|I_Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|I_Q2|MID  2e-12
I_PG2_12|_PG|I_Q2|B 0 _PG2_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|I_Q1|MID  2e-12
I_PG2_12|_PG|I_Q1|B 0 _PG2_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_PG|A1|1 _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A1|P _PG2_12|_PG|A1|MID_SERIES 0  2e-13
R_PG2_12|_PG|A1|B _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A1|RB _PG2_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A2|1 _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A2|P _PG2_12|_PG|A2|MID_SERIES 0  2e-13
R_PG2_12|_PG|A2|B _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A2|RB _PG2_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A12|1 _PG2_12|_PG|A2 _PG2_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|A12|B _PG2_12|_PG|A2 _PG2_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|A12|RB _PG2_12|_PG|A12|MID_SHUNT _PG2_12|_PG|A3  2.1704737578552e-12
B_PG2_12|_PG|B1|1 _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B1|P _PG2_12|_PG|B1|MID_SERIES 0  2e-13
R_PG2_12|_PG|B1|B _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B1|RB _PG2_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B2|1 _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B2|P _PG2_12|_PG|B2|MID_SERIES 0  2e-13
R_PG2_12|_PG|B2|B _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B2|RB _PG2_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B12|1 _PG2_12|_PG|B2 _PG2_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|B12|B _PG2_12|_PG|B2 _PG2_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|B12|RB _PG2_12|_PG|B12|MID_SHUNT _PG2_12|_PG|B3  2.1704737578552e-12
B_PG2_12|_PG|Q2|1 _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q2|P _PG2_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q2|RB _PG2_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|Q1|1 _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q1|P _PG2_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q1|RB _PG2_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_GG|I_A1|B _PG2_12|_GG|A1 _PG2_12|_GG|I_A1|MID  2e-12
I_PG2_12|_GG|I_A1|B 0 _PG2_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_B1|B _PG2_12|_GG|B1 _PG2_12|_GG|I_B1|MID  2e-12
I_PG2_12|_GG|I_B1|B 0 _PG2_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q3|B _PG2_12|_GG|Q3 _PG2_12|_GG|I_Q3|MID  2e-12
I_PG2_12|_GG|I_Q3|B 0 _PG2_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_GG|I_Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|I_Q2|MID  2e-12
I_PG2_12|_GG|I_Q2|B 0 _PG2_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|I_Q1|MID  2e-12
I_PG2_12|_GG|I_Q1|B 0 _PG2_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_GG|A1|1 _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A1|P _PG2_12|_GG|A1|MID_SERIES 0  2e-13
R_PG2_12|_GG|A1|B _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A1|RB _PG2_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A2|1 _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A2|P _PG2_12|_GG|A2|MID_SERIES 0  2e-13
R_PG2_12|_GG|A2|B _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A2|RB _PG2_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A12|1 _PG2_12|_GG|A2 _PG2_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|A12|B _PG2_12|_GG|A2 _PG2_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|A12|RB _PG2_12|_GG|A12|MID_SHUNT _PG2_12|_GG|A3  2.1704737578552e-12
B_PG2_12|_GG|B1|1 _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B1|P _PG2_12|_GG|B1|MID_SERIES 0  2e-13
R_PG2_12|_GG|B1|B _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B1|RB _PG2_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B2|1 _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B2|P _PG2_12|_GG|B2|MID_SERIES 0  2e-13
R_PG2_12|_GG|B2|B _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B2|RB _PG2_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B12|1 _PG2_12|_GG|B2 _PG2_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|B12|B _PG2_12|_GG|B2 _PG2_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|B12|RB _PG2_12|_GG|B12|MID_SHUNT _PG2_12|_GG|B3  2.1704737578552e-12
B_PG2_12|_GG|Q2|1 _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q2|P _PG2_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q2|RB _PG2_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|Q1|1 _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q1|P _PG2_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q1|RB _PG2_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_PG|I_1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|I_1|MID  2e-12
I_PG2_12|_DFF_PG|I_1|B 0 _PG2_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|I_3|MID  2e-12
I_PG2_12|_DFF_PG|I_3|B 0 _PG2_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_PG|I_T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|I_T|MID  2e-12
I_PG2_12|_DFF_PG|I_T|B 0 _PG2_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|I_6|MID  2e-12
I_PG2_12|_DFF_PG|I_6|B 0 _PG2_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_PG|1|1 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|1|P _PG2_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|1|RB _PG2_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|23|1 _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|23|B _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|23|RB _PG2_12|_DFF_PG|23|MID_SHUNT _PG2_12|_DFF_PG|A3  2.1704737578552e-12
B_PG2_12|_DFF_PG|3|1 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|3|P _PG2_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|3|RB _PG2_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|4|1 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|4|P _PG2_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|4|B _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|4|RB _PG2_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|T|1 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|T|P _PG2_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|T|RB _PG2_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|45|1 _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|45|B _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|45|RB _PG2_12|_DFF_PG|45|MID_SHUNT _PG2_12|_DFF_PG|A4  2.1704737578552e-12
B_PG2_12|_DFF_PG|6|1 _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|6|P _PG2_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|6|RB _PG2_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_GG|I_1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|I_1|MID  2e-12
I_PG2_12|_DFF_GG|I_1|B 0 _PG2_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|I_3|MID  2e-12
I_PG2_12|_DFF_GG|I_3|B 0 _PG2_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_GG|I_T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|I_T|MID  2e-12
I_PG2_12|_DFF_GG|I_T|B 0 _PG2_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|I_6|MID  2e-12
I_PG2_12|_DFF_GG|I_6|B 0 _PG2_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_GG|1|1 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|1|P _PG2_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|1|RB _PG2_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|23|1 _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|23|B _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|23|RB _PG2_12|_DFF_GG|23|MID_SHUNT _PG2_12|_DFF_GG|A3  2.1704737578552e-12
B_PG2_12|_DFF_GG|3|1 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|3|P _PG2_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|3|RB _PG2_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|4|1 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|4|P _PG2_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|4|B _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|4|RB _PG2_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|T|1 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|T|P _PG2_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|T|RB _PG2_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|45|1 _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|45|B _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|45|RB _PG2_12|_DFF_GG|45|MID_SHUNT _PG2_12|_DFF_GG|A4  2.1704737578552e-12
B_PG2_12|_DFF_GG|6|1 _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|6|P _PG2_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|6|RB _PG2_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_G|I_A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|I_A1|MID  2e-12
I_PG2_12|_AND_G|I_A1|B 0 _PG2_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|I_B1|MID  2e-12
I_PG2_12|_AND_G|I_B1|B 0 _PG2_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q3|B _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|I_Q3|MID  2e-12
I_PG2_12|_AND_G|I_Q3|B 0 _PG2_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_G|I_Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|I_Q2|MID  2e-12
I_PG2_12|_AND_G|I_Q2|B 0 _PG2_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|I_Q1|MID  2e-12
I_PG2_12|_AND_G|I_Q1|B 0 _PG2_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_G|A1|1 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A1|P _PG2_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A1|RB _PG2_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A2|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A2|P _PG2_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A2|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A2|RB _PG2_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A12|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|A12|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|A12|RB _PG2_12|_AND_G|A12|MID_SHUNT _PG2_12|_AND_G|A3  2.1704737578552e-12
B_PG2_12|_AND_G|B1|1 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B1|P _PG2_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B1|RB _PG2_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B2|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B2|P _PG2_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B2|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B2|RB _PG2_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B12|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|B12|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|B12|RB _PG2_12|_AND_G|B12|MID_SHUNT _PG2_12|_AND_G|B3  2.1704737578552e-12
B_PG2_12|_AND_G|Q2|1 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q2|P _PG2_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q2|RB _PG2_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|Q1|1 _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q1|P _PG2_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q1|RB _PG2_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_SPL_G1|I_D1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|I_D1|MID  2e-12
I_PG3_12|_SPL_G1|I_D1|B 0 _PG3_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_D2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|I_D2|MID  2e-12
I_PG3_12|_SPL_G1|I_D2|B 0 _PG3_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_12|_SPL_G1|I_Q1|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|I_Q1|MID  2e-12
I_PG3_12|_SPL_G1|I_Q1|B 0 _PG3_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_Q2|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|I_Q2|MID  2e-12
I_PG3_12|_SPL_G1|I_Q2|B 0 _PG3_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_12|_SPL_G1|1|1 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|1|P _PG3_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|1|RB _PG3_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|2|1 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|2|P _PG3_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|2|RB _PG3_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|A|1 _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|A|P _PG3_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|A|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|A|RB _PG3_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|B|1 _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|B|P _PG3_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|B|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|B|RB _PG3_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_PG|I_A1|B _PG3_12|_PG|A1 _PG3_12|_PG|I_A1|MID  2e-12
I_PG3_12|_PG|I_A1|B 0 _PG3_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_B1|B _PG3_12|_PG|B1 _PG3_12|_PG|I_B1|MID  2e-12
I_PG3_12|_PG|I_B1|B 0 _PG3_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q3|B _PG3_12|_PG|Q3 _PG3_12|_PG|I_Q3|MID  2e-12
I_PG3_12|_PG|I_Q3|B 0 _PG3_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_PG|I_Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|I_Q2|MID  2e-12
I_PG3_12|_PG|I_Q2|B 0 _PG3_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|I_Q1|MID  2e-12
I_PG3_12|_PG|I_Q1|B 0 _PG3_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_PG|A1|1 _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A1|P _PG3_12|_PG|A1|MID_SERIES 0  2e-13
R_PG3_12|_PG|A1|B _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A1|RB _PG3_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A2|1 _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A2|P _PG3_12|_PG|A2|MID_SERIES 0  2e-13
R_PG3_12|_PG|A2|B _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A2|RB _PG3_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A12|1 _PG3_12|_PG|A2 _PG3_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|A12|B _PG3_12|_PG|A2 _PG3_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|A12|RB _PG3_12|_PG|A12|MID_SHUNT _PG3_12|_PG|A3  2.1704737578552e-12
B_PG3_12|_PG|B1|1 _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B1|P _PG3_12|_PG|B1|MID_SERIES 0  2e-13
R_PG3_12|_PG|B1|B _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B1|RB _PG3_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B2|1 _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B2|P _PG3_12|_PG|B2|MID_SERIES 0  2e-13
R_PG3_12|_PG|B2|B _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B2|RB _PG3_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B12|1 _PG3_12|_PG|B2 _PG3_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|B12|B _PG3_12|_PG|B2 _PG3_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|B12|RB _PG3_12|_PG|B12|MID_SHUNT _PG3_12|_PG|B3  2.1704737578552e-12
B_PG3_12|_PG|Q2|1 _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q2|P _PG3_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q2|RB _PG3_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|Q1|1 _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q1|P _PG3_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q1|RB _PG3_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_GG|I_A1|B _PG3_12|_GG|A1 _PG3_12|_GG|I_A1|MID  2e-12
I_PG3_12|_GG|I_A1|B 0 _PG3_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_B1|B _PG3_12|_GG|B1 _PG3_12|_GG|I_B1|MID  2e-12
I_PG3_12|_GG|I_B1|B 0 _PG3_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q3|B _PG3_12|_GG|Q3 _PG3_12|_GG|I_Q3|MID  2e-12
I_PG3_12|_GG|I_Q3|B 0 _PG3_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_GG|I_Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|I_Q2|MID  2e-12
I_PG3_12|_GG|I_Q2|B 0 _PG3_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|I_Q1|MID  2e-12
I_PG3_12|_GG|I_Q1|B 0 _PG3_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_GG|A1|1 _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A1|P _PG3_12|_GG|A1|MID_SERIES 0  2e-13
R_PG3_12|_GG|A1|B _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A1|RB _PG3_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A2|1 _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A2|P _PG3_12|_GG|A2|MID_SERIES 0  2e-13
R_PG3_12|_GG|A2|B _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A2|RB _PG3_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A12|1 _PG3_12|_GG|A2 _PG3_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|A12|B _PG3_12|_GG|A2 _PG3_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|A12|RB _PG3_12|_GG|A12|MID_SHUNT _PG3_12|_GG|A3  2.1704737578552e-12
B_PG3_12|_GG|B1|1 _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B1|P _PG3_12|_GG|B1|MID_SERIES 0  2e-13
R_PG3_12|_GG|B1|B _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B1|RB _PG3_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B2|1 _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B2|P _PG3_12|_GG|B2|MID_SERIES 0  2e-13
R_PG3_12|_GG|B2|B _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B2|RB _PG3_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B12|1 _PG3_12|_GG|B2 _PG3_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|B12|B _PG3_12|_GG|B2 _PG3_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|B12|RB _PG3_12|_GG|B12|MID_SHUNT _PG3_12|_GG|B3  2.1704737578552e-12
B_PG3_12|_GG|Q2|1 _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q2|P _PG3_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q2|RB _PG3_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|Q1|1 _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q1|P _PG3_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q1|RB _PG3_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_PG|I_1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|I_1|MID  2e-12
I_PG3_12|_DFF_PG|I_1|B 0 _PG3_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|I_3|MID  2e-12
I_PG3_12|_DFF_PG|I_3|B 0 _PG3_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_PG|I_T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|I_T|MID  2e-12
I_PG3_12|_DFF_PG|I_T|B 0 _PG3_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|I_6|MID  2e-12
I_PG3_12|_DFF_PG|I_6|B 0 _PG3_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_PG|1|1 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|1|P _PG3_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|1|RB _PG3_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|23|1 _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|23|B _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|23|RB _PG3_12|_DFF_PG|23|MID_SHUNT _PG3_12|_DFF_PG|A3  2.1704737578552e-12
B_PG3_12|_DFF_PG|3|1 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|3|P _PG3_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|3|RB _PG3_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|4|1 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|4|P _PG3_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|4|B _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|4|RB _PG3_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|T|1 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|T|P _PG3_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|T|RB _PG3_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|45|1 _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|45|B _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|45|RB _PG3_12|_DFF_PG|45|MID_SHUNT _PG3_12|_DFF_PG|A4  2.1704737578552e-12
B_PG3_12|_DFF_PG|6|1 _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|6|P _PG3_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|6|RB _PG3_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_GG|I_1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|I_1|MID  2e-12
I_PG3_12|_DFF_GG|I_1|B 0 _PG3_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|I_3|MID  2e-12
I_PG3_12|_DFF_GG|I_3|B 0 _PG3_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_GG|I_T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|I_T|MID  2e-12
I_PG3_12|_DFF_GG|I_T|B 0 _PG3_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|I_6|MID  2e-12
I_PG3_12|_DFF_GG|I_6|B 0 _PG3_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_GG|1|1 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|1|P _PG3_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|1|RB _PG3_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|23|1 _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|23|B _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|23|RB _PG3_12|_DFF_GG|23|MID_SHUNT _PG3_12|_DFF_GG|A3  2.1704737578552e-12
B_PG3_12|_DFF_GG|3|1 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|3|P _PG3_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|3|RB _PG3_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|4|1 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|4|P _PG3_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|4|B _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|4|RB _PG3_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|T|1 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|T|P _PG3_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|T|RB _PG3_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|45|1 _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|45|B _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|45|RB _PG3_12|_DFF_GG|45|MID_SHUNT _PG3_12|_DFF_GG|A4  2.1704737578552e-12
B_PG3_12|_DFF_GG|6|1 _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|6|P _PG3_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|6|RB _PG3_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_G|I_A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|I_A1|MID  2e-12
I_PG3_12|_AND_G|I_A1|B 0 _PG3_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|I_B1|MID  2e-12
I_PG3_12|_AND_G|I_B1|B 0 _PG3_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q3|B _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|I_Q3|MID  2e-12
I_PG3_12|_AND_G|I_Q3|B 0 _PG3_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_G|I_Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|I_Q2|MID  2e-12
I_PG3_12|_AND_G|I_Q2|B 0 _PG3_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|I_Q1|MID  2e-12
I_PG3_12|_AND_G|I_Q1|B 0 _PG3_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_G|A1|1 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A1|P _PG3_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A1|RB _PG3_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A2|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A2|P _PG3_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A2|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A2|RB _PG3_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A12|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|A12|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|A12|RB _PG3_12|_AND_G|A12|MID_SHUNT _PG3_12|_AND_G|A3  2.1704737578552e-12
B_PG3_12|_AND_G|B1|1 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B1|P _PG3_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B1|RB _PG3_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B2|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B2|P _PG3_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B2|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B2|RB _PG3_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B12|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|B12|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|B12|RB _PG3_12|_AND_G|B12|MID_SHUNT _PG3_12|_AND_G|B3  2.1704737578552e-12
B_PG3_12|_AND_G|Q2|1 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q2|P _PG3_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q2|RB _PG3_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|Q1|1 _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q1|P _PG3_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q1|RB _PG3_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_S0
.print DEVI R_S1
.print DEVI R_S2
.print DEVI R_S3
.print DEVI R_S4
.print V IP0_0_RX
.print V G1_2
.print V G2_2
.print V S2
.print V IG0_0_TO1
.print V T07
.print V P0_2_RX
.print V IP2_0
.print V D03
.print V G0_1_RX
.print V T00
.print V P0_1
.print V IG1_0
.print V T11
.print V IP1_0_RX
.print V IP1_1_OUT
.print V B0
.print V IP3_2_OUT_RX
.print V P2_1
.print V B2_RX
.print V IP1_1_OUT_RX
.print V IP3_2_OUT
.print V P2_1_RX
.print V IG2_0
.print V G2_1_RX
.print V B3
.print V T03
.print V T15
.print V G3_1
.print V IP3_0_TO1
.print V G2_1
.print V IP2_0_TO2
.print V B2
.print V IP1_2_OUT
.print V B0_RX
.print V G1_1
.print V G0_2
.print V S3
.print V G2_2_RX
.print V IP1_0_TO1
.print V S1
.print V T14
.print V T08
.print V IG2_0_RX
.print V T02
.print V T09
.print V T16
.print V G1_2_RX
.print V IP1_2_OUT_RX
.print V IG1_0_RX
.print V G1_1_RX
.print V T04
.print V T12
.print V IG0_0_RX
.print V G1_1_TO1
.print V A2
.print V IP0_0
.print V IP3_0_OUT
.print V IG0_0_TO0
.print V P3_1
.print V G1_1_TO3
.print V S4
.print V A0
.print V A2_RX
.print V IP2_2_OUT
.print V A3
.print V IP2_0_TO3
.print V T01
.print V T10
.print V IP2_1_OUT
.print V D02
.print V B1_RX
.print V B3_RX
.print V T13
.print V IP3_1_OUT_RX
.print V IP1_0
.print V IP3_0_RX
.print V IP3_0
.print V P0_1_RX
.print V IP3_1_OUT
.print V T06
.print V G3_1_RX
.print V IG3_0
.print V A0_RX
.print V IG2_0_TO3
.print V G0_1
.print V IP2_0_RX
.print V G3_2_RX
.print V D01
.print V P0_2
.print V D13
.print V S0
.print V IG2_0_TO2
.print V G3_2
.print V A1
.print V IG3_0_RX
.print V A3_RX
.print V B1
.print V IP2_0_OUT
.print V IP2_1_OUT_RX
.print V G1_1_TO2
.print V P3_1_RX
.print V IG0_0
.print V D11
.print V D12
.print V T05
.print V A1_RX
.print V IP1_0_OUT
.print V G0_2_RX
.print V IP2_2_OUT_RX
