*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=5e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM IU=1.25e-05
.PARAM VU=0.0006857
.PARAM LU=2.632e-12
.PARAM ICRECEIVE=1.6
.PARAM ICTRANS=2.5
.PARAM RD=1.36
.PARAM OFFSET1=5e-11
.PARAM TCLOCK=2.5e-10
.PARAM DO=6.25e-11
.PARAM ZED0=5
.PARAM IMAX=0.0006
.PARAM TR=9.5e-12
.PARAM TF=9.5e-12
.PARAM PW=1e-12
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL	JJMIT	JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
TCLK  CLK_TX  0 CLK 0 LOSSLESS Z0=ZED0 TD=1P
TA    A_TX    0 A   0 LOSSLESS Z0=ZED0 TD=1P
TSUM SUM_TX  0 SUM  0  LOSSLESS Z0=ZED0 TD=1P
TCARRY CARRY_TX  0 CARRY  0  LOSSLESS Z0=ZED0 TD=1P
TCBAR CBAR_TX  0 CBAR  0  LOSSLESS Z0=ZED0 TD=1P
.TRAN 0.25E-12 2.6E-9
ICLK 0 CLK_DC  PULSE(0 IMAX OFFSET1               TR TF PW   TCLOCK)
IA1_1 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+1*TCLOCK TR TF PW 8*TCLOCK)
IA1_2 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+3*TCLOCK TR TF PW 8*TCLOCK)
IA1_3 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+5*TCLOCK TR TF PW 8*TCLOCK)
IA1_4 0 A1_DC  PULSE(0 IMAX OFFSET1+1*DO+7*TCLOCK TR TF PW 8*TCLOCK)
IA2_1 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+2*TCLOCK TR TF PW 8*TCLOCK)
IA2_2 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+3*TCLOCK TR TF PW 8*TCLOCK)
IA2_3 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+6*TCLOCK TR TF PW 8*TCLOCK)
IA2_4 0 A1_DC  PULSE(0 IMAX OFFSET1+2*DO+7*TCLOCK TR TF PW 8*TCLOCK)
IA3_1 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+4*TCLOCK TR TF PW 8*TCLOCK)
IA3_2 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+5*TCLOCK TR TF PW 8*TCLOCK)
IA3_3 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+6*TCLOCK TR TF PW 8*TCLOCK)
IA3_4 0 A1_DC  PULSE(0 IMAX OFFSET1+3*DO+7*TCLOCK TR TF PW 8*TCLOCK)
RSUM SUM 0  1
RCARRY CARRY 0  1
RCBAR CBAR 0  1
BDCSFQCLK|1 DCSFQCLK|2 DCSFQCLK|3 JJMIT AREA=2.25
BDCSFQCLK|2 DCSFQCLK|5 DCSFQCLK|6 JJMIT AREA=2.25
BDCSFQCLK|3 DCSFQCLK|7 DCSFQCLK|8 JJMIT AREA=2.5
BDCSFQCLK|4 DCSFQCLK|11 DCSFQCLK|12 JJMIT AREA=2.5
IDCSFQCLK|B1 0 DCSFQCLK|4  0.00027500000000000007
IDCSFQCLK|B2 0 DCSFQCLK|10  0.00034999999999999994
LDCSFQCLK|B1 DCSFQCLK|4 DCSFQCLK|3  2e-12
LDCSFQCLK|B2 DCSFQCLK|10 DCSFQCLK|9  2e-12
LDCSFQCLK|P2 DCSFQCLK|6 0  5e-13
LDCSFQCLK|P3 DCSFQCLK|8 0  5e-13
LDCSFQCLK|P4 DCSFQCLK|12 0  5e-13
LDCSFQCLK|1 CLK_DC DCSFQCLK|1  1e-12
LDCSFQCLK|2 DCSFQCLK|1 0  3.9e-12
LDCSFQCLK|3 DCSFQCLK|1 DCSFQCLK|2  6e-13
LDCSFQCLK|4 DCSFQCLK|3 DCSFQCLK|5  1.1e-12
LDCSFQCLK|5 DCSFQCLK|5 DCSFQCLK|7  4.5951863288888885e-12
LDCSFQCLK|6 DCSFQCLK|7 DCSFQCLK|9  2.067833848e-12
LDCSFQCLK|7 DCSFQCLK|9 DCSFQCLK|11  2.067833848e-12
LDCSFQCLK|8 DCSFQCLK|11 DCSFQCLK|13  2e-12
RDCSFQCLK|D DCSFQCLK|13 CLK_TX  1.36
RDCSFQCLK|B1 DCSFQCLK|2 DCSFQCLK|102  3.048846408
LDCSFQCLK|RB1 DCSFQCLK|102 DCSFQCLK|3  1.7225982205200002e-12
RDCSFQCLK|B2 DCSFQCLK|5 DCSFQCLK|105  3.048846408
LDCSFQCLK|RB2 DCSFQCLK|105 0  2.2225982205200003e-12
RDCSFQCLK|B3 DCSFQCLK|7 DCSFQCLK|107  2.7439617672
LDCSFQCLK|RB3 DCSFQCLK|107 0  2.050338398468e-12
RDCSFQCLK|B4 DCSFQCLK|11 DCSFQCLK|111  2.7439617672
LDCSFQCLK|RB4 DCSFQCLK|111 0  2.050338398468e-12
BDCSFQ_1|1 DCSFQ_1|2 DCSFQ_1|3 JJMIT AREA=2.25
BDCSFQ_1|2 DCSFQ_1|5 DCSFQ_1|6 JJMIT AREA=2.25
BDCSFQ_1|3 DCSFQ_1|7 DCSFQ_1|8 JJMIT AREA=2.5
BDCSFQ_1|4 DCSFQ_1|11 DCSFQ_1|12 JJMIT AREA=2.5
IDCSFQ_1|B1 0 DCSFQ_1|4  0.00027500000000000007
IDCSFQ_1|B2 0 DCSFQ_1|10  0.00034999999999999994
LDCSFQ_1|B1 DCSFQ_1|4 DCSFQ_1|3  2e-12
LDCSFQ_1|B2 DCSFQ_1|10 DCSFQ_1|9  2e-12
LDCSFQ_1|P2 DCSFQ_1|6 0  5e-13
LDCSFQ_1|P3 DCSFQ_1|8 0  5e-13
LDCSFQ_1|P4 DCSFQ_1|12 0  5e-13
LDCSFQ_1|1 A1_DC DCSFQ_1|1  1e-12
LDCSFQ_1|2 DCSFQ_1|1 0  3.9e-12
LDCSFQ_1|3 DCSFQ_1|1 DCSFQ_1|2  6e-13
LDCSFQ_1|4 DCSFQ_1|3 DCSFQ_1|5  1.1e-12
LDCSFQ_1|5 DCSFQ_1|5 DCSFQ_1|7  4.5951863288888885e-12
LDCSFQ_1|6 DCSFQ_1|7 DCSFQ_1|9  2.067833848e-12
LDCSFQ_1|7 DCSFQ_1|9 DCSFQ_1|11  2.067833848e-12
LDCSFQ_1|8 DCSFQ_1|11 DCSFQ_1|13  2e-12
RDCSFQ_1|D DCSFQ_1|13 A_TX  1.36
RDCSFQ_1|B1 DCSFQ_1|2 DCSFQ_1|102  3.048846408
LDCSFQ_1|RB1 DCSFQ_1|102 DCSFQ_1|3  1.7225982205200002e-12
RDCSFQ_1|B2 DCSFQ_1|5 DCSFQ_1|105  3.048846408
LDCSFQ_1|RB2 DCSFQ_1|105 0  2.2225982205200003e-12
RDCSFQ_1|B3 DCSFQ_1|7 DCSFQ_1|107  2.7439617672
LDCSFQ_1|RB3 DCSFQ_1|107 0  2.050338398468e-12
RDCSFQ_1|B4 DCSFQ_1|11 DCSFQ_1|111  2.7439617672
LDCSFQ_1|RB4 DCSFQ_1|111 0  2.050338398468e-12
L_TFF|6 _TFF|READOUT _TFF|1  5.26e-12
B_TFF|11 _TFF|1 _TFF|2 JJMIT 
B_TFF|10 _TFF|2 0 JJMIT 
L_TFF|8 _TFF|2 _TFF|SUM_TX  3.9e-12
B_TFF|12 _TFF|2 _TFF|4 JJMIT 
B_TFF|6 _TFF|4 _TFF|6 JJMIT 
L_TFF|1 _TFF|3 _TFF|4  5.26e-12
L_TFF|3 _TFF|3 _TFF|CBAR_TX  5.26e-12
B_TFF|1 _TFF|3 0 JJMIT 
B_TFF|2 _TFF|3 _TFF|5 JJMIT 
B_TFF|5 _TFF|5 _TFF|6 JJMIT 
L_TFF|4 _TFF|6 _TFF|CARRY_TX  5.26e-12
B_TFF|4 _TFF|6 0 JJMIT 
L_TFF|2 _TFF|5 _TFF|7  1.3e-12
B_TFF|3 _TFF|7 0 JJMIT 
L_TFF|7 _TFF|7 _TFF|TOGGLE  2.63e-12
B_TFF|_READOUT|1 _TFF|_READOUT|1 _TFF|_READOUT|2 JJMIT AREA=1.6
B_TFF|_READOUT|2 _TFF|_READOUT|4 _TFF|_READOUT|5 JJMIT AREA=2.0
B_TFF|_READOUT|3 _TFF|_READOUT|7 _TFF|_READOUT|8 JJMIT AREA=2.5
I_TFF|_READOUT|B1 0 _TFF|_READOUT|3  0.000112
I_TFF|_READOUT|B2 0 _TFF|_READOUT|6  0.0002
I_TFF|_READOUT|B3 0 _TFF|_READOUT|9  0.00017499999999999997
L_TFF|_READOUT|B1 _TFF|_READOUT|3 _TFF|_READOUT|1  2e-12
L_TFF|_READOUT|B2 _TFF|_READOUT|6 _TFF|_READOUT|4  2e-12
L_TFF|_READOUT|B3 _TFF|_READOUT|9 _TFF|_READOUT|7  2e-12
L_TFF|_READOUT|1 CLK _TFF|_READOUT|1  2e-12
L_TFF|_READOUT|2 _TFF|_READOUT|1 _TFF|_READOUT|4  6.461980775e-12
L_TFF|_READOUT|3 _TFF|_READOUT|4 _TFF|_READOUT|7  5.16958462e-12
L_TFF|_READOUT|4 _TFF|_READOUT|7 _TFF|READOUT  2.067833848e-12
L_TFF|_READOUT|P1 _TFF|_READOUT|2 0  5e-13
L_TFF|_READOUT|P2 _TFF|_READOUT|5 0  5e-13
L_TFF|_READOUT|P3 _TFF|_READOUT|8 0  5e-13
R_TFF|_READOUT|B1 _TFF|_READOUT|1 _TFF|_READOUT|101  4.2874402612499996
L_TFF|_READOUT|RB1 _TFF|_READOUT|101 0  2.92240374760625e-12
R_TFF|_READOUT|B2 _TFF|_READOUT|4 _TFF|_READOUT|104  3.429952209
L_TFF|_READOUT|RB2 _TFF|_READOUT|104 0  2.437922998085e-12
R_TFF|_READOUT|B3 _TFF|_READOUT|7 _TFF|_READOUT|107  2.7439617672
L_TFF|_READOUT|RB3 _TFF|_READOUT|107 0  2.050338398468e-12
B_TFF|_TOGGLE|1 _TFF|_TOGGLE|1 _TFF|_TOGGLE|2 JJMIT AREA=1.6
B_TFF|_TOGGLE|2 _TFF|_TOGGLE|4 _TFF|_TOGGLE|5 JJMIT AREA=2.0
B_TFF|_TOGGLE|3 _TFF|_TOGGLE|7 _TFF|_TOGGLE|8 JJMIT AREA=2.5
I_TFF|_TOGGLE|B1 0 _TFF|_TOGGLE|3  0.000112
I_TFF|_TOGGLE|B2 0 _TFF|_TOGGLE|6  0.0002
I_TFF|_TOGGLE|B3 0 _TFF|_TOGGLE|9  0.00017499999999999997
L_TFF|_TOGGLE|B1 _TFF|_TOGGLE|3 _TFF|_TOGGLE|1  2e-12
L_TFF|_TOGGLE|B2 _TFF|_TOGGLE|6 _TFF|_TOGGLE|4  2e-12
L_TFF|_TOGGLE|B3 _TFF|_TOGGLE|9 _TFF|_TOGGLE|7  2e-12
L_TFF|_TOGGLE|1 A _TFF|_TOGGLE|1  2e-12
L_TFF|_TOGGLE|2 _TFF|_TOGGLE|1 _TFF|_TOGGLE|4  6.461980775e-12
L_TFF|_TOGGLE|3 _TFF|_TOGGLE|4 _TFF|_TOGGLE|7  5.16958462e-12
L_TFF|_TOGGLE|4 _TFF|_TOGGLE|7 _TFF|TOGGLE  2.067833848e-12
L_TFF|_TOGGLE|P1 _TFF|_TOGGLE|2 0  5e-13
L_TFF|_TOGGLE|P2 _TFF|_TOGGLE|5 0  5e-13
L_TFF|_TOGGLE|P3 _TFF|_TOGGLE|8 0  5e-13
R_TFF|_TOGGLE|B1 _TFF|_TOGGLE|1 _TFF|_TOGGLE|101  4.2874402612499996
L_TFF|_TOGGLE|RB1 _TFF|_TOGGLE|101 0  2.92240374760625e-12
R_TFF|_TOGGLE|B2 _TFF|_TOGGLE|4 _TFF|_TOGGLE|104  3.429952209
L_TFF|_TOGGLE|RB2 _TFF|_TOGGLE|104 0  2.437922998085e-12
R_TFF|_TOGGLE|B3 _TFF|_TOGGLE|7 _TFF|_TOGGLE|107  2.7439617672
L_TFF|_TOGGLE|RB3 _TFF|_TOGGLE|107 0  2.050338398468e-12
B_TFF|_SUM|1 _TFF|_SUM|1 _TFF|_SUM|2 JJMIT AREA=2.5
B_TFF|_SUM|2 _TFF|_SUM|4 _TFF|_SUM|5 JJMIT AREA=2.5
I_TFF|_SUM|B1 0 _TFF|_SUM|3  0.00017499999999999997
I_TFF|_SUM|B2 0 _TFF|_SUM|6  0.00017499999999999997
L_TFF|_SUM|B1 _TFF|_SUM|3 _TFF|_SUM|1  2e-12
L_TFF|_SUM|B2 _TFF|_SUM|6 _TFF|_SUM|4  2e-12
L_TFF|_SUM|1 _TFF|SUM_TX _TFF|_SUM|1  2.067833848e-12
L_TFF|_SUM|2 _TFF|_SUM|1 _TFF|_SUM|4  4.135667696e-12
L_TFF|_SUM|3 _TFF|_SUM|4 _TFF|_SUM|7  2e-12
L_TFF|_SUM|P1 _TFF|_SUM|2 0  5e-13
L_TFF|_SUM|P2 _TFF|_SUM|5 0  5e-13
R_TFF|_SUM|D _TFF|_SUM|7 SUM_TX  1.36
R_TFF|_SUM|B1 _TFF|_SUM|1 _TFF|_SUM|101  2.7439617672
L_TFF|_SUM|RB1 _TFF|_SUM|101 0  2.050338398468e-12
R_TFF|_SUM|B2 _TFF|_SUM|4 _TFF|_SUM|104  2.7439617672
L_TFF|_SUM|RB2 _TFF|_SUM|104 0  2.050338398468e-12
B_TFF|_CARRY|1 _TFF|_CARRY|1 _TFF|_CARRY|2 JJMIT AREA=2.5
B_TFF|_CARRY|2 _TFF|_CARRY|4 _TFF|_CARRY|5 JJMIT AREA=2.5
I_TFF|_CARRY|B1 0 _TFF|_CARRY|3  0.00017499999999999997
I_TFF|_CARRY|B2 0 _TFF|_CARRY|6  0.00017499999999999997
L_TFF|_CARRY|B1 _TFF|_CARRY|3 _TFF|_CARRY|1  2e-12
L_TFF|_CARRY|B2 _TFF|_CARRY|6 _TFF|_CARRY|4  2e-12
L_TFF|_CARRY|1 _TFF|CARRY_TX _TFF|_CARRY|1  2.067833848e-12
L_TFF|_CARRY|2 _TFF|_CARRY|1 _TFF|_CARRY|4  4.135667696e-12
L_TFF|_CARRY|3 _TFF|_CARRY|4 _TFF|_CARRY|7  2e-12
L_TFF|_CARRY|P1 _TFF|_CARRY|2 0  5e-13
L_TFF|_CARRY|P2 _TFF|_CARRY|5 0  5e-13
R_TFF|_CARRY|D _TFF|_CARRY|7 CARRY_TX  1.36
R_TFF|_CARRY|B1 _TFF|_CARRY|1 _TFF|_CARRY|101  2.7439617672
L_TFF|_CARRY|RB1 _TFF|_CARRY|101 0  2.050338398468e-12
R_TFF|_CARRY|B2 _TFF|_CARRY|4 _TFF|_CARRY|104  2.7439617672
L_TFF|_CARRY|RB2 _TFF|_CARRY|104 0  2.050338398468e-12
B_TFF|_CBAR|1 _TFF|_CBAR|1 _TFF|_CBAR|2 JJMIT AREA=2.5
B_TFF|_CBAR|2 _TFF|_CBAR|4 _TFF|_CBAR|5 JJMIT AREA=2.5
I_TFF|_CBAR|B1 0 _TFF|_CBAR|3  0.00017499999999999997
I_TFF|_CBAR|B2 0 _TFF|_CBAR|6  0.00017499999999999997
L_TFF|_CBAR|B1 _TFF|_CBAR|3 _TFF|_CBAR|1  2e-12
L_TFF|_CBAR|B2 _TFF|_CBAR|6 _TFF|_CBAR|4  2e-12
L_TFF|_CBAR|1 _TFF|CBAR_TX _TFF|_CBAR|1  2.067833848e-12
L_TFF|_CBAR|2 _TFF|_CBAR|1 _TFF|_CBAR|4  4.135667696e-12
L_TFF|_CBAR|3 _TFF|_CBAR|4 _TFF|_CBAR|7  2e-12
L_TFF|_CBAR|P1 _TFF|_CBAR|2 0  5e-13
L_TFF|_CBAR|P2 _TFF|_CBAR|5 0  5e-13
R_TFF|_CBAR|D _TFF|_CBAR|7 CBAR_TX  1.36
R_TFF|_CBAR|B1 _TFF|_CBAR|1 _TFF|_CBAR|101  2.7439617672
L_TFF|_CBAR|RB1 _TFF|_CBAR|101 0  2.050338398468e-12
R_TFF|_CBAR|B2 _TFF|_CBAR|4 _TFF|_CBAR|104  2.7439617672
L_TFF|_CBAR|RB2 _TFF|_CBAR|104 0  2.050338398468e-12
L_TFF|I1|B _TFF|3 _TFF|I1|MID  2e-12
I_TFF|I1|B 0 _TFF|I1|MID  PWL(0 0 5e-12 0.00019)
L_TFF|I2|B _TFF|7 _TFF|I2|MID  2e-12
I_TFF|I2|B 0 _TFF|I2|MID  PWL(0 0 5e-12 0.00019)
.print DEVI ICLK
.print DEVI IA1_1
.print DEVI IA1_2
.print DEVI IA1_3
.print DEVI IA1_4
.print DEVI IA2_1
.print DEVI IA2_2
.print DEVI IA2_3
.print DEVI IA2_4
.print DEVI IA3_1
.print DEVI IA3_2
.print DEVI IA3_3
.print DEVI IA3_4
.print DEVI RSUM
.print DEVI RCARRY
.print DEVI RCBAR
.print DEVI BDCSFQCLK|1
.print DEVI BDCSFQCLK|2
.print DEVI BDCSFQCLK|3
.print DEVI BDCSFQCLK|4
.print DEVI IDCSFQCLK|B1
.print DEVI IDCSFQCLK|B2
.print DEVI LDCSFQCLK|B1
.print DEVI LDCSFQCLK|B2
.print DEVI LDCSFQCLK|P2
.print DEVI LDCSFQCLK|P3
.print DEVI LDCSFQCLK|P4
.print DEVI LDCSFQCLK|1
.print DEVI LDCSFQCLK|2
.print DEVI LDCSFQCLK|3
.print DEVI LDCSFQCLK|4
.print DEVI LDCSFQCLK|5
.print DEVI LDCSFQCLK|6
.print DEVI LDCSFQCLK|7
.print DEVI LDCSFQCLK|8
.print DEVI RDCSFQCLK|D
.print DEVI RDCSFQCLK|B1
.print DEVI LDCSFQCLK|RB1
.print DEVI RDCSFQCLK|B2
.print DEVI LDCSFQCLK|RB2
.print DEVI RDCSFQCLK|B3
.print DEVI LDCSFQCLK|RB3
.print DEVI RDCSFQCLK|B4
.print DEVI LDCSFQCLK|RB4
.print DEVI BDCSFQ_1|1
.print DEVI BDCSFQ_1|2
.print DEVI BDCSFQ_1|3
.print DEVI BDCSFQ_1|4
.print DEVI IDCSFQ_1|B1
.print DEVI IDCSFQ_1|B2
.print DEVI LDCSFQ_1|B1
.print DEVI LDCSFQ_1|B2
.print DEVI LDCSFQ_1|P2
.print DEVI LDCSFQ_1|P3
.print DEVI LDCSFQ_1|P4
.print DEVI LDCSFQ_1|1
.print DEVI LDCSFQ_1|2
.print DEVI LDCSFQ_1|3
.print DEVI LDCSFQ_1|4
.print DEVI LDCSFQ_1|5
.print DEVI LDCSFQ_1|6
.print DEVI LDCSFQ_1|7
.print DEVI LDCSFQ_1|8
.print DEVI RDCSFQ_1|D
.print DEVI RDCSFQ_1|B1
.print DEVI LDCSFQ_1|RB1
.print DEVI RDCSFQ_1|B2
.print DEVI LDCSFQ_1|RB2
.print DEVI RDCSFQ_1|B3
.print DEVI LDCSFQ_1|RB3
.print DEVI RDCSFQ_1|B4
.print DEVI LDCSFQ_1|RB4
.print DEVI L_TFF|6
.print DEVI B_TFF|11
.print DEVI B_TFF|10
.print DEVI L_TFF|8
.print DEVI B_TFF|12
.print DEVI B_TFF|6
.print DEVI L_TFF|1
.print DEVI L_TFF|3
.print DEVI B_TFF|1
.print DEVI B_TFF|2
.print DEVI B_TFF|5
.print DEVI L_TFF|4
.print DEVI B_TFF|4
.print DEVI L_TFF|2
.print DEVI B_TFF|3
.print DEVI L_TFF|7
.print V DCSFQCLK|111
.print V DCSFQCLK|13
.print V DCSFQ_1|2
.print V _TFF|READOUT
.print V DCSFQCLK|2
.print V SUM_TX
.print V _TFF|4
.print V SUM
.print V _TFF|5
.print V CLK_TX
.print V _TFF|TOGGLE
.print V DCSFQ_1|11
.print V DCSFQCLK|8
.print V CBAR_TX
.print V DCSFQ_1|5
.print V DCSFQ_1|6
.print V DCSFQ_1|102
.print V _TFF|SUM_TX
.print V DCSFQCLK|12
.print V DCSFQ_1|8
.print V DCSFQCLK|107
.print V A_TX
.print V DCSFQCLK|102
.print V DCSFQ_1|107
.print V DCSFQ_1|7
.print V DCSFQCLK|6
.print V _TFF|7
.print V CARRY
.print V _TFF|CBAR_TX
.print V DCSFQCLK|1
.print V DCSFQ_1|111
.print V DCSFQCLK|4
.print V _TFF|6
.print V CLK
.print V DCSFQCLK|105
.print V CBAR
.print V A1_DC
.print V DCSFQ_1|105
.print V DCSFQ_1|9
.print V DCSFQ_1|4
.print V _TFF|CARRY_TX
.print V CARRY_TX
.print V DCSFQCLK|9
.print V DCSFQ_1|3
.print V _TFF|1
.print V _TFF|3
.print V DCSFQ_1|1
.print V DCSFQ_1|13
.print V DCSFQCLK|5
.print V DCSFQCLK|11
.print V DCSFQCLK|7
.print V DCSFQCLK|10
.print V DCSFQCLK|3
.print V A
.print V CLK_DC
.print V DCSFQ_1|10
.print V _TFF|2
.print V DCSFQ_1|12
.print DEVP BDCSFQCLK|1
.print DEVP BDCSFQCLK|2
.print DEVP BDCSFQCLK|3
.print DEVP BDCSFQCLK|4
.print DEVP BDCSFQ_1|1
.print DEVP BDCSFQ_1|2
.print DEVP BDCSFQ_1|3
.print DEVP BDCSFQ_1|4
.print DEVP B_TFF|11
.print DEVP B_TFF|10
.print DEVP B_TFF|12
.print DEVP B_TFF|6
.print DEVP B_TFF|1
.print DEVP B_TFF|2
.print DEVP B_TFF|5
.print DEVP B_TFF|4
.print DEVP B_TFF|3
.print DEVP B_TFF|_READOUT|1
.print DEVP B_TFF|_READOUT|2
.print DEVP B_TFF|_READOUT|3
.print DEVP B_TFF|_TOGGLE|1
.print DEVP B_TFF|_TOGGLE|2
.print DEVP B_TFF|_TOGGLE|3
.print DEVP B_TFF|_SUM|1
.print DEVP B_TFF|_SUM|2
.print DEVP B_TFF|_CARRY|1
.print DEVP B_TFF|_CARRY|2
.print DEVP B_TFF|_CBAR|1
.print DEVP B_TFF|_CBAR|2
