
* .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.subckt LSMITLL_JTL a q BiasScale=1
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2
  .param Lsheet=1.13e-12
  .param LP=0.2p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.7

  .param B1=IC
  .param B2=IC
  .param IB1=(B1+B2)*Ic0*BiasCoef
  .param LB1=LB
  .param L1=Phi0/(4*B1*Ic0)
  .param L2=Phi0/(4*B1*Ic0)
  .param L3=Phi0/(4*B1*Ic0)
  .param L4=Phi0/(4*B2*Ic0)
  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param LRB1=(RB1/Rsheet)*Lsheet+LP
  .param LRB2=(RB2/Rsheet)*Lsheet+LP
  .param LP1=LP
  .param LP2=LP

  B1 1 2 jjmit area=B1
  B2 6 7 jjmit area=B2
  IB1 0 5 pwl(0 0 5p IB1*BiasScale)
  L1 a 1 L1
  L2 1 4 L2
  L3 4 6 L3
  L4 6 q L4
  LP1 2 0 LP1
  LP2 7 0 LP2
  LB1 5 4 LB1
  RB1 1 3 RB1
  RB2 6 8 RB2
  LRB1 3 0 LRB1
  LRB2 8 0 LRB2
.ends

.subckt LSmitll_XOR	a	b	clk 	q
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2
  .param Lsheet=1.13e-12
  .param LP=0.5p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.70
  .param B1=IC
  .param B2=IC
  .param B3=IC
  .param B4=B1
  .param B5=B2
  .param B6=B3
  .param B7=IC/1.25
  .param B8=IC
  .param B9=IC/1.25
  .param B10=IC
  .param B11=IC
  .param IB1=BiasCoef*Ic0*B1
  .param IB2=BiasCoef*Ic0*B2
  .param IB3=IB1
  .param IB4=IB2
  .param IB5=BiasCoef*Ic0*B8
  .param IB6=BiasCoef*Ic0*B11
  .param L1=Phi0/(4*IC*Ic0)
  .param L2=Phi0/(2*B1*Ic0)
  .param L3=1.2p
  .param L4=Phi0/(B2*Ic0)
  .param L5=L1
  .param L6=L2
  .param L7=L3
  .param L8=L4
  .param L9=1.2p
  .param L10=Phi0/(4*IC*Ic0)
  .param L11=Phi0/(2*B8*Ic0)
  .param L12=Phi0/(2*B10*Ic0)
  .param L13=Phi0/(4*IC*Ic0)
  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3
  .param RB4=B0Rs/B4
  .param RB5=B0Rs/B5
  .param RB6=B0Rs/B6
  .param RB7=B0Rs/B7
  .param RB8=B0Rs/B8
  .param RB9=B0Rs/B9
  .param RB10=B0Rs/B10
  .param RB11=B0Rs/B11
  .param LRB1=(RB1/Rsheet)*Lsheet+LP
  .param LRB2=(RB2/Rsheet)*Lsheet+LP
  .param LRB3=(RB3/Rsheet)*Lsheet+LP
  .param LRB4=(RB4/Rsheet)*Lsheet+LP
  .param LRB5=(RB5/Rsheet)*Lsheet+LP
  .param LRB6=(RB6/Rsheet)*Lsheet+LP
  .param LRB7=(RB7/Rsheet)*Lsheet+LP
  .param LRB8=(RB8/Rsheet)*Lsheet+LP
  .param LRB9=(RB9/Rsheet)*Lsheet+LP
  .param LRB10=(RB10/Rsheet)*Lsheet+LP
  .param LRB11=(RB11/Rsheet)*Lsheet+LP
  B1 1 2 jjmit area=B1
  B2 4 5 jjmit area=B2
  B3 25 6 jjmit area=B3
  B4 9 10 jjmit area=B4
  B5 12 13 jjmit area=B5
  B6 26 14 jjmit area=B6
  B7 27 16 jjmit area=B7
  B8 17 18 jjmit area=B8
  B9 20 16 jjmit area=B9
  B10 16 21 jjmit area=B10
  B11 22 23 jjmit area=B11
  IB1 0 3 pwl(0 0 5p IB1)
  IB2 0 7 pwl(0 0 5p IB2)
  IB3 0 11 pwl(0 0 5p IB3)
  IB4 0 15 pwl(0 0 5p IB4)
  IB5 0 19 pwl(0 0 5p IB5)
  IB6 0 24 pwl(0 0 5p IB6)
  LB1 3 1 LB
  LB2 7 6 LB
  LB3 11 9 LB
  LB4 15 14 LB
  LB5 19 17 LB
  LB6 24 22 LB
  L1 a 1 L1
  L2 1 4 L2
  L3 4 25 L3
  L4 6 8 L4
  L5 b 9 L5
  L6 9 12 L6
  L7 12 26 L7
  L8 14 8 L8
  L9 8 27 L9
  L10 clk 17 L10
  L11 17 20 L11
  L12 16 22 L12
  L13 22 q L13
  LP1 2 0 LP
  LP2 5 0 LP
  LP4 10 0 LP
  LP5 13 0 LP
  LP8 18 0 LP
  LP10 21 0 LP
  LP11 23 0 LP
  RB1 1 101 RB1
  LRB1 101 0 LRB1
  RB2 4 104 RB2
  LRB2 104 0 LRB2
  RB3 4 106 RB3
  LRB3 106 6 LRB3
  RB4 9 109 RB4
  LRB4 109 0 LRB4
  RB5 12 112 RB5
  LRB5 112 0 LRB5
  RB6 12 114 RB6
  LRB6 114 14 LRB6
  RB7 8 108 RB7
  LRB7 108 16 LRB7
  RB8 17 117 RB8
  LRB8 117 0 LRB8
  RB9 20 120 RB9
  LRB9 120 16 LRB9
  RB10 16 116 RB10
  LRB10 116 0 LRB10
  RB11 22 122 RB11
  LRB11 122 0 LRB11
.ends

.subckt LSMITLL_NOT a clk q BiasScale=1
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2
  .param Lsheet=1.13e-12
  .param LP=0.2p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.7

  .param B1=IC
  .param B2=IC
  .param B3=IC/1.4
  .param B4=IC
  .param B5=IC/1.4
  .param B6=IC
  .param B7=IC/1.4
  .param B8=IC
  .param B9=IC

  .param IB1=BiasCoef*Ic0*B1
  .param IB2=0.5*Ic0*B2
  .param IB3=BiasCoef*Ic0*B6
  .param IB4=BiasCoef*Ic0*B4
  .param IB5=BiasCoef*Ic0*B9

  .param LB1=LB
  .param LB2=LB
  .param LB3=LB
  .param LB4=LB
  .param LB5=LB

  .param L1=Phi0/(4*IC*Ic0)
  .param L2=Phi0/(2*B1*Ic0)
  .param L3=Phi0/(2*B2*Ic0)
  .param L4=Phi0/(4*IC*Ic0)
  .param L5=1p
  .param L6=Phi0/(2*B4*Ic0)
  .param L7=2p
  .param L8=1p
  .param L9=Phi0/(B6*Ic0)
  .param L10=1p
  .param L11=Phi0/(2*B8*Ic0)
  .param L12=Phi0/(4*IC*Ic0)

  .param LP1=LP
  .param LP2=LP
  .param LP4=LP
  .param LP6=LP
  .param LP8=LP
  .param LP9=LP

  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3
  .param RB4=B0Rs/B4
  .param RB5=B0Rs/B5
  .param RB6=B0Rs/B6
  .param RB7=B0Rs/B7
  .param RB8=B0Rs/B8
  .param RB9=B0Rs/B9

  .param LRB1=(RB1/Rsheet)*Lsheet
  .param LRB2=(RB2/Rsheet)*Lsheet
  .param LRB3=(RB3/Rsheet)*Lsheet
  .param LRB4=(RB4/Rsheet)*Lsheet
  .param LRB5=(RB5/Rsheet)*Lsheet
  .param LRB6=(RB6/Rsheet)*Lsheet
  .param LRB7=(RB7/Rsheet)*Lsheet
  .param LRB8=(RB8/Rsheet)*Lsheet
  .param LRB9=(RB9/Rsheet)*Lsheet

  .param RD=4
  .param LRD=2p

  B1 1 2 jjmit area=B1
  B2 4 5 jjmit area=B2
  B3 7 8 jjmit area=B3
  B4 13 14 jjmit area=B4
  B5 17 18 jjmit area=B5
  B6 10 11 jjmit area=B6
  B7 20 18 jjmit area=B7
  B8 18 19 jjmit area=B8
  B9 21 22 jjmit area=B9

  IB1 0 3 pwl(0 0 5p IB1*BiasScale)
  IB2 0 6 pwl(0 0 5p IB2*BiasScale)
  IB3 0 9 pwl(0 0 5p IB3*BiasScale)
  IB4 0 15 pwl(0 0 5p IB4*BiasScale)
  IB5 0 23 pwl(0 0 5p IB5*BiasScale)

  LB1 3 1 LB1
  LB2 6 4 LB2
  LB3 8 9 LB3
  LB4 13 15 LB4
  LB5 21 23 LB5

  L1 a 1 L1
  L2 1 4 L2
  L3 4 7 L3
  L4 clk 13 L4
  L5 13 16 L5
  L6 16 17 L6
  L7 16 12 L7
  L8 10 12 L8
  L9 10 8 L9
  L10 8 20 L10
  L11 18 21 L11
  L12 21 q L12

  LP1 2 0 LP1
  LP2 5 0 LP2
  LP4 14 0 LP4
  LP6 11 0 LP6
  LP8 19 0 LP8
  LP9 22 0 LP9

  RB1 1 101 RB1
  LRB1 101 0 LRB1
  RB2 4 104 RB2
  LRB2 104 5 LRB2
  RB3 7 107 RB3
  LRB3 107 8 LRB3
  RB4 13 113 RB4
  LRB4 113 0 LRB4
  RB5 17 117 RB5
  LRB5 117 18 LRB5
  RB6 10 110 RB6
  LRB6 110 0 LRB6
  RB7 20 120 RB7
  LRB7 120 18 LRB7
  RB8 18 118 RB8
  LRB8 118 0 LRB8
  RB9 21 121 RB9
  LRB9 121 0 LRB9
  LRD 12 112 LRD
  RD 112 0 RD
.ends

.subckt LSmitll_XOR_opt	a	b	clk 	q   BiasScale=1
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2
  .param Lsheet=1.13e-12
  .param LP=0.5p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.70
  .param B1=2.5
  .param B2=2.09
  .param B3=1.71
  .param B4=B1
  .param B5=B2
  .param B6=B3
  .param B7=1.62
  .param B8=2.5
  .param B9=1.45
  .param B10=0.89
  .param B11=2.5
  .param IB1=175u
  .param IB2=112u
  .param IB3=IB1
  .param IB4=IB2
  .param IB5=175u
  .param IB6=175u
  .param L1=Phi0/(4*IC*Ic0)
  .param L2=Phi0/(2*B1*Ic0)
  .param L3=1.2p
  .param L4=Phi0/(B2*Ic0)
  .param L5=L1
  .param L6=L2
  .param L7=L3
  .param L8=L4
  .param L9=1.2p
  .param L10=Phi0/(4*IC*Ic0)
  .param L11=Phi0/(2*B8*Ic0)
  .param L12=Phi0/(2*B10*Ic0)
  .param L13=Phi0/(4*IC*Ic0)
  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3
  .param RB4=B0Rs/B4
  .param RB5=B0Rs/B5
  .param RB6=B0Rs/B6
  .param RB7=B0Rs/B7
  .param RB8=B0Rs/B8
  .param RB9=B0Rs/B9
  .param RB10=B0Rs/B10
  .param RB11=B0Rs/B11
  .param LRB1=(RB1/Rsheet)*Lsheet+LP
  .param LRB2=(RB2/Rsheet)*Lsheet+LP
  .param LRB3=(RB3/Rsheet)*Lsheet+LP
  .param LRB4=(RB4/Rsheet)*Lsheet+LP
  .param LRB5=(RB5/Rsheet)*Lsheet+LP
  .param LRB6=(RB6/Rsheet)*Lsheet+LP
  .param LRB7=(RB7/Rsheet)*Lsheet+LP
  .param LRB8=(RB8/Rsheet)*Lsheet+LP
  .param LRB9=(RB9/Rsheet)*Lsheet+LP
  .param LRB10=(RB10/Rsheet)*Lsheet+LP
  .param LRB11=(RB11/Rsheet)*Lsheet+LP
  B1 1 2 jjmit area=B1
  B2 4 5 jjmit area=B2
  B3 25 6 jjmit area=B3
  B4 9 10 jjmit area=B4
  B5 12 13 jjmit area=B5
  B6 26 14 jjmit area=B6
  B7 27 16 jjmit area=B7
  B8 17 18 jjmit area=B8
  B9 20 16 jjmit area=B9
  B10 16 21 jjmit area=B10
  B11 22 23 jjmit area=B11
  IB1 0 3 pwl(0 0 5p IB1*BiasScale)
  IB2 0 7 pwl(0 0 5p IB2*BiasScale)
  IB3 0 11 pwl(0 0 5p IB3*BiasScale)
  IB4 0 15 pwl(0 0 5p IB4*BiasScale)
  IB5 0 19 pwl(0 0 5p IB5*BiasScale)
  IB6 0 24 pwl(0 0 5p IB6*BiasScale)
  LB1 3 1 LB
  LB2 7 6 LB
  LB3 11 9 LB
  LB4 15 14 LB
  LB5 19 17 LB
  LB6 24 22 LB
  L1 a 1 2.06E-12
  L2 1 4 3.233E-12
  L3 4 25 1.419E-12
  L4 6 8 6.051E-12
  L5 b 9 2.092E-12
  L6 9 12 3.221E-12
  L7 12 26 1.384E-12
  L8 14 8 6.059E-12
  L9 8 27 1.301E-12
  L10 clk 17 2.082E-12
  L11 17 20 1.43E-12
  L12 16 22 3.892E-12
  L13 22 q 2.077E-12
  LP1 2 0 5.508E-13
  LP2 5 0 4.769E-13
  LP4 10 0 4.767E-13
  LP5 13 0 4.812E-13
  LP8 18 0 4.526E-13
  LP10 21 0 5.69E-13
  LP11 23 0 4.746E-13
  RB1 1 101 RB1
  LRB1 101 0 LRB1
  RB2 4 104 RB2
  LRB2 104 0 LRB2
  RB3 4 106 RB3
  LRB3 106 6 LRB3
  RB4 9 109 RB4
  LRB4 109 0 LRB4
  RB5 12 112 RB5
  LRB5 112 0 LRB5
  RB6 12 114 RB6
  LRB6 114 14 LRB6
  RB7 8 108 RB7
  LRB7 108 16 LRB7
  RB8 17 117 RB8
  LRB8 117 0 LRB8
  RB9 20 120 RB9
  LRB9 120 16 LRB9
  RB10 16 116 RB10
  LRB10 116 0 LRB10
  RB11 22 122 RB11
  LRB11 122 0 LRB11
.ends

.subckt LSMITLL_NOT_opt a clk q BiasScale=1
  .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2
  .param Lsheet=1.13e-12
  .param LP=0.2p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.7

  .param B1=IC
  .param B2=2.57
  .param B3=1.07
  .param B4=IC
  .param B5=1.34
  .param B6=3.03
  .param B7=1.38
  .param B8=0.8
  .param B9=IC

  .param IB1=BiasCoef*Ic0*B1
  .param IB2=87u
  .param IB3=257u
  .param IB4=BiasCoef*Ic0*B4
  .param IB5=BiasCoef*Ic0*B9

  .param LB1=LB
  .param LB2=LB
  .param LB3=LB
  .param LB4=LB
  .param LB5=LB

  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3
  .param RB4=B0Rs/B4
  .param RB5=B0Rs/B5
  .param RB6=B0Rs/B6
  .param RB7=B0Rs/B7
  .param RB8=B0Rs/B8
  .param RB9=B0Rs/B9

  .param LRB1=(RB1/Rsheet)*Lsheet
  .param LRB2=(RB2/Rsheet)*Lsheet
  .param LRB3=(RB3/Rsheet)*Lsheet
  .param LRB4=(RB4/Rsheet)*Lsheet
  .param LRB5=(RB5/Rsheet)*Lsheet
  .param LRB6=(RB6/Rsheet)*Lsheet
  .param LRB7=(RB7/Rsheet)*Lsheet
  .param LRB8=(RB8/Rsheet)*Lsheet
  .param LRB9=(RB9/Rsheet)*Lsheet

  .param RD=4
  .param LRD=2p

  B1 1 2 jjmit area=B1
  B2 4 5 jjmit area=B2
  B3 7 8 jjmit area=B3
  B4 13 14 jjmit area=B4
  B5 17 18 jjmit area=B5
  B6 10 11 jjmit area=B6
  B7 20 18 jjmit area=B7
  B8 18 19 jjmit area=B8
  B9 21 22 jjmit area=B9

  IB1 0 3 pwl(0 0 5p IB1*BiasScale)
  IB2 0 6 pwl(0 0 5p IB2*BiasScale)
  IB3 0 9 pwl(0 0 5p IB3*BiasScale)
  IB4 0 15 pwl(0 0 5p IB4*BiasScale)
  IB5 0 23 pwl(0 0 5p IB5*BiasScale)

  LB1 3 1 LB1
  LB2 6 4 LB2
  LB3 8 9 LB3
  LB4 13 15 LB4
  LB5 21 23 LB5

  L1 a 1 2.062E-12
  L2 1 4 1.889E-12
  L3 4 7 2.72E-12
  L4 clk 13 2.057E-12
  L5 13 16 1.029E-12
  L6 16 17 1.241E-12
  L7 16 12 1.973E-12
  L8 10 12 1.003E-12
  L9 10 8 7.524E-12
  L10 8 20 1.234E-12
  L11 18 21 2.607E-12
  L12 21 q 2.062E-12

  LP1 2 0 5.271E-13
  LP2 5 0 5.237E-13
  LP4 14 0 4.759E-13
  LP6 11 0 5.021E-13
  LP8 19 0 6.33E-13
  LP9 22 0 4.749E-13

  RB1 1 101 RB1
  LRB1 101 0 LRB1
  RB2 4 104 RB2
  LRB2 104 5 LRB2
  RB3 7 107 RB3
  LRB3 107 8 LRB3
  RB4 13 113 RB4
  LRB4 113 0 LRB4
  RB5 17 117 RB5
  LRB5 117 18 LRB5
  RB6 10 110 RB6
  LRB6 110 0 LRB6
  RB7 20 120 RB7
  LRB7 120 18 LRB7
  RB8 18 118 RB8
  LRB8 118 0 LRB8
  RB9 21 121 RB9
  LRB9 121 0 LRB9
  LRD 12 112 LRD
  RD 112 0 RD
.ends

.subckt LSMITLL_AND_opt a b clk q
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2 
  .param Lsheet=1.13e-12 
  .param LP=0.2p
  .param IC=2.5
  .param Lptl=2p
  .param LB=2p
  .param BiasCoef=0.7

  .param B1=IC
  .param B2=2.01
  .param B3=1.91
  .param B4=1.26
  .param B5=1.57
  .param B6=1.19
  .param B7=B1
  .param B8=B2
  .param B9=B3
  .param B10=B4
  .param B11=B5
  .param B12=B6
  .param B13=IC
  .param B14=2.06
  .param B15=IC

  .param IB1=BiasCoef*Ic0*B1
  .param IB2=123u
  .param IB3=IB1
  .param IB4=IB2
  .param IB5=BiasCoef*Ic0*B13
  .param IB6=133u
  .param IB7=BiasCoef*Ic0*B15

  .param LB1=LB
  .param LB2=LB
  .param LB3=LB
  .param LB4=LB
  .param LB5=LB
  .param LB6=LB
  .param LB7=LB

  .param L1=Phi0/(4*IC*Ic0)
  .param L2=Phi0/(2*B1*Ic0)
  .param L3=Phi0/(B3*Ic0)
  .param L4=1p
  .param L5=Phi0/(2*B5*Ic0)
  .param L6=L1
  .param L7=L2
  .param L8=L3
  .param L9=L4
  .param L10=L5
  .param L11=Phi0/(4*IC*Ic0)
  .param L12=Phi0/(2*B13*Ic0)
  .param L13=1p
  .param L14=1p
  .param L15=Phi0/(4*IC*Ic0)

  .param LP1=LP
  .param LP3=LP
  .param LP5=LP
  .param LP7=LP
  .param LP9=LP
  .param LP11=LP
  .param LP13=LP
  .param LP14=LP
  .param LP15=LP

  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3
  .param RB4=B0Rs/B4
  .param RB5=B0Rs/B5
  .param RB6=B0Rs/B6
  .param RB7=B0Rs/B7
  .param RB8=B0Rs/B8
  .param RB9=B0Rs/B9
  .param RB10=B0Rs/B10
  .param RB11=B0Rs/B11
  .param RB12=B0Rs/B12
  .param RB13=B0Rs/B13
  .param RB14=B0Rs/B14
  .param RB15=B0Rs/B15
  .param LRB1=(RB1/Rsheet)*Lsheet
  .param LRB2=(RB2/Rsheet)*Lsheet
  .param LRB3=(RB3/Rsheet)*Lsheet
  .param LRB4=(RB4/Rsheet)*Lsheet
  .param LRB5=(RB5/Rsheet)*Lsheet
  .param LRB6=(RB6/Rsheet)*Lsheet
  .param LRB7=(RB7/Rsheet)*Lsheet
  .param LRB8=(RB8/Rsheet)*Lsheet
  .param LRB9=(RB9/Rsheet)*Lsheet
  .param LRB10=(RB10/Rsheet)*Lsheet
  .param LRB11=(RB11/Rsheet)*Lsheet
  .param LRB12=(RB12/Rsheet)*Lsheet
  .param LRB13=(RB13/Rsheet)*Lsheet
  .param LRB14=(RB14/Rsheet)*Lsheet
  .param LRB15=(RB15/Rsheet)*Lsheet

  B1 1 2 jjmit area=B1
  B2 4 5 jjmit area=B2
  B3 5 6 jjmit area=B3
  B4 8 9 jjmit area=B4
  B5 8 11 jjmit area=B5
  B6 12 13 jjmit area=B6
  B7 14 15 jjmit area=B7
  B8 17 18 jjmit area=B8
  B9 18 19 jjmit area=B9
  B10 21 22 jjmit area=B10
  B11 21 23 jjmit area=B11
  B12 24 13 jjmit area=B12
  B13 25 26 jjmit area=B13
  B14 31 32 jjmit area=B14
  B15 28 29 jjmit area=B15

  IB1 0 3 pwl(0 0 5p IB1)
  IB2 0 7 pwl(0 0 5p IB2)
  IB3 0 16 pwl(0 0 5p IB3)
  IB4 0 20 pwl(0 0 5p IB4)
  IB5 0 27 pwl(0 0 5p IB5)
  IB6 0 33 pwl(0 0 5p IB6)
  IB7 0 30 pwl(0 0 5p IB7)

  LB1 3 1 LB1
  LB2 7 5 LB2
  LB3 16 14 LB3
  LB4 20 18 LB4
  LB5 27 25 LB5
  LB6 30 28 LB6
  LB7 33 31 LB7

  LP1 2 0 4.864E-13
  LP3 6 0 5.474E-13
  LP5 11 0 5.279E-13
  LP7 15 0 4.901E-13
  LP9 19 0 5.414E-13
  LP11 23 0 5.306E-13
  LP13 26 0 5.084E-13
  LP14 32 0 5.329E-13
  LP15 29 0 4.92E-13

  L1 a 1 2.075E-12
  L2 1 4 2.812E-12
  L3 5 8 9.756E-12
  L4 9 10 1.079E-12
  L5 8 12 3.105E-12
  L6 b 14 2.073E-12
  L7 14 17 2.811E-12
  L8 18 21 9.768E-12
  L9 22 10 1.084E-12
  L10 21 24 3.095E-12
  L11 clk 25 2.063E-12
  L12 25 31 2.96E-12
  L13 31 10 1.002E-12
  L14 13 28 1.06E-12
  L15 28 q 2.069E-12

  RB1 1 101 RB1
  LRB1 101 0 LRB1
  RB2 4 104 RB2
  LRB2 104 5 LRB2
  RB3 5 105 RB3
  LRB3 105 0 LRB3
  RB4 8 109 RB4
  LRB4 109 9 LRB4
  RB5 8 108 RB5
  LRB5 108 0 LRB5
  RB6 12 112 RB6
  LRB6 112 13 LRB6
  RB7 14 114 RB7
  LRB7 114 0 LRB7
  RB8 17 117 RB8
  LRB8 117 18 LRB8
  RB9 18 118 RB9
  LRB9 118 0 LRB9
  RB10 21 122 RB10
  LRB10 122 22 LRB10
  RB11 21 121 RB11
  LRB11 121 0 LRB11
  RB12 24 124 RB12
  LRB12 124 13 LRB12
  RB13 25 125 RB13
  LRB13 125 0 LRB13
  RB14 31 131 RB14
  LRB14 131 0 LRB14
  RB15 28 128 RB15
  LRB15 128 0 LRB15
.ends

.subckt LSMITLL_AND2 a b clk q
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.2p
    .param IC=2.5
    .param LB=2p
    .param BiasCoef=0.7

    .param B1=IC
    .param B2=IC/1.4
    .param B3=IC
    .param B4=IC/1.4
    .param B5=IC
    .param B6=IC/1.4
    .param B7=B1
    .param B8=B2
    .param B9=B3
    .param B10=B4
    .param B11=B5
    .param B12=B6
    .param B13=IC
    .param B14=IC
    .param B15=IC

    .param IB1=BiasCoef*Ic0*B1
    .param IB2=BiasCoef*Ic0*B3
    .param IB3=IB1
    .param IB4=IB2
    .param IB5=BiasCoef*Ic0*B13
    .param IB6=BiasCoef*Ic0*B14
    .param IB7=BiasCoef*Ic0*B15

    .param LB1=LB
    .param LB2=LB
    .param LB3=LB
    .param LB4=LB
    .param LB5=LB
    .param LB6=LB
    .param LB7=LB

    .param L1=Phi0/(4*IC*Ic0)
    .param L2=Phi0/(2*B1*Ic0)
    .param L3=Phi0/(B3*Ic0)
    .param L4=1p
    .param L5=Phi0/(2*B5*Ic0)
    .param L6=L1
    .param L7=L2
    .param L8=L3
    .param L9=L4
    .param L10=L5
    .param L11=Phi0/(4*IC*Ic0)
    .param L12=Phi0/(2*B13*Ic0)
    .param L13=1p
    .param L14=1p
    .param L15=Phi0/(4*IC*Ic0)

    .param LP1=LP
    .param LP3=LP
    .param LP5=LP
    .param LP7=LP
    .param LP9=LP
    .param LP11=LP
    .param LP13=LP
    .param LP14=LP
    .param LP15=LP

    .param RB1=B0Rs/B1
    .param RB2=B0Rs/B2
    .param RB3=B0Rs/B3
    .param RB4=B0Rs/B4
    .param RB5=B0Rs/B5
    .param RB6=B0Rs/B6
    .param RB7=B0Rs/B7
    .param RB8=B0Rs/B8
    .param RB9=B0Rs/B9
    .param RB10=B0Rs/B10
    .param RB11=B0Rs/B11
    .param RB12=B0Rs/B12
    .param RB13=B0Rs/B13
    .param RB14=B0Rs/B14
    .param RB15=B0Rs/B15
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet
    .param LRB3=(RB3/Rsheet)*Lsheet
    .param LRB4=(RB4/Rsheet)*Lsheet
    .param LRB5=(RB5/Rsheet)*Lsheet
    .param LRB6=(RB6/Rsheet)*Lsheet
    .param LRB7=(RB7/Rsheet)*Lsheet
    .param LRB8=(RB8/Rsheet)*Lsheet
    .param LRB9=(RB9/Rsheet)*Lsheet
    .param LRB10=(RB10/Rsheet)*Lsheet
    .param LRB11=(RB11/Rsheet)*Lsheet
    .param LRB12=(RB12/Rsheet)*Lsheet
    .param LRB13=(RB13/Rsheet)*Lsheet
    .param LRB14=(RB14/Rsheet)*Lsheet
    .param LRB15=(RB15/Rsheet)*Lsheet

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 5 6 jjmit area=B3
    B4 8 9 jjmit area=B4
    B5 8 11 jjmit area=B5
    B6 12 13 jjmit area=B6
    B7 14 15 jjmit area=B7
    B8 17 18 jjmit area=B8
    B9 18 19 jjmit area=B9
    B10 21 22 jjmit area=B10
    B11 21 23 jjmit area=B11
    B12 24 13 jjmit area=B12
    B13 25 26 jjmit area=B13
    B14 31 32 jjmit area=B14
    B15 28 29 jjmit area=B15

    IB1 0 3 pwl(0 0 5p IB1)
    IB2 0 7 pwl(0 0 5p IB2)
    IB3 0 16 pwl(0 0 5p IB3)
    IB4 0 20 pwl(0 0 5p IB4)
    IB5 0 27 pwl(0 0 5p IB5)
    IB6 0 33 pwl(0 0 5p IB6)
    IB7 0 30 pwl(0 0 5p IB7)

    LB1 3 1 LB1
    LB2 7 5 LB2
    LB3 16 14 LB3
    LB4 20 18 LB4
    LB5 27 25 LB5
    LB6 30 28 LB6
    LB7 33 31 LB7

    LP1 2 0 LP1
    LP3 6 0 LP3
    LP5 11 0 LP5
    LP7 15 0 LP7
    LP9 19 0 LP9
    LP11 23 0 LP11
    LP13 26 0 LP13
    LP14 32 0 LP14
    LP15 29 0 LP15

    L1 a 1 L1
    L2 1 4 L2
    L3 5 8 L3
    L4 9 10 L4
    L5 8 12 L5
    L6 b 14 L6
    L7 14 17 L7
    L8 18 21 L8
    L9 22 10 L9
    L10 21 24 L10
    L11 clk 25 L11
    L12 25 31 L12
    L13 31 10 L13
    L14 13 28 L14
    L15 28 q L15

    RB1 1 101 RB1
    LRB1 101 0 LRB1
    RB2 4 104 RB2
    LRB2 104 5 LRB2
    RB3 5 105 RB3
    LRB3 105 0 LRB3
    RB4 8 109 RB4
    LRB4 109 9 LRB4
    RB5 8 108 RB5
    LRB5 108 0 LRB5
    RB6 12 112 RB6
    LRB6 112 13 LRB6
    RB7 14 114 RB7
    LRB7 114 0 LRB7
    RB8 17 117 RB8
    LRB8 117 18 LRB8
    RB9 18 118 RB9
    LRB9 118 0 LRB9
    RB10 21 122 RB10
    LRB10 122 22 LRB10
    RB11 21 121 RB11
    LRB11 121 0 LRB11
    RB12 24 124 RB12
    LRB12 124 13 LRB12
    RB13 25 125 RB13
    LRB13 125 0 LRB13
    RB14 31 131 RB14
    LRB14 131 0 LRB14
    RB15 28 128 RB15
    LRB15 128 0 LRB15
.ends

.subckt LSmitll_XOR_2	a	b	clk 	q
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2
  .param Lsheet=1.13e-12
  .param LP=0.5p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.70
  .param B1=IC
  .param B2=IC
  .param B3=IC
  .param B4=B1
  .param B5=B2
  .param B6=B3
  .param B7=IC/1.25
  .param B8=IC
  .param B9=IC/1.25
  .param B10=IC
  .param B11=IC
  .param IB1=BiasCoef*Ic0*B1
  .param IB2=BiasCoef*Ic0*B2
  .param IB3=IB1
  .param IB4=IB2
  .param IB5=BiasCoef*Ic0*B8
  .param IB6=BiasCoef*Ic0*B11
  .param L1=Phi0/(4*IC*Ic0)
  .param L2=Phi0/(2*B1*Ic0)
  .param L3=1.2p
  .param L4=Phi0/(B2*Ic0)
  .param L5=L1
  .param L6=L2
  .param L7=L3
  .param L8=L4
  .param L9=1.2p
  .param L10=Phi0/(4*IC*Ic0)
  .param L11=Phi0/(2*B8*Ic0)
  .param L12=Phi0/(2*B10*Ic0)
  .param L13=Phi0/(4*IC*Ic0)
  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3
  .param RB4=B0Rs/B4
  .param RB5=B0Rs/B5
  .param RB6=B0Rs/B6
  .param RB7=B0Rs/B7
  .param RB8=B0Rs/B8
  .param RB9=B0Rs/B9
  .param RB10=B0Rs/B10
  .param RB11=B0Rs/B11
  .param LRB1=(RB1/Rsheet)*Lsheet+LP
  .param LRB2=(RB2/Rsheet)*Lsheet+LP
  .param LRB3=(RB3/Rsheet)*Lsheet+LP
  .param LRB4=(RB4/Rsheet)*Lsheet+LP
  .param LRB5=(RB5/Rsheet)*Lsheet+LP
  .param LRB6=(RB6/Rsheet)*Lsheet+LP
  .param LRB7=(RB7/Rsheet)*Lsheet+LP
  .param LRB8=(RB8/Rsheet)*Lsheet+LP
  .param LRB9=(RB9/Rsheet)*Lsheet+LP
  .param LRB10=(RB10/Rsheet)*Lsheet+LP
  .param LRB11=(RB11/Rsheet)*Lsheet+LP
  B1 1 2 jjmit area=B1
  B2 4 5 jjmit area=B2
  B3 25 6 jjmit area=B3
  B4 9 10 jjmit area=B4
  B5 12 13 jjmit area=B5
  B6 26 14 jjmit area=B6
  B7 27 16 jjmit area=B7
  B8 17 18 jjmit area=B8
  B9 20 16 jjmit area=B9
  B10 16 21 jjmit area=B10
  B11 22 23 jjmit area=B11
  IB1 0 3 pwl(0 0 5p IB1)
  IB2 0 7 pwl(0 0 5p IB2)
  IB3 0 11 pwl(0 0 5p IB3)
  IB4 0 15 pwl(0 0 5p IB4)
  IB5 0 19 pwl(0 0 5p IB5)
  IB6 0 24 pwl(0 0 5p IB6)
  LB1 3 1 LB
  LB2 7 6 LB
  LB3 11 9 LB
  LB4 15 14 LB
  LB5 19 17 LB
  LB6 24 22 LB
  L1 a 1 L1
  L2 1 4 L2
  L3 4 25 L3
  L4 6 8 L4
  L5 b 9 L5
  L6 9 12 L6
  L7 12 26 L7
  L8 14 8 L8
  L9 8 27 L9
  L10 clk 17 L10
  L11 17 20 L11
  L12 16 22 L12
  L13 22 q L13
  LP1 2 0 LP
  LP2 5 0 LP
  LP4 10 0 LP
  LP5 13 0 LP
  LP8 18 0 LP
  LP10 21 0 LP
  LP11 23 0 LP
  RB1 1 101 RB1
  LRB1 101 0 LRB1
  RB2 4 104 RB2
  LRB2 104 0 LRB2
  RB3 4 106 RB3
  LRB3 106 6 LRB3
  RB4 9 109 RB4
  LRB4 109 0 LRB4
  RB5 12 112 RB5
  LRB5 112 0 LRB5
  RB6 12 114 RB6
  LRB6 114 14 LRB6
  RB7 8 108 RB7
  LRB7 108 16 LRB7
  RB8 17 117 RB8
  LRB8 117 0 LRB8
  RB9 20 120 RB9
  LRB9 120 16 LRB9
  RB10 16 116 RB10
  LRB10 116 0 LRB10
  RB11 22 122 RB11
  LRB11 122 0 LRB11
.ends

.subckt LSMITLL_BUFF a q
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.5p
    .param IC=2.5
    .param Lptl=2p
    .param LB=2p
    .param BiasCoef=0.7

    .param B1=IC
    .param B2=IC
    .param B3=IC
    .param B4=IC
    .param IB1=B1*Ic0*BiasCoef
    .param IB2=B2*Ic0*0.95
    .param IB3=B3*Ic0*0.95
    .param IB4=B4*Ic0*BiasCoef
    .param LB1=LB
    .param LB2=LB
    .param LB3=LB
    .param LB4=LB
    .param L1=Phi0/(4*IC*Ic0)
    .param L2=Phi0/(2*B1*Ic0)
    .param L3=Phi0/(2*B2*Ic0)
    .param L4=Phi0/(2*B3*Ic0)
    .param L5=Phi0/(4*IC*Ic0)
    .param RB1=B0Rs/B1   
    .param RB2=B0Rs/B2
    .param RB3=B0Rs/B3
    .param RB4=B0Rs/B4
    .param LRB1=(RB1/Rsheet)*Lsheet+LP
    .param LRB2=(RB2/Rsheet)*Lsheet+LP
    .param LRB3=(RB3/Rsheet)*Lsheet+LP
    .param LRB4=(RB4/Rsheet)*Lsheet+LP
    .param LP1=LP
    .param LP2=LP
    .param LP3=LP
    .param LP4=LP

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 7 8 jjmit area=B3
    B4 10 11 jjmit area=B4

    IB1 0 3 pwl(0 0 5p IB1)
    IB2 0 6 pwl(0 0 5p IB2)
    IB3 0 9 pwl(0 0 5p IB3)
    IB4 0 12 pwl(0 0 5p IB4)

    L1 a 1 L1
    L2 1 4 L2
    L3 4 7 L3
    L4 7 10 L4
    L5 10 q L5

    LP1 2 0 LP1
    LP2 5 0 LP2
    LP3 8 0 LP3
    LP4 11 0 LP4

    LB1 1 3 LB1
    LB2 4 6 LB2
    LB3 7 9 LB3
    LB4 10 12 LB4

    RB1 1 101 RB1
    RB2 4 104 RB2
    RB3 7 107 RB3
    RB4 10 110 RB4

    LRB1 101 0 LRB1
    LRB2 104 0 LRB2
    LRB3 107 0 LRB3
    LRB4 110 0 LRB4
.ends


*$Ports a q0 q1
.subckt LSmitll_SPLIT a q0 q1
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.2p
    .param IC=2.5
    .param Lptl=2p
    .param LB=2p
    .param BiasCoef=0.7
    .param RD=1.36

    .param B1=IC
    .param B2=1.4*IC
    .param B3=IC
    .param B4=IC

    .param IB1=BiasCoef*Ic0*B1
    .param IB2=BiasCoef*Ic0*B2
    .param IB3=BiasCoef*Ic0*B3
    .param IB4=IB3

    .param L1=Lptl
    .param L2=Phi0/(2*B1*Ic0)
    .param L3=(Phi0/(2*B2*Ic0))/2
    .param L4=L3
    .param L5=Lptl
    .param L6=L3
    .param L7=Lptl

    .param RB1=B0Rs/B1
    .param RB2=B0Rs/B2
    .param RB3=B0Rs/B3
    .param RB4=B0Rs/B4
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet
    .param LRB3=(RB3/Rsheet)*Lsheet
    .param LRB4=(RB4/Rsheet)*Lsheet

    IB1 0 3 pwl(0 0 5p IB1)
    IB2 0 6 pwl(0 0 5p IB2)
    IB3 0 10 pwl(0 0 5p IB3)
    IB4 0 13 pwl(0 0 5p IB4)
    LB1 3 1 LB
    LB2 6 4 LB
    LB3 10 8 LB
    LB4 13 11 LB

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 8 9 jjmit area=B3
    B4 11 12 jjmit area=B4
    L1 a 1 L1
    L2 1 4 L2
    L3 4 7 L3
    L4 7 8 L4
    L5 8 q0 L5
    L6 7 11 L6
    L7 11 q1 L7

    LP1 2 0 0.2p
    LP2 5 0 0.2p
    LP3 9 0 0.2p
    LP4 12 0 0.2p
    RB1 1 101 RB1
    LRB1 101 0 LRB1
    RB2 4 104 RB2
    LRB2 104 0 LRB2
    RB3 8 108 RB3
    LRB3 108 0 LRB3
    RB4 11 111 RB4
    LRB4 111 0 LRB4
.ends

.subckt LSmitll_DFF_opt	  a	clk q	BiasScale=1
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.2p
    .param IC=2.5
    .param LB=2p
    .param BiasCoef=0.70

    .param B1=2.5
    .param B2=1.61
    .param B3=1.54
    .param B4=1.69
    .param B5=1.38
    .param B6=2.5
    .param B7=2.5

    .param IB1=175u     
    .param IB2=173u      
    .param IB3=175u            
    .param IB4=175u        

    .param L1=Phi0/(4*IC*Ic0)               
    .param L2=Phi0/(2*B1*Ic0)         
    .param L3=Phi0/(B3*Ic0)       
    .param L4=Phi0/(2*B6*Ic0)      
    .param L5=Phi0/(4*IC*Ic0)     
    .param L6=Phi0/(2*B4*Ic0)       
    .param L7=Phi0/(4*B7*Ic0)         
    .param LB1=LB            
    .param LB2=LB           
    .param LB3=LB           
    .param LB4=LB        
    .param LP1=LP         
    .param LP3=LP          
    .param LP4=LP         
    .param LP6=LP          
    .param LP7=LP          
    .param RB1=B0Rs/B1       
    .param RB2=B0Rs/B2       
    .param RB3=B0Rs/B3          
    .param RB4=B0Rs/B4         
    .param RB5=B0Rs/B5         
    .param RB6=B0Rs/B6          
    .param RB7=B0Rs/B7
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet
    .param LRB3=(RB3/Rsheet)*Lsheet
    .param LRB4=(RB4/Rsheet)*Lsheet
    .param LRB5=(RB5/Rsheet)*Lsheet
    .param LRB6=(RB6/Rsheet)*Lsheet
    .param LRB7=(RB7/Rsheet)*Lsheet

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 5 6 jjmit area=B3
    B4 8 9 jjmit area=B4
    B5 10 8 jjmit area=B5
    B6 11 12 jjmit area=B6
    B7 14 15 jjmit area=B7

    IB1 0 3 pwl(0 0 5p IB1*BiasScale)
    IB2 0 7 pwl(0 0 5p IB2*BiasScale)
    IB3 0 13 pwl(0 0 5p IB3*BiasScale)
    IB4 0 16 pwl(0 0 5p IB4*BiasScale)

    LB1 3 1 LB1
    LB2 7 5 LB2
    LB3 11 13 LB3
    LB4 16 14 LB4

    L1 a 1 2.059E-12
    L2 1 4 4.123E-12
    L3 5 8 6.873E-12
    L4 10 11 5.195E-12
    L5 clk 11 2.071E-12
    L6 8 14 3.287E-12
    L7 14 q 2.066E-12

    LP1 2 0 5.042E-13    
    LP3 6 0 5.799E-13    
    LP4 9 0 5.733E-13    
    LP6 12 0 4.605E-13    
    LP7 15 0 4.961E-13    

    RB1 1 101 RB1
    LRB1 101 0 LRB1
    RB2 4 104 RB2
    LRB2 104 5 LRB2
    RB3 5 105 RB3
    LRB3 105 0 LRB3
    RB4 8 108 RB4
    LRB4 108 0 LRB4
    RB5 10 110 RB5
    LRB5 110 8 LRB5
    RB6 11 111 RB6
    LRB6 111 0 LRB6
    RB7 14 114 RB7
    LRB7 114 0 LRB7
.ends

.subckt LSmitll_MERGE_opt a b q mbias=1 BiasScale=1
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.2p
    .param IC=2.5
    .param LB=2p
    .param BiasCoef=0.70
    .param RD=1.36

    .param B1=IC
    .param B2=2.5
    .param B3=1.92
    .param B4=B1
    .param B5=B2
    .param B6=B3
    .param B7=2.53
    .param B8=IC

    .param IB1=BiasCoef*Ic0*B1
    .param IB2=IB1
    .param IB3=254E-6
    .param IB4=192E-6
    .param IB5=BiasCoef*Ic0*B8

    .param L1=Phi0/(4*IC*Ic0)
    .param L2=3.173E-12
    .param L3=1.2E-12
    .param L4=L1
    .param L5=L2
    .param L6=L3
    .param L7=5.354E-12
    .param L8=4.456E-12
    .param L9=Phi0/(4*B8*Ic0)

    .param LB1=LB
    .param LB2=LB
    .param LB3=LB
    .param LB4=LB
    .param LB5=LB

    .param LP1=LP
    .param LP2=LP
    .param LP4=LP
    .param LP5=LP
    .param LP7=LP
    .param LP8=LP

    .param RB1=B0Rs/B1
    .param RB2=B0Rs/B2
    .param RB3=B0Rs/B3
    .param RB4=B0Rs/B4
    .param RB5=B0Rs/B5
    .param RB6=B0Rs/B6
    .param RB7=B0Rs/B7
    .param RB8=B0Rs/B8
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet
    .param LRB3=(RB3/Rsheet)*Lsheet
    .param LRB4=(RB4/Rsheet)*Lsheet
    .param LRB5=(RB5/Rsheet)*Lsheet
    .param LRB6=(RB6/Rsheet)*Lsheet
    .param LRB7=(RB7/Rsheet)*Lsheet
    .param LRB8=(RB8/Rsheet)*Lsheet

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 4 6 jjmit area=B3
    B4 8 9 jjmit area=B4
    B5 11 12 jjmit area=B5
    B6 11 13 jjmit area=B6
    B7 15 16 jjmit area=B7
    B8 18 19 jjmit area=B8

    IB1 0 3 pwl(0 0 5p IB1*BiasScale)
    IB2 0 10 pwl(0 0 5p IB2*BiasScale)
    IB3 0 14 pwl(0 0 5p IB3*mbias*BiasScale)
    IB4 0 17 pwl(0 0 5p IB4*BiasScale)
    IB5 0 20 pwl(0 0 5p IB5*BiasScale)

    L1 a 1 2.117E-12
    L2 1 4 3.17E-12
    L3 6 7 1.234E-12

    L4 b 8 2.082E-12
    L5 8 11 3.165E-12
    L6 13 7 1.224E-12

    L7 7 15 5.299E-12
    L8 15 18 4.489E-12
    L9 18 q 2.077E-12

    LP1 2 0 4.652E-13
    LP2 5 0 4.457E-13
    LP4 9 0 5.293E-13
    LP5 12 0 4.452E-13
    LP7 16 0 5.039E-13
    LP8 19 0 4.984E-13

    LB1 1 3 LB1
    LB2 8 10 LB2
    LB3 7 14 LB3
    LB4 15 17 LB4
    LB5 18 20 LB5

    RB1 1 101 RB1
    LRB1 101 0 LRB1
    RB2 4 104 RB2
    LRB2 104 0 LRB2
    RB3 4 106 RB3
    LRB3 106 6 LRB3
    RB4 8 108 RB4
    LRB4 108 0 LRB4
    RB5 11 111 RB5
    LRB5 111 0 LRB5
    RB6 11 113 RB6
    LRB6 113 13 LRB6
    RB7 15 115 RB7
    LRB7 115 0 LRB7
    RB8 18 118 RB8
    LRB8 118 0 LRB8
.ends

.subckt LSmitll_SPLIT_opt a q0 q1 BiasScale=1
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.2p
    .param IC=2.5
    .param Lptl=2p
    .param LB=2p
    .param BiasCoef=0.7
    .param RD=1.36

    .param B1=2.5
    .param B2=3.0
    .param B3=2.5
    .param B4=2.5

    .param IB1=175u
    .param IB2=280u
    .param IB3=175u
    .param IB4=175u

    .param L1=Lptl
    .param L2=Phi0/(2*B1*Ic0)
    .param L3=(Phi0/(2*B2*Ic0))/2
    .param L4=L3
    .param L5=Lptl
    .param L6=L3
    .param L7=Lptl

    .param RB1=B0Rs/B1
    .param RB2=B0Rs/B2
    .param RB3=B0Rs/B3
    .param RB4=B0Rs/B4
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet
    .param LRB3=(RB3/Rsheet)*Lsheet
    .param LRB4=(RB4/Rsheet)*Lsheet

    IB1 0 3 pwl(0 0 5p IB1*BiasScale)
    IB2 0 6 pwl(0 0 5p IB2*BiasScale)
    IB3 0 10 pwl(0 0 5p IB3*BiasScale)
    IB4 0 13 pwl(0 0 5p IB4*BiasScale)
    LB1 3 1 9.175E-13
    LB2 6 4 7.666E-13
    LB3 10 8 1.928E-12
    LB4 13 11 8.786E-13

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 8 9 jjmit area=B3
    B4 11 12 jjmit area=B4
    L1 a 1 2.063E-12
    L2 1 4 3.637E-12
    L3 4 7 1.278E-12
    L4 7 8 1.305E-12
    L5 8 q0 2.05E-12
    L6 7 11 1.315E-12
    L7 11 q1 2.06E-12

    LP1 2 0 4.676E-13
    LP2 5 0 4.498E-13
    LP3 9 0 5.183E-13
    LP4 12 0 4.639E-13
    RB1 1 101 RB1
    LRB1 101 0 LRB1
    RB2 4 104 RB2
    LRB2 104 0 LRB2
    RB3 8 108 RB3
    LRB3 108 0 LRB3
    RB4 11 111 RB4
    LRB4 111 0 LRB4
.ends

.subckt LSmitll_PTLTX a q
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.5p
    .param LB=2p
    .param Lptl=2p
    .param RD=1.36
    .param IC=2.5
    .param BiasCoef=0.7

    .param B1=IC
    .param B2=IC
    .param IB1=BiasCoef*Ic0*B1      
    .param IB2=BiasCoef*Ic0*B2
    .param L1=Phi0/(4*B1*Ic0)         
    .param L2=Phi0/(2*B1*Ic0)     
    .param L3=Lptl
    .param LB1=LB           
    .param LB2=LB   
    .param LP1=LP         
    .param LP2=LP 
    .param RB1=B0Rs/B1       
    .param RB2=B0Rs/B2   
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    IB1 0 3 pwl(0 0 5p IB1)
    IB2 0 6 pwl(0 0 5p IB2)
    LB1 1 3 1.684E-012
    LB2 4 6 3.596E-012
    L1 a 1 2.063E-012
    L2 1 4 4.123E-012
    L3 4 7 2.193E-012
    RD 7 q RD
    LP1 2 0 5.254E-013
    LP2 5 0 5.141E-013
    RB1 1 101 RB1
    RB2 4 104 RB2
    LRB1 101 0 LRB1
    LRB2 104 0 LRB2
.ends

.subckt LSmitll_PTLRX a q
    .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
    .param Phi0=2.067833848E-15
    .param B0=1
    .param Ic0=0.0001
    .param IcRs=100u*6.859904418
    .param B0Rs=IcRs/Ic0*B0
    .param Rsheet=2 
    .param Lsheet=1.13e-12 
    .param LP=0.5p
    .param LB=2p
    .param Lptl=2p
    .param IC=2.5
    .param BiasCoef=0.7

    .param B1=IC/1.54
    .param B2=IC/1.25
    .param B3=IC
    .param IB1=Ic0*B1
    .param IB2=BiasCoef*Ic0*B2
    .param IB3=BiasCoef*Ic0*B3
    .param L1=Lptl
    .param L2=Phi0/(2*B1*Ic0)
    .param L3=Phi0/(2*B2*Ic0)
    .param L4=Phi0/(4*IC*Ic0)

    .param LB1=LB
    .param LB2=LB
    .param LB3=LB
    .param LP1=LP         
    .param LP2=LP          
    .param LP3=LP  
    .param RB1=B0Rs/B1       
    .param RB2=B0Rs/B2       
    .param RB3=B0Rs/B3   
    .param LRB1=(RB1/Rsheet)*Lsheet
    .param LRB2=(RB2/Rsheet)*Lsheet
    .param LRB3=(RB3/Rsheet)*Lsheet

    B1 1 2 jjmit area=B1
    B2 4 5 jjmit area=B2
    B3 7 8 jjmit area=B3
    IB1 0 3 pwl(0 0 5p IB1)
    LB1 1 3 2.777E-012
    IB2 0 6 pwl(0 0 5p IB2)
    LB2 4 6 2.685E-012
    IB3 0 9 pwl(0 0 5p IB3)
    LB3 7 9 2.764E-012
    L1 a 1 1.346E-012
    L2 1 4 6.348E-012
    L3 4 7 5.197E-012
    L4 7 q 2.058E-012

    LP1 2 0 4.795E-013
    LP2 5 0 5.431E-013
    LP3 8 0 5.339E-013
    RB1 1 101 RB1
    RB2 4 104 RB2
    RB3 7 107 RB3
    LRB1 101 0 LRB1
    LRB2 104 0 LRB2
    LRB3 107 0 LRB3
.ends

.subckt LSMITLL_DCSFQ a q
  .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
  .param Phi0=2.067833848E-15
  .param B0=1
  .param Ic0=0.0001
  .param IcRs=100u*6.859904418
  .param B0Rs=IcRs/Ic0*B0
  .param Rsheet=2 
  .param Lsheet=1.13e-12 
  .param LP=0.5p
  .param IC=2.5
  .param LB=2p
  .param BiasCoef=0.7

  .param B1=2.25
  .param B2=2.25
  .param B3=IC

  .param IB1=275u/1.4
  .param IB2=B3*Ic0*BiasCoef

  .param LB1=LB
  .param LB2=LB

  .param L1=1p
  .param L2=3.9p
  .param L3=0.6p
  .param L4=1.1p
  .param L5=4.5p
  .param L6=Phi0/(4*IC*Ic0)

  .param LP2=LP
  .param LP3=LP

  .param RB1=B0Rs/B1
  .param RB2=B0Rs/B2
  .param RB3=B0Rs/B3

  .param LRB1=(RB1/Rsheet)*Lsheet
  .param LRB2=(RB2/Rsheet)*Lsheet+LP
  .param LRB3=(RB3/Rsheet)*Lsheet+LP

  * Input
  L1 a 1 L1
  L2 1 0 L2 
  L3 1 2 L3 

  B1 2 3 jjmit  area=B1 
  RB1 2 102 RB1  
  LRB1 102 3 LRB1 

  L4 3 5 L4 

  * grounded
  B2 5 6 jjmit  area=B2 
  LP2 6 0 LP2 
  RB2 5 105 RB2  
  LRB2 105 0 LRB2 

  L5 5 7 L5 

  * grounded
  B3 7 8 jjmit  area=B3 
  LP3 8 0 LP3 
  RB3 7 107 RB3  
  LRB3 107 0 LRB3

  IB1 0 4 pwl(0 0 5p IB1)
  LB1 4 3 LB1 
  IB2 0 9 pwl(0 0 5p IB2)
  LB2 9 7 LB2 

  L6 7 q L6 


.ends