*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PRINT DEVI ROUT_936C
.PRINT DEVI I33CC
.PRINT DEVI I5F5F
.PRINT V 33CC
.PRINT V 5F5F
.PRINT V 6C93
.PRINT V 936C
.PRINT DEVI IT1
.PRINT DEVI IT2
.TRAN 1E-12 8.250000000000001E-09
ROUT_936C 936C 0  1
I33CC 0 33CC  PWL(0 0 2.97E-10 0 3E-10 0.0005 3.03E-10 0 7.97E-10 0 8E-10 0.0005 8.03E-10 0 1.297E-09 0 1.3E-09 0.0005 1.303E-09 0 1.797E-09 0 1.8E-09 0.0005 1.803E-09 0 2.297E-09 0 2.3E-09 0.0005 2.303E-09 0 2.797E-09 0 2.8E-09 0.0005 2.803E-09 0 3.297E-09 0 3.3E-09 0.0005 3.303E-09 0 3.797E-09 0 3.8E-09 0.0005 3.803E-09 0 4.297E-09 0 4.3E-09 0.0005 4.303E-09 0 4.797E-09 0 4.8E-09 0.0005 4.803E-09 0 5.297E-09 0 5.3E-09 0.0005 5.303E-09 0 5.797E-09 0 5.8E-09 0.0005 5.803E-09 0 6.297E-09 0 6.3E-09 0.0005 6.303E-09 0 6.797E-09 0 6.8E-09 0.0005 6.803E-09 0 7.297E-09 0 7.3E-09 0.0005 7.303E-09 0 7.797E-09 0 7.8E-09 0.0005 7.803E-09 0)
I5F5F 0 5F5F  PWL(0 0 5.97E-10 0 6E-10 0.0005 6.03E-10 0 8.47E-10 0 8.5E-10 0.0005 8.53E-10 0 1.597E-09 0 1.6E-09 0.0005 1.603E-09 0 1.847E-09 0 1.85E-09 0.0005 1.853E-09 0 2.597E-09 0 2.6E-09 0.0005 2.603E-09 0 2.847E-09 0 2.85E-09 0.0005 2.853E-09 0 3.597E-09 0 3.6E-09 0.0005 3.603E-09 0 3.847E-09 0 3.85E-09 0.0005 3.853E-09 0 4.597E-09 0 4.6E-09 0.0005 4.603E-09 0 4.847E-09 0 4.85E-09 0.0005 4.853E-09 0 5.597E-09 0 5.6E-09 0.0005 5.603E-09 0 5.847E-09 0 5.85E-09 0.0005 5.853E-09 0 6.597E-09 0 6.6E-09 0.0005 6.603E-09 0 6.847E-09 0 6.85E-09 0.0005 6.853E-09 0 7.597E-09 0 7.6E-09 0.0005 7.603E-09 0 7.847E-09 0 7.85E-09 0.0005 7.853E-09 0)
IT1 0 T1  PWL(0 0  2.4700000000000003E-10 0 2.5E-10 0.0005 2.53E-10 0 4.97E-10 0 5E-10 0.0005 5.03E-10 0 7.470000000000001E-10 0 7.500000000000001E-10 0.0005 7.530000000000001E-10 0 9.97E-10 0 1E-09 0.0005 1.0030000000000002E-09 0 1.247E-09 0 1.25E-09 0.0005 1.2530000000000001E-09 0 1.4970000000000001E-09 0 1.5000000000000002E-09 0.0005 1.5030000000000003E-09 0 1.747E-09 0 1.7500000000000002E-09 0.0005 1.7530000000000003E-09 0 1.997E-09 0 2E-09 0.0005 2.0030000000000002E-09 0 2.247E-09 0 2.2500000000000003E-09 0.0005 2.2530000000000004E-09 0 2.497E-09 0 2.5E-09 0.0005 2.503E-09 0 2.747E-09 0 2.7500000000000002E-09 0.0005 2.7530000000000003E-09 0 2.9970000000000003E-09 0 3.0000000000000004E-09 0.0005 3.0030000000000005E-09 0 3.247E-09 0 3.25E-09 0.0005 3.2530000000000002E-09 0 3.4970000000000002E-09 0 3.5000000000000003E-09 0.0005 3.5030000000000004E-09 0 3.747E-09 0 3.7500000000000005E-09 0.0005 3.7530000000000006E-09 0 3.997E-09 0 4E-09 0.0005 4.003E-09 0 4.247E-09 0 4.25E-09 0.0005 4.253E-09 0 4.4970000000000005E-09 0 4.500000000000001E-09 0.0005 4.503000000000001E-09 0 4.747E-09 0 4.75E-09 0.0005 4.7530000000000004E-09 0 4.997E-09 0 5E-09 0.0005 5.003E-09 0 5.247000000000001E-09 0 5.250000000000001E-09 0.0005 5.253000000000001E-09 0 5.497E-09 0 5.5000000000000004E-09 0.0005 5.5030000000000005E-09 0 5.747E-09 0 5.75E-09 0.0005 5.753E-09 0 5.997000000000001E-09 0 6.000000000000001E-09 0.0005 6.003000000000001E-09 0 6.2470000000000005E-09 0 6.2500000000000005E-09 0.0005 6.253000000000001E-09 0 6.497E-09 0 6.5E-09 0.0005 6.503E-09 0 6.747E-09 0 6.75E-09 0.0005 6.753E-09 0 6.9970000000000005E-09 0 7.000000000000001E-09 0.0005 7.003000000000001E-09 0 7.247E-09 0 7.25E-09 0.0005 7.2530000000000005E-09 0 7.497000000000001E-09 0 7.500000000000001E-09 0.0005 7.503000000000001E-09 0 7.747E-09 0 7.75E-09 0.0005 7.753E-09 0 7.997E-09 0 8E-09 0.0005 8.003E-09 0 )
IT2 0 T2  PWL(0 0  2.4700000000000003E-10 0 2.5E-10 0.0005 2.53E-10 0 4.97E-10 0 5E-10 0.0005 5.03E-10 0 7.470000000000001E-10 0 7.500000000000001E-10 0.0005 7.530000000000001E-10 0 9.97E-10 0 1E-09 0.0005 1.0030000000000002E-09 0 1.247E-09 0 1.25E-09 0.0005 1.2530000000000001E-09 0 1.4970000000000001E-09 0 1.5000000000000002E-09 0.0005 1.5030000000000003E-09 0 1.747E-09 0 1.7500000000000002E-09 0.0005 1.7530000000000003E-09 0 1.997E-09 0 2E-09 0.0005 2.0030000000000002E-09 0 2.247E-09 0 2.2500000000000003E-09 0.0005 2.2530000000000004E-09 0 2.497E-09 0 2.5E-09 0.0005 2.503E-09 0 2.747E-09 0 2.7500000000000002E-09 0.0005 2.7530000000000003E-09 0 2.9970000000000003E-09 0 3.0000000000000004E-09 0.0005 3.0030000000000005E-09 0 3.247E-09 0 3.25E-09 0.0005 3.2530000000000002E-09 0 3.4970000000000002E-09 0 3.5000000000000003E-09 0.0005 3.5030000000000004E-09 0 3.747E-09 0 3.7500000000000005E-09 0.0005 3.7530000000000006E-09 0 3.997E-09 0 4E-09 0.0005 4.003E-09 0 4.247E-09 0 4.25E-09 0.0005 4.253E-09 0 4.4970000000000005E-09 0 4.500000000000001E-09 0.0005 4.503000000000001E-09 0 4.747E-09 0 4.75E-09 0.0005 4.7530000000000004E-09 0 4.997E-09 0 5E-09 0.0005 5.003E-09 0 5.247000000000001E-09 0 5.250000000000001E-09 0.0005 5.253000000000001E-09 0 5.497E-09 0 5.5000000000000004E-09 0.0005 5.5030000000000005E-09 0 5.747E-09 0 5.75E-09 0.0005 5.753E-09 0 5.997000000000001E-09 0 6.000000000000001E-09 0.0005 6.003000000000001E-09 0 6.2470000000000005E-09 0 6.2500000000000005E-09 0.0005 6.253000000000001E-09 0 6.497E-09 0 6.5E-09 0.0005 6.503E-09 0 6.747E-09 0 6.75E-09 0.0005 6.753E-09 0 6.9970000000000005E-09 0 7.000000000000001E-09 0.0005 7.003000000000001E-09 0 7.247E-09 0 7.25E-09 0.0005 7.2530000000000005E-09 0 7.497000000000001E-09 0 7.500000000000001E-09 0.0005 7.503000000000001E-09 0 7.747E-09 0 7.75E-09 0.0005 7.753E-09 0 7.997E-09 0 8E-09 0.0005 8.003E-09 0 )
L6C93|A1 33CC 6C93|A1  2.067833848e-12
L6C93|A2 6C93|A1 6C93|A2  4.135667696e-12
L6C93|A3 6C93|A3 6C93|AB  8.271335392e-12
L6C93|B1 5F5F 6C93|B1  2.067833848e-12
L6C93|B2 6C93|B1 6C93|B2  4.135667696e-12
L6C93|B3 6C93|B3 6C93|AB  8.271335392e-12
L6C93|T1 T1 6C93|T1  2.067833848e-12
L6C93|T2 6C93|T1 6C93|T2  4.135667696e-12
L6C93|Q2 6C93|ABTQ 6C93|Q1  4.135667696e-12
L6C93|Q1 6C93|Q1 6C93_O  2.067833848e-12
LJTL1|1 6C93_O JTL1|1  2.067833848e-12
LJTL1|2 JTL1|1 JTL1|4  2.067833848e-12
LJTL1|3 JTL1|4 JTL1|6  2.067833848e-12
LJTL1|4 JTL1|6 6C93_1  2.067833848e-12
LJTL2|1 6C93_1 JTL2|1  2.067833848e-12
LJTL2|2 JTL2|1 JTL2|4  2.067833848e-12
LJTL2|3 JTL2|4 JTL2|6  2.067833848e-12
LJTL2|4 JTL2|6 6C93_2  2.067833848e-12
LJTL3|1 6C93_2 JTL3|1  2.067833848e-12
LJTL3|2 JTL3|1 JTL3|4  2.067833848e-12
LJTL3|3 JTL3|4 JTL3|6  2.067833848e-12
LJTL3|4 JTL3|6 6C93_3  2.067833848e-12
LJTL4|1 6C93_3 JTL4|1  2.067833848e-12
LJTL4|2 JTL4|1 JTL4|4  2.067833848e-12
LJTL4|3 JTL4|4 JTL4|6  2.067833848e-12
LJTL4|4 JTL4|6 6C93_I  2.067833848e-12
L936C|1 6C93_I 936C|A1  2.067833848e-12
L936C|2 936C|A1 936C|A2  4.135667696e-12
L936C|3 936C|A2 936C|A3  4.135667696e-12
L936C|4 T2 936C|T1  2.067833848e-12
L936C|5 936C|T1 936C|T2  1e-12
L936C|7 936C|T2 936C|CW1  2e-12
L936C|8 936C|CW1 936C|CW2  1e-12
L936C|9 936C|CW2 936C|A4  8.271335392e-12
L936C|10 936C|A4 936C|CW3  1e-12
L936C|6 936C|T2 936C|CCW  4.135667696e-12
L936C|11 936C|Q2 936C|Q1  4.135667696e-12
L936C|12 936C|Q1 936C  2.067833848e-12
L936C|RD 936C|CW1 936C|112  2e-12
R936C|D 936C|112 0  4
L6C93|I_A1|B 6C93|A1 6C93|I_A1|MID  2e-12
I6C93|I_A1|B 0 6C93|I_A1|MID  0.000175
L6C93|I_A3|B 6C93|A3 6C93|I_A3|MID  2e-12
I6C93|I_A3|B 0 6C93|I_A3|MID  0.000175
L6C93|I_B1|B 6C93|B1 6C93|I_B1|MID  2e-12
I6C93|I_B1|B 0 6C93|I_B1|MID  0.000175
L6C93|I_B3|B 6C93|B3 6C93|I_B3|MID  2e-12
I6C93|I_B3|B 0 6C93|I_B3|MID  0.000175
L6C93|I_T1|B 6C93|T1 6C93|I_T1|MID  2e-12
I6C93|I_T1|B 0 6C93|I_T1|MID  0.000175
L6C93|I_Q1|B 6C93|Q1 6C93|I_Q1|MID  2e-12
I6C93|I_Q1|B 0 6C93|I_Q1|MID  0.000175
B6C93|A1|1 6C93|A1 6C93|A1|MID_SERIES JJMIT AREA=2.5
L6C93|A1|P 6C93|A1|MID_SERIES 0  5e-13
R6C93|A1|B 6C93|A1 6C93|A1|MID_SHUNT  2.7439617672
L6C93|A1|RB 6C93|A1|MID_SHUNT 0  2.050338398468e-12
B6C93|A2|1 6C93|A2 6C93|A2|MID_SERIES JJMIT AREA=2.5
L6C93|A2|P 6C93|A2|MID_SERIES 0  5e-13
R6C93|A2|B 6C93|A2 6C93|A2|MID_SHUNT  2.7439617672
L6C93|A2|RB 6C93|A2|MID_SHUNT 0  2.050338398468e-12
B6C93|A3|1 6C93|A2 6C93|A3|MID_SERIES JJMIT AREA=2.5
L6C93|A3|P 6C93|A3|MID_SERIES 6C93|A3  1.2e-12
R6C93|A3|B 6C93|A2 6C93|A3|MID_SHUNT  2.7439617672
L6C93|A3|RB 6C93|A3|MID_SHUNT 6C93|A3  2.050338398468e-12
B6C93|B1|1 6C93|B1 6C93|B1|MID_SERIES JJMIT AREA=2.5
L6C93|B1|P 6C93|B1|MID_SERIES 0  5e-13
R6C93|B1|B 6C93|B1 6C93|B1|MID_SHUNT  2.7439617672
L6C93|B1|RB 6C93|B1|MID_SHUNT 0  2.050338398468e-12
B6C93|B2|1 6C93|B2 6C93|B2|MID_SERIES JJMIT AREA=2.5
L6C93|B2|P 6C93|B2|MID_SERIES 0  5e-13
R6C93|B2|B 6C93|B2 6C93|B2|MID_SHUNT  2.7439617672
L6C93|B2|RB 6C93|B2|MID_SHUNT 0  2.050338398468e-12
B6C93|B3|1 6C93|B2 6C93|B3|MID_SERIES JJMIT AREA=2.5
L6C93|B3|P 6C93|B3|MID_SERIES 6C93|B3  1.2e-12
R6C93|B3|B 6C93|B2 6C93|B3|MID_SHUNT  2.7439617672
L6C93|B3|RB 6C93|B3|MID_SHUNT 6C93|B3  2.050338398468e-12
B6C93|T1|1 6C93|T1 6C93|T1|MID_SERIES JJMIT AREA=2.5
L6C93|T1|P 6C93|T1|MID_SERIES 0  5e-13
R6C93|T1|B 6C93|T1 6C93|T1|MID_SHUNT  2.7439617672
L6C93|T1|RB 6C93|T1|MID_SHUNT 0  2.050338398468e-12
B6C93|T2|1 6C93|T2 6C93|ABTQ JJMIT AREA=2.0
R6C93|T2|B 6C93|T2 6C93|T2|MID_SHUNT  3.429952209
L6C93|T2|RB 6C93|T2|MID_SHUNT 6C93|ABTQ  2.437922998085e-12
B6C93|AB|1 6C93|AB 6C93|AB|MID_SERIES JJMIT AREA=2.0
L6C93|AB|P 6C93|AB|MID_SERIES 6C93|ABTQ  1.2e-12
R6C93|AB|B 6C93|AB 6C93|AB|MID_SHUNT  3.429952209
L6C93|AB|RB 6C93|AB|MID_SHUNT 6C93|ABTQ  2.437922998085e-12
B6C93|ABTQ|1 6C93|ABTQ 6C93|ABTQ|MID_SERIES JJMIT AREA=2.5
L6C93|ABTQ|P 6C93|ABTQ|MID_SERIES 0  5e-13
R6C93|ABTQ|B 6C93|ABTQ 6C93|ABTQ|MID_SHUNT  2.7439617672
L6C93|ABTQ|RB 6C93|ABTQ|MID_SHUNT 0  2.050338398468e-12
B6C93|Q1|1 6C93|Q1 6C93|Q1|MID_SERIES JJMIT AREA=2.5
L6C93|Q1|P 6C93|Q1|MID_SERIES 0  5e-13
R6C93|Q1|B 6C93|Q1 6C93|Q1|MID_SHUNT  2.7439617672
L6C93|Q1|RB 6C93|Q1|MID_SHUNT 0  2.050338398468e-12
BJTL1|1|1 JTL1|1 JTL1|1|MID_SERIES JJMIT AREA=2.5
LJTL1|1|P JTL1|1|MID_SERIES 0  2e-13
RJTL1|1|B JTL1|1 JTL1|1|MID_SHUNT  2.7439617672
LJTL1|1|RB JTL1|1|MID_SHUNT 0  1.750338398468e-12
LJTL1|B|B JTL1|4 JTL1|B|MID  2e-12
IJTL1|B|B 0 JTL1|B|MID  0.0005
BJTL1|2|1 JTL1|6 JTL1|2|MID_SERIES JJMIT AREA=2.5
LJTL1|2|P JTL1|2|MID_SERIES 0  2e-13
RJTL1|2|B JTL1|6 JTL1|2|MID_SHUNT  2.7439617672
LJTL1|2|RB JTL1|2|MID_SHUNT 0  1.750338398468e-12
BJTL2|1|1 JTL2|1 JTL2|1|MID_SERIES JJMIT AREA=2.5
LJTL2|1|P JTL2|1|MID_SERIES 0  2e-13
RJTL2|1|B JTL2|1 JTL2|1|MID_SHUNT  2.7439617672
LJTL2|1|RB JTL2|1|MID_SHUNT 0  1.750338398468e-12
LJTL2|B|B JTL2|4 JTL2|B|MID  2e-12
IJTL2|B|B 0 JTL2|B|MID  0.0005
BJTL2|2|1 JTL2|6 JTL2|2|MID_SERIES JJMIT AREA=2.5
LJTL2|2|P JTL2|2|MID_SERIES 0  2e-13
RJTL2|2|B JTL2|6 JTL2|2|MID_SHUNT  2.7439617672
LJTL2|2|RB JTL2|2|MID_SHUNT 0  1.750338398468e-12
BJTL3|1|1 JTL3|1 JTL3|1|MID_SERIES JJMIT AREA=2.5
LJTL3|1|P JTL3|1|MID_SERIES 0  2e-13
RJTL3|1|B JTL3|1 JTL3|1|MID_SHUNT  2.7439617672
LJTL3|1|RB JTL3|1|MID_SHUNT 0  1.750338398468e-12
LJTL3|B|B JTL3|4 JTL3|B|MID  2e-12
IJTL3|B|B 0 JTL3|B|MID  0.0005
BJTL3|2|1 JTL3|6 JTL3|2|MID_SERIES JJMIT AREA=2.5
LJTL3|2|P JTL3|2|MID_SERIES 0  2e-13
RJTL3|2|B JTL3|6 JTL3|2|MID_SHUNT  2.7439617672
LJTL3|2|RB JTL3|2|MID_SHUNT 0  1.750338398468e-12
BJTL4|1|1 JTL4|1 JTL4|1|MID_SERIES JJMIT AREA=2.5
LJTL4|1|P JTL4|1|MID_SERIES 0  2e-13
RJTL4|1|B JTL4|1 JTL4|1|MID_SHUNT  2.7439617672
LJTL4|1|RB JTL4|1|MID_SHUNT 0  1.750338398468e-12
LJTL4|B|B JTL4|4 JTL4|B|MID  2e-12
IJTL4|B|B 0 JTL4|B|MID  0.0005
BJTL4|2|1 JTL4|6 JTL4|2|MID_SERIES JJMIT AREA=2.5
LJTL4|2|P JTL4|2|MID_SERIES 0  2e-13
RJTL4|2|B JTL4|6 JTL4|2|MID_SHUNT  2.7439617672
LJTL4|2|RB JTL4|2|MID_SHUNT 0  1.750338398468e-12
B936C|1|1 936C|A1 936C|1|MID_SERIES JJMIT AREA=2.5
L936C|1|P 936C|1|MID_SERIES 0  2e-13
R936C|1|B 936C|A1 936C|1|MID_SHUNT  2.7439617672
L936C|1|RB 936C|1|MID_SHUNT 0  1.550338398468e-12
B936C|2|1 936C|A2 936C|2|B_JCT JJMIT AREA=1.7857142857142858
R936C|2|B 936C|A2 936C|2|MID_SHUNT  3.84154647408
L936C|2|RB 936C|2|MID_SHUNT 936C|2|B_JCT  2.1704737578552e-12
L936C|2|P_SERIES 936C|2|B_JCT 0  2e-13
B936C|3|1 936C|A3 936C|A4 JJMIT AREA=1.7857142857142858
R936C|3|B 936C|A3 936C|3|MID_SHUNT  3.84154647408
L936C|3|RB 936C|3|MID_SHUNT 936C|A4  2.1704737578552e-12
B936C|4|1 936C|T1 936C|4|MID_SERIES JJMIT AREA=2.5
L936C|4|P 936C|4|MID_SERIES 0  2e-13
R936C|4|B 936C|T1 936C|4|MID_SHUNT  2.7439617672
L936C|4|RB 936C|4|MID_SHUNT 0  1.550338398468e-12
B936C|6|1 936C|CW2 936C|6|MID_SERIES JJMIT AREA=2.5
L936C|6|P 936C|6|MID_SERIES 0  2e-13
R936C|6|B 936C|CW2 936C|6|MID_SHUNT  2.7439617672
L936C|6|RB 936C|6|MID_SHUNT 0  1.550338398468e-12
B936C|7|1 936C|CW3 936C|Q2 JJMIT AREA=1.7857142857142858
R936C|7|B 936C|CW3 936C|7|MID_SHUNT  3.84154647408
L936C|7|RB 936C|7|MID_SHUNT 936C|Q2  2.1704737578552e-12
B936C|5|1 936C|CCW 936C|Q2 JJMIT AREA=1.7857142857142858
R936C|5|B 936C|CCW 936C|5|MID_SHUNT  3.84154647408
L936C|5|RB 936C|5|MID_SHUNT 936C|Q2  2.1704737578552e-12
B936C|8|1 936C|Q2 936C|8|MID_SERIES JJMIT AREA=2.5
L936C|8|P 936C|8|MID_SERIES 0  2e-13
R936C|8|B 936C|Q2 936C|8|MID_SHUNT  2.7439617672
L936C|8|RB 936C|8|MID_SHUNT 0  1.550338398468e-12
B936C|9|1 936C|Q1 936C|9|MID_SERIES JJMIT AREA=2.5
L936C|9|P 936C|9|MID_SERIES 0  2e-13
R936C|9|B 936C|Q1 936C|9|MID_SHUNT  2.7439617672
L936C|9|RB 936C|9|MID_SHUNT 0  1.550338398468e-12
L936C|I_A1|B 936C|A1 936C|I_A1|MID  2e-12
I936C|I_A1|B 0 936C|I_A1|MID  0.000175
L936C|I_A2|B 936C|A2 936C|I_A2|MID  2e-12
I936C|I_A2|B 0 936C|I_A2|MID  0.000125
L936C|I_A4|B 936C|A4 936C|I_A4|MID  2e-12
I936C|I_A4|B 0 936C|I_A4|MID  0.000175
L936C|I_T1|B 936C|T1 936C|I_T1|MID  2e-12
I936C|I_T1|B 0 936C|I_T1|MID  0.000175
L936C|I_Q1|B 936C|Q1 936C|I_Q1|MID  2e-12
I936C|I_Q1|B 0 936C|I_Q1|MID  0.000175
