*
.include /Users/brainkz/Documents/GitHub/SFQ_gate_Exploration/jj_library.cir
.include /Users/brainkz/Documents/GitHub/SFQ/sunmagnetics_library.cir

.param offset1=0

.param tclock=10e-11

Xt1       clk  clk_sig    clk_offset=offset1 factor=1    Tck=tclock

Xdata_a1  a  data_signal_a   clk_offset=offset1 do_factor=0.1 Tck=tclock
Xdata_b1  b  data_signal_b   clk_offset=offset1 do_factor=0.7 Tck=tclock
Xdata_c1  c  data_signal_c_r clk_offset=offset1 do_factor=0.4 Tck=tclock

X_merge a      b a_or_b    merge mbias=1
X_xor a_or_b c clk q xor t_scaling=1 main_scaling=1 bottom_scaling=1

ROUT q  0  1  

.tran 0.1e-12 0.45e-09

.end
