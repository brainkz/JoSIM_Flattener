*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM TCLOCK=2e-10
.PARAM OS=1.0000000000000001e-11
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.5E-12 2000E-12
R_S0 S0_5 0  1
R_S1 S1_5 0  1
R_S2 S2_5 0  1
R_S3 S3_5 0  1
R_S4 S4_5 0  1
R_S5 S5_5 0  1
R_S6 S6_5 0  1
R_S7 S7_5 0  1
R_S8 S8_5 0  1
IA0|A 0 A0_TX  PWL(0 0 2.63e-10 0 2.66e-10 0.0007 2.69e-10 0 6.63e-10 0 6.66e-10 0.0007 6.69e-10 0 1.063e-09 0 1.066e-09 0.0007 1.069e-09 0 1.463e-09 0 1.466e-09 0.0007 1.469e-09 0 1.863e-09 0 1.866e-09 0.0007 1.869e-09 0 2.263e-09 0 2.266e-09 0.0007 2.269e-09 0 2.663e-09 0 2.666e-09 0.0007 2.669e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 3.463e-09 0 3.466e-09 0.0007 3.469e-09 0 3.863e-09 0 3.866e-09 0.0007 3.869e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.663e-09 0 4.666e-09 0.0007 4.669e-09 0 5.063e-09 0 5.066e-09 0.0007 5.069e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.863e-09 0 5.866e-09 0.0007 5.869e-09 0 6.263e-09 0 6.266e-09 0.0007 6.269e-09 0 6.663e-09 0 6.666e-09 0.0007 6.669e-09 0 7.063e-09 0 7.066e-09 0.0007 7.069e-09 0 7.463e-09 0 7.466e-09 0.0007 7.469e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 8.263e-09 0 8.266e-09 0.0007 8.269e-09 0 8.663e-09 0 8.666e-09 0.0007 8.669e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.463e-09 0 9.466e-09 0.0007 9.469e-09 0 9.863e-09 0 9.866e-09 0.0007 9.869e-09 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0663e-08 0 1.0666e-08 0.0007 1.0669e-08 0 1.1063e-08 0 1.1066e-08 0.0007 1.1069e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1863e-08 0 1.1866e-08 0.0007 1.1869e-08 0 1.2263e-08 0 1.2266e-08 0.0007 1.2269e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.3063e-08 0 1.3066e-08 0.0007 1.3069e-08 0 1.3463e-08 0 1.3466e-08 0.0007 1.3469e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.4263e-08 0 1.4266e-08 0.0007 1.4269e-08 0 1.4663e-08 0 1.4666e-08 0.0007 1.4669e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5463e-08 0 1.5466e-08 0.0007 1.5469e-08 0 1.5863e-08 0 1.5866e-08 0.0007 1.5869e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6663e-08 0 1.6666e-08 0.0007 1.6669e-08 0 1.7063e-08 0 1.7066e-08 0.0007 1.7069e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7863e-08 0 1.7866e-08 0.0007 1.7869e-08 0 1.8263e-08 0 1.8266e-08 0.0007 1.8269e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.9063e-08 0 1.9066e-08 0.0007 1.9069e-08 0 1.9463e-08 0 1.9466e-08 0.0007 1.9469e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 2.0263e-08 0 2.0266e-08 0.0007 2.0269e-08 0 2.0663e-08 0 2.0666e-08 0.0007 2.0669e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1463e-08 0 2.1466e-08 0.0007 2.1469e-08 0 2.1863e-08 0 2.1866e-08 0.0007 2.1869e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2663e-08 0 2.2666e-08 0.0007 2.2669e-08 0 2.3063e-08 0 2.3066e-08 0.0007 2.3069e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3863e-08 0 2.3866e-08 0.0007 2.3869e-08 0 2.4263e-08 0 2.4266e-08 0.0007 2.4269e-08 0 2.4663e-08 0 2.4666e-08 0.0007 2.4669e-08 0 2.5063e-08 0 2.5066e-08 0.0007 2.5069e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 2.5863e-08 0 2.5866e-08 0.0007 2.5869e-08 0 2.6263e-08 0 2.6266e-08 0.0007 2.6269e-08 0 2.6663e-08 0 2.6666e-08 0.0007 2.6669e-08 0 2.7063e-08 0 2.7066e-08 0.0007 2.7069e-08 0 2.7463e-08 0 2.7466e-08 0.0007 2.7469e-08 0 2.7863e-08 0 2.7866e-08 0.0007 2.7869e-08 0 2.8263e-08 0 2.8266e-08 0.0007 2.8269e-08 0 2.8663e-08 0 2.8666e-08 0.0007 2.8669e-08 0 2.9063e-08 0 2.9066e-08 0.0007 2.9069e-08 0 2.9463e-08 0 2.9466e-08 0.0007 2.9469e-08 0 2.9863e-08 0 2.9866e-08 0.0007 2.9869e-08 0 3.0263e-08 0 3.0266e-08 0.0007 3.0269e-08 0 3.0663e-08 0 3.0666e-08 0.0007 3.0669e-08 0 3.1063e-08 0 3.1066e-08 0.0007 3.1069e-08 0 3.1463e-08 0 3.1466e-08 0.0007 3.1469e-08 0 3.1863e-08 0 3.1866e-08 0.0007 3.1869e-08 0 3.2263e-08 0 3.2266e-08 0.0007 3.2269e-08 0 3.2663e-08 0 3.2666e-08 0.0007 3.2669e-08 0 3.3063e-08 0 3.3066e-08 0.0007 3.3069e-08 0 3.3463e-08 0 3.3466e-08 0.0007 3.3469e-08 0 3.3863e-08 0 3.3866e-08 0.0007 3.3869e-08 0 3.4263e-08 0 3.4266e-08 0.0007 3.4269e-08 0 3.4663e-08 0 3.4666e-08 0.0007 3.4669e-08 0 3.5063e-08 0 3.5066e-08 0.0007 3.5069e-08 0 3.5463e-08 0 3.5466e-08 0.0007 3.5469e-08 0 3.5863e-08 0 3.5866e-08 0.0007 3.5869e-08 0 3.6263e-08 0 3.6266e-08 0.0007 3.6269e-08 0 3.6663e-08 0 3.6666e-08 0.0007 3.6669e-08 0 3.7063e-08 0 3.7066e-08 0.0007 3.7069e-08 0 3.7463e-08 0 3.7466e-08 0.0007 3.7469e-08 0 3.7863e-08 0 3.7866e-08 0.0007 3.7869e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 3.8663e-08 0 3.8666e-08 0.0007 3.8669e-08 0 3.9063e-08 0 3.9066e-08 0.0007 3.9069e-08 0 3.9463e-08 0 3.9466e-08 0.0007 3.9469e-08 0 3.9863e-08 0 3.9866e-08 0.0007 3.9869e-08 0 4.0263e-08 0 4.0266e-08 0.0007 4.0269e-08 0 4.0663e-08 0 4.0666e-08 0.0007 4.0669e-08 0 4.1063e-08 0 4.1066e-08 0.0007 4.1069e-08 0 4.1463e-08 0 4.1466e-08 0.0007 4.1469e-08 0 4.1863e-08 0 4.1866e-08 0.0007 4.1869e-08 0 4.2263e-08 0 4.2266e-08 0.0007 4.2269e-08 0 4.2663e-08 0 4.2666e-08 0.0007 4.2669e-08 0 4.3063e-08 0 4.3066e-08 0.0007 4.3069e-08 0 4.3463e-08 0 4.3466e-08 0.0007 4.3469e-08 0 4.3863e-08 0 4.3866e-08 0.0007 4.3869e-08 0 4.4263e-08 0 4.4266e-08 0.0007 4.4269e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.5063e-08 0 4.5066e-08 0.0007 4.5069e-08 0 4.5463e-08 0 4.5466e-08 0.0007 4.5469e-08 0 4.5863e-08 0 4.5866e-08 0.0007 4.5869e-08 0 4.6263e-08 0 4.6266e-08 0.0007 4.6269e-08 0 4.6663e-08 0 4.6666e-08 0.0007 4.6669e-08 0 4.7063e-08 0 4.7066e-08 0.0007 4.7069e-08 0 4.7463e-08 0 4.7466e-08 0.0007 4.7469e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.8263e-08 0 4.8266e-08 0.0007 4.8269e-08 0 4.8663e-08 0 4.8666e-08 0.0007 4.8669e-08 0 4.9063e-08 0 4.9066e-08 0.0007 4.9069e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 4.9863e-08 0 4.9866e-08 0.0007 4.9869e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA1|B 0 A1_TX  PWL(0 0 4.63e-10 0 4.66e-10 0.0007 4.69e-10 0 6.63e-10 0 6.66e-10 0.0007 6.69e-10 0 1.263e-09 0 1.266e-09 0.0007 1.269e-09 0 1.463e-09 0 1.466e-09 0.0007 1.469e-09 0 2.063e-09 0 2.066e-09 0.0007 2.069e-09 0 2.263e-09 0 2.266e-09 0.0007 2.269e-09 0 2.863e-09 0 2.866e-09 0.0007 2.869e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 3.663e-09 0 3.666e-09 0.0007 3.669e-09 0 3.863e-09 0 3.866e-09 0.0007 3.869e-09 0 4.463e-09 0 4.466e-09 0.0007 4.469e-09 0 4.663e-09 0 4.666e-09 0.0007 4.669e-09 0 5.263e-09 0 5.266e-09 0.0007 5.269e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.263e-09 0 6.266e-09 0.0007 6.269e-09 0 6.863e-09 0 6.866e-09 0.0007 6.869e-09 0 7.063e-09 0 7.066e-09 0.0007 7.069e-09 0 7.663e-09 0 7.666e-09 0.0007 7.669e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.663e-09 0 8.666e-09 0.0007 8.669e-09 0 9.263e-09 0 9.266e-09 0.0007 9.269e-09 0 9.463e-09 0 9.466e-09 0.0007 9.469e-09 0 1.0063e-08 0 1.0066e-08 0.0007 1.0069e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.1063e-08 0 1.1066e-08 0.0007 1.1069e-08 0 1.1663e-08 0 1.1666e-08 0.0007 1.1669e-08 0 1.1863e-08 0 1.1866e-08 0.0007 1.1869e-08 0 1.2463e-08 0 1.2466e-08 0.0007 1.2469e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.3263e-08 0 1.3266e-08 0.0007 1.3269e-08 0 1.3463e-08 0 1.3466e-08 0.0007 1.3469e-08 0 1.4063e-08 0 1.4066e-08 0.0007 1.4069e-08 0 1.4263e-08 0 1.4266e-08 0.0007 1.4269e-08 0 1.4863e-08 0 1.4866e-08 0.0007 1.4869e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5863e-08 0 1.5866e-08 0.0007 1.5869e-08 0 1.6463e-08 0 1.6466e-08 0.0007 1.6469e-08 0 1.6663e-08 0 1.6666e-08 0.0007 1.6669e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.7269e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8263e-08 0 1.8266e-08 0.0007 1.8269e-08 0 1.8863e-08 0 1.8866e-08 0.0007 1.8869e-08 0 1.9063e-08 0 1.9066e-08 0.0007 1.9069e-08 0 1.9663e-08 0 1.9666e-08 0.0007 1.9669e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0663e-08 0 2.0666e-08 0.0007 2.0669e-08 0 2.1263e-08 0 2.1266e-08 0.0007 2.1269e-08 0 2.1463e-08 0 2.1466e-08 0.0007 2.1469e-08 0 2.2063e-08 0 2.2066e-08 0.0007 2.2069e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.3063e-08 0 2.3066e-08 0.0007 2.3069e-08 0 2.3663e-08 0 2.3666e-08 0.0007 2.3669e-08 0 2.3863e-08 0 2.3866e-08 0.0007 2.3869e-08 0 2.4463e-08 0 2.4466e-08 0.0007 2.4469e-08 0 2.4663e-08 0 2.4666e-08 0.0007 2.4669e-08 0 2.5263e-08 0 2.5266e-08 0.0007 2.5269e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 2.6063e-08 0 2.6066e-08 0.0007 2.6069e-08 0 2.6263e-08 0 2.6266e-08 0.0007 2.6269e-08 0 2.6863e-08 0 2.6866e-08 0.0007 2.6869e-08 0 2.7063e-08 0 2.7066e-08 0.0007 2.7069e-08 0 2.7663e-08 0 2.7666e-08 0.0007 2.7669e-08 0 2.7863e-08 0 2.7866e-08 0.0007 2.7869e-08 0 2.8463e-08 0 2.8466e-08 0.0007 2.8469e-08 0 2.8663e-08 0 2.8666e-08 0.0007 2.8669e-08 0 2.9263e-08 0 2.9266e-08 0.0007 2.9269e-08 0 2.9463e-08 0 2.9466e-08 0.0007 2.9469e-08 0 3.0063e-08 0 3.0066e-08 0.0007 3.0069e-08 0 3.0263e-08 0 3.0266e-08 0.0007 3.0269e-08 0 3.0863e-08 0 3.0866e-08 0.0007 3.0869e-08 0 3.1063e-08 0 3.1066e-08 0.0007 3.1069e-08 0 3.1663e-08 0 3.1666e-08 0.0007 3.1669e-08 0 3.1863e-08 0 3.1866e-08 0.0007 3.1869e-08 0 3.2463e-08 0 3.2466e-08 0.0007 3.2469e-08 0 3.2663e-08 0 3.2666e-08 0.0007 3.2669e-08 0 3.3263e-08 0 3.3266e-08 0.0007 3.3269e-08 0 3.3463e-08 0 3.3466e-08 0.0007 3.3469e-08 0 3.4063e-08 0 3.4066e-08 0.0007 3.4069e-08 0 3.4263e-08 0 3.4266e-08 0.0007 3.4269e-08 0 3.4863e-08 0 3.4866e-08 0.0007 3.4869e-08 0 3.5063e-08 0 3.5066e-08 0.0007 3.5069e-08 0 3.5663e-08 0 3.5666e-08 0.0007 3.5669e-08 0 3.5863e-08 0 3.5866e-08 0.0007 3.5869e-08 0 3.6463e-08 0 3.6466e-08 0.0007 3.6469e-08 0 3.6663e-08 0 3.6666e-08 0.0007 3.6669e-08 0 3.7263e-08 0 3.7266e-08 0.0007 3.7269e-08 0 3.7463e-08 0 3.7466e-08 0.0007 3.7469e-08 0 3.8063e-08 0 3.8066e-08 0.0007 3.8069e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 3.8863e-08 0 3.8866e-08 0.0007 3.8869e-08 0 3.9063e-08 0 3.9066e-08 0.0007 3.9069e-08 0 3.9663e-08 0 3.9666e-08 0.0007 3.9669e-08 0 3.9863e-08 0 3.9866e-08 0.0007 3.9869e-08 0 4.0463e-08 0 4.0466e-08 0.0007 4.0469e-08 0 4.0663e-08 0 4.0666e-08 0.0007 4.0669e-08 0 4.1263e-08 0 4.1266e-08 0.0007 4.1269e-08 0 4.1463e-08 0 4.1466e-08 0.0007 4.1469e-08 0 4.2063e-08 0 4.2066e-08 0.0007 4.2069e-08 0 4.2263e-08 0 4.2266e-08 0.0007 4.2269e-08 0 4.2863e-08 0 4.2866e-08 0.0007 4.2869e-08 0 4.3063e-08 0 4.3066e-08 0.0007 4.3069e-08 0 4.3663e-08 0 4.3666e-08 0.0007 4.3669e-08 0 4.3863e-08 0 4.3866e-08 0.0007 4.3869e-08 0 4.4463e-08 0 4.4466e-08 0.0007 4.4469e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.5263e-08 0 4.5266e-08 0.0007 4.5269e-08 0 4.5463e-08 0 4.5466e-08 0.0007 4.5469e-08 0 4.6063e-08 0 4.6066e-08 0.0007 4.6069e-08 0 4.6263e-08 0 4.6266e-08 0.0007 4.6269e-08 0 4.6863e-08 0 4.6866e-08 0.0007 4.6869e-08 0 4.7063e-08 0 4.7066e-08 0.0007 4.7069e-08 0 4.7663e-08 0 4.7666e-08 0.0007 4.7669e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.8463e-08 0 4.8466e-08 0.0007 4.8469e-08 0 4.8663e-08 0 4.8666e-08 0.0007 4.8669e-08 0 4.9263e-08 0 4.9266e-08 0.0007 4.9269e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 5.0063e-08 0 5.0066e-08 0.0007 5.0069e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA2|C 0 A2_TX  PWL(0 0 8.63e-10 0 8.66e-10 0.0007 8.69e-10 0 1.063e-09 0 1.066e-09 0.0007 1.069e-09 0 1.263e-09 0 1.266e-09 0.0007 1.269e-09 0 1.463e-09 0 1.466e-09 0.0007 1.469e-09 0 2.463e-09 0 2.466e-09 0.0007 2.469e-09 0 2.663e-09 0 2.666e-09 0.0007 2.669e-09 0 2.863e-09 0 2.866e-09 0.0007 2.869e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 4.063e-09 0 4.066e-09 0.0007 4.069e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.463e-09 0 4.466e-09 0.0007 4.469e-09 0 4.663e-09 0 4.666e-09 0.0007 4.669e-09 0 5.663e-09 0 5.666e-09 0.0007 5.669e-09 0 5.863e-09 0 5.866e-09 0.0007 5.869e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.263e-09 0 6.266e-09 0.0007 6.269e-09 0 7.263e-09 0 7.266e-09 0.0007 7.269e-09 0 7.463e-09 0 7.466e-09 0.0007 7.469e-09 0 7.663e-09 0 7.666e-09 0.0007 7.669e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 8.863e-09 0 8.866e-09 0.0007 8.869e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.263e-09 0 9.266e-09 0.0007 9.269e-09 0 9.463e-09 0 9.466e-09 0.0007 9.469e-09 0 1.0463e-08 0 1.0466e-08 0.0007 1.0469e-08 0 1.0663e-08 0 1.0666e-08 0.0007 1.0669e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.1063e-08 0 1.1066e-08 0.0007 1.1069e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2263e-08 0 1.2266e-08 0.0007 1.2269e-08 0 1.2463e-08 0 1.2466e-08 0.0007 1.2469e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.3663e-08 0 1.3666e-08 0.0007 1.3669e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.4063e-08 0 1.4066e-08 0.0007 1.4069e-08 0 1.4263e-08 0 1.4266e-08 0.0007 1.4269e-08 0 1.5263e-08 0 1.5266e-08 0.0007 1.5269e-08 0 1.5463e-08 0 1.5466e-08 0.0007 1.5469e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5863e-08 0 1.5866e-08 0.0007 1.5869e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.7063e-08 0 1.7066e-08 0.0007 1.7069e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.7269e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.8463e-08 0 1.8466e-08 0.0007 1.8469e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8863e-08 0 1.8866e-08 0.0007 1.8869e-08 0 1.9063e-08 0 1.9066e-08 0.0007 1.9069e-08 0 2.0063e-08 0 2.0066e-08 0.0007 2.0069e-08 0 2.0263e-08 0 2.0266e-08 0.0007 2.0269e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0663e-08 0 2.0666e-08 0.0007 2.0669e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1863e-08 0 2.1866e-08 0.0007 2.1869e-08 0 2.2063e-08 0 2.2066e-08 0.0007 2.2069e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.3263e-08 0 2.3266e-08 0.0007 2.3269e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3663e-08 0 2.3666e-08 0.0007 2.3669e-08 0 2.3863e-08 0 2.3866e-08 0.0007 2.3869e-08 0 2.4863e-08 0 2.4866e-08 0.0007 2.4869e-08 0 2.5063e-08 0 2.5066e-08 0.0007 2.5069e-08 0 2.5263e-08 0 2.5266e-08 0.0007 2.5269e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 2.6463e-08 0 2.6466e-08 0.0007 2.6469e-08 0 2.6663e-08 0 2.6666e-08 0.0007 2.6669e-08 0 2.6863e-08 0 2.6866e-08 0.0007 2.6869e-08 0 2.7063e-08 0 2.7066e-08 0.0007 2.7069e-08 0 2.8063e-08 0 2.8066e-08 0.0007 2.8069e-08 0 2.8263e-08 0 2.8266e-08 0.0007 2.8269e-08 0 2.8463e-08 0 2.8466e-08 0.0007 2.8469e-08 0 2.8663e-08 0 2.8666e-08 0.0007 2.8669e-08 0 2.9663e-08 0 2.9666e-08 0.0007 2.9669e-08 0 2.9863e-08 0 2.9866e-08 0.0007 2.9869e-08 0 3.0063e-08 0 3.0066e-08 0.0007 3.0069e-08 0 3.0263e-08 0 3.0266e-08 0.0007 3.0269e-08 0 3.1263e-08 0 3.1266e-08 0.0007 3.1269e-08 0 3.1463e-08 0 3.1466e-08 0.0007 3.1469e-08 0 3.1663e-08 0 3.1666e-08 0.0007 3.1669e-08 0 3.1863e-08 0 3.1866e-08 0.0007 3.1869e-08 0 3.2863e-08 0 3.2866e-08 0.0007 3.2869e-08 0 3.3063e-08 0 3.3066e-08 0.0007 3.3069e-08 0 3.3263e-08 0 3.3266e-08 0.0007 3.3269e-08 0 3.3463e-08 0 3.3466e-08 0.0007 3.3469e-08 0 3.4463e-08 0 3.4466e-08 0.0007 3.4469e-08 0 3.4663e-08 0 3.4666e-08 0.0007 3.4669e-08 0 3.4863e-08 0 3.4866e-08 0.0007 3.4869e-08 0 3.5063e-08 0 3.5066e-08 0.0007 3.5069e-08 0 3.6063e-08 0 3.6066e-08 0.0007 3.6069e-08 0 3.6263e-08 0 3.6266e-08 0.0007 3.6269e-08 0 3.6463e-08 0 3.6466e-08 0.0007 3.6469e-08 0 3.6663e-08 0 3.6666e-08 0.0007 3.6669e-08 0 3.7663e-08 0 3.7666e-08 0.0007 3.7669e-08 0 3.7863e-08 0 3.7866e-08 0.0007 3.7869e-08 0 3.8063e-08 0 3.8066e-08 0.0007 3.8069e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 3.9263e-08 0 3.9266e-08 0.0007 3.9269e-08 0 3.9463e-08 0 3.9466e-08 0.0007 3.9469e-08 0 3.9663e-08 0 3.9666e-08 0.0007 3.9669e-08 0 3.9863e-08 0 3.9866e-08 0.0007 3.9869e-08 0 4.0863e-08 0 4.0866e-08 0.0007 4.0869e-08 0 4.1063e-08 0 4.1066e-08 0.0007 4.1069e-08 0 4.1263e-08 0 4.1266e-08 0.0007 4.1269e-08 0 4.1463e-08 0 4.1466e-08 0.0007 4.1469e-08 0 4.2463e-08 0 4.2466e-08 0.0007 4.2469e-08 0 4.2663e-08 0 4.2666e-08 0.0007 4.2669e-08 0 4.2863e-08 0 4.2866e-08 0.0007 4.2869e-08 0 4.3063e-08 0 4.3066e-08 0.0007 4.3069e-08 0 4.4063e-08 0 4.4066e-08 0.0007 4.4069e-08 0 4.4263e-08 0 4.4266e-08 0.0007 4.4269e-08 0 4.4463e-08 0 4.4466e-08 0.0007 4.4469e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.5663e-08 0 4.5666e-08 0.0007 4.5669e-08 0 4.5863e-08 0 4.5866e-08 0.0007 4.5869e-08 0 4.6063e-08 0 4.6066e-08 0.0007 4.6069e-08 0 4.6263e-08 0 4.6266e-08 0.0007 4.6269e-08 0 4.7263e-08 0 4.7266e-08 0.0007 4.7269e-08 0 4.7463e-08 0 4.7466e-08 0.0007 4.7469e-08 0 4.7663e-08 0 4.7666e-08 0.0007 4.7669e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.8863e-08 0 4.8866e-08 0.0007 4.8869e-08 0 4.9063e-08 0 4.9066e-08 0.0007 4.9069e-08 0 4.9263e-08 0 4.9266e-08 0.0007 4.9269e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 5.0463e-08 0 5.0466e-08 0.0007 5.0469e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA3|D 0 A3_TX  PWL(0 0 1.663e-09 0 1.666e-09 0.0007 1.669e-09 0 1.863e-09 0 1.866e-09 0.0007 1.869e-09 0 2.063e-09 0 2.066e-09 0.0007 2.069e-09 0 2.263e-09 0 2.266e-09 0.0007 2.269e-09 0 2.463e-09 0 2.466e-09 0.0007 2.469e-09 0 2.663e-09 0 2.666e-09 0.0007 2.669e-09 0 2.863e-09 0 2.866e-09 0.0007 2.869e-09 0 3.063e-09 0 3.066e-09 0.0007 3.069e-09 0 4.863e-09 0 4.866e-09 0.0007 4.869e-09 0 5.063e-09 0 5.066e-09 0.0007 5.069e-09 0 5.263e-09 0 5.266e-09 0.0007 5.269e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.663e-09 0 5.666e-09 0.0007 5.669e-09 0 5.863e-09 0 5.866e-09 0.0007 5.869e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.263e-09 0 6.266e-09 0.0007 6.269e-09 0 8.063e-09 0 8.066e-09 0.0007 8.069e-09 0 8.263e-09 0 8.266e-09 0.0007 8.269e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.663e-09 0 8.666e-09 0.0007 8.669e-09 0 8.863e-09 0 8.866e-09 0.0007 8.869e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.263e-09 0 9.266e-09 0.0007 9.269e-09 0 9.463e-09 0 9.466e-09 0.0007 9.469e-09 0 1.1263e-08 0 1.1266e-08 0.0007 1.1269e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1663e-08 0 1.1666e-08 0.0007 1.1669e-08 0 1.1863e-08 0 1.1866e-08 0.0007 1.1869e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2263e-08 0 1.2266e-08 0.0007 1.2269e-08 0 1.2463e-08 0 1.2466e-08 0.0007 1.2469e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.4463e-08 0 1.4466e-08 0.0007 1.4469e-08 0 1.4663e-08 0 1.4666e-08 0.0007 1.4669e-08 0 1.4863e-08 0 1.4866e-08 0.0007 1.4869e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5263e-08 0 1.5266e-08 0.0007 1.5269e-08 0 1.5463e-08 0 1.5466e-08 0.0007 1.5469e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5863e-08 0 1.5866e-08 0.0007 1.5869e-08 0 1.7663e-08 0 1.7666e-08 0.0007 1.7669e-08 0 1.7863e-08 0 1.7866e-08 0.0007 1.7869e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8263e-08 0 1.8266e-08 0.0007 1.8269e-08 0 1.8463e-08 0 1.8466e-08 0.0007 1.8469e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8863e-08 0 1.8866e-08 0.0007 1.8869e-08 0 1.9063e-08 0 1.9066e-08 0.0007 1.9069e-08 0 2.0863e-08 0 2.0866e-08 0.0007 2.0869e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1263e-08 0 2.1266e-08 0.0007 2.1269e-08 0 2.1463e-08 0 2.1466e-08 0.0007 2.1469e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1863e-08 0 2.1866e-08 0.0007 2.1869e-08 0 2.2063e-08 0 2.2066e-08 0.0007 2.2069e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.4063e-08 0 2.4066e-08 0.0007 2.4069e-08 0 2.4263e-08 0 2.4266e-08 0.0007 2.4269e-08 0 2.4463e-08 0 2.4466e-08 0.0007 2.4469e-08 0 2.4663e-08 0 2.4666e-08 0.0007 2.4669e-08 0 2.4863e-08 0 2.4866e-08 0.0007 2.4869e-08 0 2.5063e-08 0 2.5066e-08 0.0007 2.5069e-08 0 2.5263e-08 0 2.5266e-08 0.0007 2.5269e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 2.7263e-08 0 2.7266e-08 0.0007 2.7269e-08 0 2.7463e-08 0 2.7466e-08 0.0007 2.7469e-08 0 2.7663e-08 0 2.7666e-08 0.0007 2.7669e-08 0 2.7863e-08 0 2.7866e-08 0.0007 2.7869e-08 0 2.8063e-08 0 2.8066e-08 0.0007 2.8069e-08 0 2.8263e-08 0 2.8266e-08 0.0007 2.8269e-08 0 2.8463e-08 0 2.8466e-08 0.0007 2.8469e-08 0 2.8663e-08 0 2.8666e-08 0.0007 2.8669e-08 0 3.0463e-08 0 3.0466e-08 0.0007 3.0469e-08 0 3.0663e-08 0 3.0666e-08 0.0007 3.0669e-08 0 3.0863e-08 0 3.0866e-08 0.0007 3.0869e-08 0 3.1063e-08 0 3.1066e-08 0.0007 3.1069e-08 0 3.1263e-08 0 3.1266e-08 0.0007 3.1269e-08 0 3.1463e-08 0 3.1466e-08 0.0007 3.1469e-08 0 3.1663e-08 0 3.1666e-08 0.0007 3.1669e-08 0 3.1863e-08 0 3.1866e-08 0.0007 3.1869e-08 0 3.3663e-08 0 3.3666e-08 0.0007 3.3669e-08 0 3.3863e-08 0 3.3866e-08 0.0007 3.3869e-08 0 3.4063e-08 0 3.4066e-08 0.0007 3.4069e-08 0 3.4263e-08 0 3.4266e-08 0.0007 3.4269e-08 0 3.4463e-08 0 3.4466e-08 0.0007 3.4469e-08 0 3.4663e-08 0 3.4666e-08 0.0007 3.4669e-08 0 3.4863e-08 0 3.4866e-08 0.0007 3.4869e-08 0 3.5063e-08 0 3.5066e-08 0.0007 3.5069e-08 0 3.6863e-08 0 3.6866e-08 0.0007 3.6869e-08 0 3.7063e-08 0 3.7066e-08 0.0007 3.7069e-08 0 3.7263e-08 0 3.7266e-08 0.0007 3.7269e-08 0 3.7463e-08 0 3.7466e-08 0.0007 3.7469e-08 0 3.7663e-08 0 3.7666e-08 0.0007 3.7669e-08 0 3.7863e-08 0 3.7866e-08 0.0007 3.7869e-08 0 3.8063e-08 0 3.8066e-08 0.0007 3.8069e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 4.0063e-08 0 4.0066e-08 0.0007 4.0069e-08 0 4.0263e-08 0 4.0266e-08 0.0007 4.0269e-08 0 4.0463e-08 0 4.0466e-08 0.0007 4.0469e-08 0 4.0663e-08 0 4.0666e-08 0.0007 4.0669e-08 0 4.0863e-08 0 4.0866e-08 0.0007 4.0869e-08 0 4.1063e-08 0 4.1066e-08 0.0007 4.1069e-08 0 4.1263e-08 0 4.1266e-08 0.0007 4.1269e-08 0 4.1463e-08 0 4.1466e-08 0.0007 4.1469e-08 0 4.3263e-08 0 4.3266e-08 0.0007 4.3269e-08 0 4.3463e-08 0 4.3466e-08 0.0007 4.3469e-08 0 4.3663e-08 0 4.3666e-08 0.0007 4.3669e-08 0 4.3863e-08 0 4.3866e-08 0.0007 4.3869e-08 0 4.4063e-08 0 4.4066e-08 0.0007 4.4069e-08 0 4.4263e-08 0 4.4266e-08 0.0007 4.4269e-08 0 4.4463e-08 0 4.4466e-08 0.0007 4.4469e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.6463e-08 0 4.6466e-08 0.0007 4.6469e-08 0 4.6663e-08 0 4.6666e-08 0.0007 4.6669e-08 0 4.6863e-08 0 4.6866e-08 0.0007 4.6869e-08 0 4.7063e-08 0 4.7066e-08 0.0007 4.7069e-08 0 4.7263e-08 0 4.7266e-08 0.0007 4.7269e-08 0 4.7463e-08 0 4.7466e-08 0.0007 4.7469e-08 0 4.7663e-08 0 4.7666e-08 0.0007 4.7669e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.9663e-08 0 4.9666e-08 0.0007 4.9669e-08 0 4.9863e-08 0 4.9866e-08 0.0007 4.9869e-08 0 5.0063e-08 0 5.0066e-08 0.0007 5.0069e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0463e-08 0 5.0466e-08 0.0007 5.0469e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA4|E 0 A4_TX  PWL(0 0 3.263e-09 0 3.266e-09 0.0007 3.269e-09 0 3.463e-09 0 3.466e-09 0.0007 3.469e-09 0 3.663e-09 0 3.666e-09 0.0007 3.669e-09 0 3.863e-09 0 3.866e-09 0.0007 3.869e-09 0 4.063e-09 0 4.066e-09 0.0007 4.069e-09 0 4.263e-09 0 4.266e-09 0.0007 4.269e-09 0 4.463e-09 0 4.466e-09 0.0007 4.469e-09 0 4.663e-09 0 4.666e-09 0.0007 4.669e-09 0 4.863e-09 0 4.866e-09 0.0007 4.869e-09 0 5.063e-09 0 5.066e-09 0.0007 5.069e-09 0 5.263e-09 0 5.266e-09 0.0007 5.269e-09 0 5.463e-09 0 5.466e-09 0.0007 5.469e-09 0 5.663e-09 0 5.666e-09 0.0007 5.669e-09 0 5.863e-09 0 5.866e-09 0.0007 5.869e-09 0 6.063e-09 0 6.066e-09 0.0007 6.069e-09 0 6.263e-09 0 6.266e-09 0.0007 6.269e-09 0 9.663e-09 0 9.666e-09 0.0007 9.669e-09 0 9.863e-09 0 9.866e-09 0.0007 9.869e-09 0 1.0063e-08 0 1.0066e-08 0.0007 1.0069e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0463e-08 0 1.0466e-08 0.0007 1.0469e-08 0 1.0663e-08 0 1.0666e-08 0.0007 1.0669e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.1063e-08 0 1.1066e-08 0.0007 1.1069e-08 0 1.1263e-08 0 1.1266e-08 0.0007 1.1269e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1663e-08 0 1.1666e-08 0.0007 1.1669e-08 0 1.1863e-08 0 1.1866e-08 0.0007 1.1869e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2263e-08 0 1.2266e-08 0.0007 1.2269e-08 0 1.2463e-08 0 1.2466e-08 0.0007 1.2469e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.6063e-08 0 1.6066e-08 0.0007 1.6069e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6463e-08 0 1.6466e-08 0.0007 1.6469e-08 0 1.6663e-08 0 1.6666e-08 0.0007 1.6669e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.7063e-08 0 1.7066e-08 0.0007 1.7069e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.7269e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7663e-08 0 1.7666e-08 0.0007 1.7669e-08 0 1.7863e-08 0 1.7866e-08 0.0007 1.7869e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8263e-08 0 1.8266e-08 0.0007 1.8269e-08 0 1.8463e-08 0 1.8466e-08 0.0007 1.8469e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8863e-08 0 1.8866e-08 0.0007 1.8869e-08 0 1.9063e-08 0 1.9066e-08 0.0007 1.9069e-08 0 2.2463e-08 0 2.2466e-08 0.0007 2.2469e-08 0 2.2663e-08 0 2.2666e-08 0.0007 2.2669e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.3063e-08 0 2.3066e-08 0.0007 2.3069e-08 0 2.3263e-08 0 2.3266e-08 0.0007 2.3269e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3663e-08 0 2.3666e-08 0.0007 2.3669e-08 0 2.3863e-08 0 2.3866e-08 0.0007 2.3869e-08 0 2.4063e-08 0 2.4066e-08 0.0007 2.4069e-08 0 2.4263e-08 0 2.4266e-08 0.0007 2.4269e-08 0 2.4463e-08 0 2.4466e-08 0.0007 2.4469e-08 0 2.4663e-08 0 2.4666e-08 0.0007 2.4669e-08 0 2.4863e-08 0 2.4866e-08 0.0007 2.4869e-08 0 2.5063e-08 0 2.5066e-08 0.0007 2.5069e-08 0 2.5263e-08 0 2.5266e-08 0.0007 2.5269e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 2.8863e-08 0 2.8866e-08 0.0007 2.8869e-08 0 2.9063e-08 0 2.9066e-08 0.0007 2.9069e-08 0 2.9263e-08 0 2.9266e-08 0.0007 2.9269e-08 0 2.9463e-08 0 2.9466e-08 0.0007 2.9469e-08 0 2.9663e-08 0 2.9666e-08 0.0007 2.9669e-08 0 2.9863e-08 0 2.9866e-08 0.0007 2.9869e-08 0 3.0063e-08 0 3.0066e-08 0.0007 3.0069e-08 0 3.0263e-08 0 3.0266e-08 0.0007 3.0269e-08 0 3.0463e-08 0 3.0466e-08 0.0007 3.0469e-08 0 3.0663e-08 0 3.0666e-08 0.0007 3.0669e-08 0 3.0863e-08 0 3.0866e-08 0.0007 3.0869e-08 0 3.1063e-08 0 3.1066e-08 0.0007 3.1069e-08 0 3.1263e-08 0 3.1266e-08 0.0007 3.1269e-08 0 3.1463e-08 0 3.1466e-08 0.0007 3.1469e-08 0 3.1663e-08 0 3.1666e-08 0.0007 3.1669e-08 0 3.1863e-08 0 3.1866e-08 0.0007 3.1869e-08 0 3.5263e-08 0 3.5266e-08 0.0007 3.5269e-08 0 3.5463e-08 0 3.5466e-08 0.0007 3.5469e-08 0 3.5663e-08 0 3.5666e-08 0.0007 3.5669e-08 0 3.5863e-08 0 3.5866e-08 0.0007 3.5869e-08 0 3.6063e-08 0 3.6066e-08 0.0007 3.6069e-08 0 3.6263e-08 0 3.6266e-08 0.0007 3.6269e-08 0 3.6463e-08 0 3.6466e-08 0.0007 3.6469e-08 0 3.6663e-08 0 3.6666e-08 0.0007 3.6669e-08 0 3.6863e-08 0 3.6866e-08 0.0007 3.6869e-08 0 3.7063e-08 0 3.7066e-08 0.0007 3.7069e-08 0 3.7263e-08 0 3.7266e-08 0.0007 3.7269e-08 0 3.7463e-08 0 3.7466e-08 0.0007 3.7469e-08 0 3.7663e-08 0 3.7666e-08 0.0007 3.7669e-08 0 3.7863e-08 0 3.7866e-08 0.0007 3.7869e-08 0 3.8063e-08 0 3.8066e-08 0.0007 3.8069e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 4.1663e-08 0 4.1666e-08 0.0007 4.1669e-08 0 4.1863e-08 0 4.1866e-08 0.0007 4.1869e-08 0 4.2063e-08 0 4.2066e-08 0.0007 4.2069e-08 0 4.2263e-08 0 4.2266e-08 0.0007 4.2269e-08 0 4.2463e-08 0 4.2466e-08 0.0007 4.2469e-08 0 4.2663e-08 0 4.2666e-08 0.0007 4.2669e-08 0 4.2863e-08 0 4.2866e-08 0.0007 4.2869e-08 0 4.3063e-08 0 4.3066e-08 0.0007 4.3069e-08 0 4.3263e-08 0 4.3266e-08 0.0007 4.3269e-08 0 4.3463e-08 0 4.3466e-08 0.0007 4.3469e-08 0 4.3663e-08 0 4.3666e-08 0.0007 4.3669e-08 0 4.3863e-08 0 4.3866e-08 0.0007 4.3869e-08 0 4.4063e-08 0 4.4066e-08 0.0007 4.4069e-08 0 4.4263e-08 0 4.4266e-08 0.0007 4.4269e-08 0 4.4463e-08 0 4.4466e-08 0.0007 4.4469e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.8063e-08 0 4.8066e-08 0.0007 4.8069e-08 0 4.8263e-08 0 4.8266e-08 0.0007 4.8269e-08 0 4.8463e-08 0 4.8466e-08 0.0007 4.8469e-08 0 4.8663e-08 0 4.8666e-08 0.0007 4.8669e-08 0 4.8863e-08 0 4.8866e-08 0.0007 4.8869e-08 0 4.9063e-08 0 4.9066e-08 0.0007 4.9069e-08 0 4.9263e-08 0 4.9266e-08 0.0007 4.9269e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 4.9663e-08 0 4.9666e-08 0.0007 4.9669e-08 0 4.9863e-08 0 4.9866e-08 0.0007 4.9869e-08 0 5.0063e-08 0 5.0066e-08 0.0007 5.0069e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0463e-08 0 5.0466e-08 0.0007 5.0469e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA5|F 0 A5_TX  PWL(0 0 6.463e-09 0 6.466e-09 0.0007 6.469e-09 0 6.663e-09 0 6.666e-09 0.0007 6.669e-09 0 6.863e-09 0 6.866e-09 0.0007 6.869e-09 0 7.063e-09 0 7.066e-09 0.0007 7.069e-09 0 7.263e-09 0 7.266e-09 0.0007 7.269e-09 0 7.463e-09 0 7.466e-09 0.0007 7.469e-09 0 7.663e-09 0 7.666e-09 0.0007 7.669e-09 0 7.863e-09 0 7.866e-09 0.0007 7.869e-09 0 8.063e-09 0 8.066e-09 0.0007 8.069e-09 0 8.263e-09 0 8.266e-09 0.0007 8.269e-09 0 8.463e-09 0 8.466e-09 0.0007 8.469e-09 0 8.663e-09 0 8.666e-09 0.0007 8.669e-09 0 8.863e-09 0 8.866e-09 0.0007 8.869e-09 0 9.063e-09 0 9.066e-09 0.0007 9.069e-09 0 9.263e-09 0 9.266e-09 0.0007 9.269e-09 0 9.463e-09 0 9.466e-09 0.0007 9.469e-09 0 9.663e-09 0 9.666e-09 0.0007 9.669e-09 0 9.863e-09 0 9.866e-09 0.0007 9.869e-09 0 1.0063e-08 0 1.0066e-08 0.0007 1.0069e-08 0 1.0263e-08 0 1.0266e-08 0.0007 1.0269e-08 0 1.0463e-08 0 1.0466e-08 0.0007 1.0469e-08 0 1.0663e-08 0 1.0666e-08 0.0007 1.0669e-08 0 1.0863e-08 0 1.0866e-08 0.0007 1.0869e-08 0 1.1063e-08 0 1.1066e-08 0.0007 1.1069e-08 0 1.1263e-08 0 1.1266e-08 0.0007 1.1269e-08 0 1.1463e-08 0 1.1466e-08 0.0007 1.1469e-08 0 1.1663e-08 0 1.1666e-08 0.0007 1.1669e-08 0 1.1863e-08 0 1.1866e-08 0.0007 1.1869e-08 0 1.2063e-08 0 1.2066e-08 0.0007 1.2069e-08 0 1.2263e-08 0 1.2266e-08 0.0007 1.2269e-08 0 1.2463e-08 0 1.2466e-08 0.0007 1.2469e-08 0 1.2663e-08 0 1.2666e-08 0.0007 1.2669e-08 0 1.9263e-08 0 1.9266e-08 0.0007 1.9269e-08 0 1.9463e-08 0 1.9466e-08 0.0007 1.9469e-08 0 1.9663e-08 0 1.9666e-08 0.0007 1.9669e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 2.0063e-08 0 2.0066e-08 0.0007 2.0069e-08 0 2.0263e-08 0 2.0266e-08 0.0007 2.0269e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0663e-08 0 2.0666e-08 0.0007 2.0669e-08 0 2.0863e-08 0 2.0866e-08 0.0007 2.0869e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1263e-08 0 2.1266e-08 0.0007 2.1269e-08 0 2.1463e-08 0 2.1466e-08 0.0007 2.1469e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1863e-08 0 2.1866e-08 0.0007 2.1869e-08 0 2.2063e-08 0 2.2066e-08 0.0007 2.2069e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2463e-08 0 2.2466e-08 0.0007 2.2469e-08 0 2.2663e-08 0 2.2666e-08 0.0007 2.2669e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.3063e-08 0 2.3066e-08 0.0007 2.3069e-08 0 2.3263e-08 0 2.3266e-08 0.0007 2.3269e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3663e-08 0 2.3666e-08 0.0007 2.3669e-08 0 2.3863e-08 0 2.3866e-08 0.0007 2.3869e-08 0 2.4063e-08 0 2.4066e-08 0.0007 2.4069e-08 0 2.4263e-08 0 2.4266e-08 0.0007 2.4269e-08 0 2.4463e-08 0 2.4466e-08 0.0007 2.4469e-08 0 2.4663e-08 0 2.4666e-08 0.0007 2.4669e-08 0 2.4863e-08 0 2.4866e-08 0.0007 2.4869e-08 0 2.5063e-08 0 2.5066e-08 0.0007 2.5069e-08 0 2.5263e-08 0 2.5266e-08 0.0007 2.5269e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 3.2063e-08 0 3.2066e-08 0.0007 3.2069e-08 0 3.2263e-08 0 3.2266e-08 0.0007 3.2269e-08 0 3.2463e-08 0 3.2466e-08 0.0007 3.2469e-08 0 3.2663e-08 0 3.2666e-08 0.0007 3.2669e-08 0 3.2863e-08 0 3.2866e-08 0.0007 3.2869e-08 0 3.3063e-08 0 3.3066e-08 0.0007 3.3069e-08 0 3.3263e-08 0 3.3266e-08 0.0007 3.3269e-08 0 3.3463e-08 0 3.3466e-08 0.0007 3.3469e-08 0 3.3663e-08 0 3.3666e-08 0.0007 3.3669e-08 0 3.3863e-08 0 3.3866e-08 0.0007 3.3869e-08 0 3.4063e-08 0 3.4066e-08 0.0007 3.4069e-08 0 3.4263e-08 0 3.4266e-08 0.0007 3.4269e-08 0 3.4463e-08 0 3.4466e-08 0.0007 3.4469e-08 0 3.4663e-08 0 3.4666e-08 0.0007 3.4669e-08 0 3.4863e-08 0 3.4866e-08 0.0007 3.4869e-08 0 3.5063e-08 0 3.5066e-08 0.0007 3.5069e-08 0 3.5263e-08 0 3.5266e-08 0.0007 3.5269e-08 0 3.5463e-08 0 3.5466e-08 0.0007 3.5469e-08 0 3.5663e-08 0 3.5666e-08 0.0007 3.5669e-08 0 3.5863e-08 0 3.5866e-08 0.0007 3.5869e-08 0 3.6063e-08 0 3.6066e-08 0.0007 3.6069e-08 0 3.6263e-08 0 3.6266e-08 0.0007 3.6269e-08 0 3.6463e-08 0 3.6466e-08 0.0007 3.6469e-08 0 3.6663e-08 0 3.6666e-08 0.0007 3.6669e-08 0 3.6863e-08 0 3.6866e-08 0.0007 3.6869e-08 0 3.7063e-08 0 3.7066e-08 0.0007 3.7069e-08 0 3.7263e-08 0 3.7266e-08 0.0007 3.7269e-08 0 3.7463e-08 0 3.7466e-08 0.0007 3.7469e-08 0 3.7663e-08 0 3.7666e-08 0.0007 3.7669e-08 0 3.7863e-08 0 3.7866e-08 0.0007 3.7869e-08 0 3.8063e-08 0 3.8066e-08 0.0007 3.8069e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 4.4863e-08 0 4.4866e-08 0.0007 4.4869e-08 0 4.5063e-08 0 4.5066e-08 0.0007 4.5069e-08 0 4.5263e-08 0 4.5266e-08 0.0007 4.5269e-08 0 4.5463e-08 0 4.5466e-08 0.0007 4.5469e-08 0 4.5663e-08 0 4.5666e-08 0.0007 4.5669e-08 0 4.5863e-08 0 4.5866e-08 0.0007 4.5869e-08 0 4.6063e-08 0 4.6066e-08 0.0007 4.6069e-08 0 4.6263e-08 0 4.6266e-08 0.0007 4.6269e-08 0 4.6463e-08 0 4.6466e-08 0.0007 4.6469e-08 0 4.6663e-08 0 4.6666e-08 0.0007 4.6669e-08 0 4.6863e-08 0 4.6866e-08 0.0007 4.6869e-08 0 4.7063e-08 0 4.7066e-08 0.0007 4.7069e-08 0 4.7263e-08 0 4.7266e-08 0.0007 4.7269e-08 0 4.7463e-08 0 4.7466e-08 0.0007 4.7469e-08 0 4.7663e-08 0 4.7666e-08 0.0007 4.7669e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.8063e-08 0 4.8066e-08 0.0007 4.8069e-08 0 4.8263e-08 0 4.8266e-08 0.0007 4.8269e-08 0 4.8463e-08 0 4.8466e-08 0.0007 4.8469e-08 0 4.8663e-08 0 4.8666e-08 0.0007 4.8669e-08 0 4.8863e-08 0 4.8866e-08 0.0007 4.8869e-08 0 4.9063e-08 0 4.9066e-08 0.0007 4.9069e-08 0 4.9263e-08 0 4.9266e-08 0.0007 4.9269e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 4.9663e-08 0 4.9666e-08 0.0007 4.9669e-08 0 4.9863e-08 0 4.9866e-08 0.0007 4.9869e-08 0 5.0063e-08 0 5.0066e-08 0.0007 5.0069e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0463e-08 0 5.0466e-08 0.0007 5.0469e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA6|G 0 A6_TX  PWL(0 0 1.2863e-08 0 1.2866e-08 0.0007 1.2869e-08 0 1.3063e-08 0 1.3066e-08 0.0007 1.3069e-08 0 1.3263e-08 0 1.3266e-08 0.0007 1.3269e-08 0 1.3463e-08 0 1.3466e-08 0.0007 1.3469e-08 0 1.3663e-08 0 1.3666e-08 0.0007 1.3669e-08 0 1.3863e-08 0 1.3866e-08 0.0007 1.3869e-08 0 1.4063e-08 0 1.4066e-08 0.0007 1.4069e-08 0 1.4263e-08 0 1.4266e-08 0.0007 1.4269e-08 0 1.4463e-08 0 1.4466e-08 0.0007 1.4469e-08 0 1.4663e-08 0 1.4666e-08 0.0007 1.4669e-08 0 1.4863e-08 0 1.4866e-08 0.0007 1.4869e-08 0 1.5063e-08 0 1.5066e-08 0.0007 1.5069e-08 0 1.5263e-08 0 1.5266e-08 0.0007 1.5269e-08 0 1.5463e-08 0 1.5466e-08 0.0007 1.5469e-08 0 1.5663e-08 0 1.5666e-08 0.0007 1.5669e-08 0 1.5863e-08 0 1.5866e-08 0.0007 1.5869e-08 0 1.6063e-08 0 1.6066e-08 0.0007 1.6069e-08 0 1.6263e-08 0 1.6266e-08 0.0007 1.6269e-08 0 1.6463e-08 0 1.6466e-08 0.0007 1.6469e-08 0 1.6663e-08 0 1.6666e-08 0.0007 1.6669e-08 0 1.6863e-08 0 1.6866e-08 0.0007 1.6869e-08 0 1.7063e-08 0 1.7066e-08 0.0007 1.7069e-08 0 1.7263e-08 0 1.7266e-08 0.0007 1.7269e-08 0 1.7463e-08 0 1.7466e-08 0.0007 1.7469e-08 0 1.7663e-08 0 1.7666e-08 0.0007 1.7669e-08 0 1.7863e-08 0 1.7866e-08 0.0007 1.7869e-08 0 1.8063e-08 0 1.8066e-08 0.0007 1.8069e-08 0 1.8263e-08 0 1.8266e-08 0.0007 1.8269e-08 0 1.8463e-08 0 1.8466e-08 0.0007 1.8469e-08 0 1.8663e-08 0 1.8666e-08 0.0007 1.8669e-08 0 1.8863e-08 0 1.8866e-08 0.0007 1.8869e-08 0 1.9063e-08 0 1.9066e-08 0.0007 1.9069e-08 0 1.9263e-08 0 1.9266e-08 0.0007 1.9269e-08 0 1.9463e-08 0 1.9466e-08 0.0007 1.9469e-08 0 1.9663e-08 0 1.9666e-08 0.0007 1.9669e-08 0 1.9863e-08 0 1.9866e-08 0.0007 1.9869e-08 0 2.0063e-08 0 2.0066e-08 0.0007 2.0069e-08 0 2.0263e-08 0 2.0266e-08 0.0007 2.0269e-08 0 2.0463e-08 0 2.0466e-08 0.0007 2.0469e-08 0 2.0663e-08 0 2.0666e-08 0.0007 2.0669e-08 0 2.0863e-08 0 2.0866e-08 0.0007 2.0869e-08 0 2.1063e-08 0 2.1066e-08 0.0007 2.1069e-08 0 2.1263e-08 0 2.1266e-08 0.0007 2.1269e-08 0 2.1463e-08 0 2.1466e-08 0.0007 2.1469e-08 0 2.1663e-08 0 2.1666e-08 0.0007 2.1669e-08 0 2.1863e-08 0 2.1866e-08 0.0007 2.1869e-08 0 2.2063e-08 0 2.2066e-08 0.0007 2.2069e-08 0 2.2263e-08 0 2.2266e-08 0.0007 2.2269e-08 0 2.2463e-08 0 2.2466e-08 0.0007 2.2469e-08 0 2.2663e-08 0 2.2666e-08 0.0007 2.2669e-08 0 2.2863e-08 0 2.2866e-08 0.0007 2.2869e-08 0 2.3063e-08 0 2.3066e-08 0.0007 2.3069e-08 0 2.3263e-08 0 2.3266e-08 0.0007 2.3269e-08 0 2.3463e-08 0 2.3466e-08 0.0007 2.3469e-08 0 2.3663e-08 0 2.3666e-08 0.0007 2.3669e-08 0 2.3863e-08 0 2.3866e-08 0.0007 2.3869e-08 0 2.4063e-08 0 2.4066e-08 0.0007 2.4069e-08 0 2.4263e-08 0 2.4266e-08 0.0007 2.4269e-08 0 2.4463e-08 0 2.4466e-08 0.0007 2.4469e-08 0 2.4663e-08 0 2.4666e-08 0.0007 2.4669e-08 0 2.4863e-08 0 2.4866e-08 0.0007 2.4869e-08 0 2.5063e-08 0 2.5066e-08 0.0007 2.5069e-08 0 2.5263e-08 0 2.5266e-08 0.0007 2.5269e-08 0 2.5463e-08 0 2.5466e-08 0.0007 2.5469e-08 0 3.8463e-08 0 3.8466e-08 0.0007 3.8469e-08 0 3.8663e-08 0 3.8666e-08 0.0007 3.8669e-08 0 3.8863e-08 0 3.8866e-08 0.0007 3.8869e-08 0 3.9063e-08 0 3.9066e-08 0.0007 3.9069e-08 0 3.9263e-08 0 3.9266e-08 0.0007 3.9269e-08 0 3.9463e-08 0 3.9466e-08 0.0007 3.9469e-08 0 3.9663e-08 0 3.9666e-08 0.0007 3.9669e-08 0 3.9863e-08 0 3.9866e-08 0.0007 3.9869e-08 0 4.0063e-08 0 4.0066e-08 0.0007 4.0069e-08 0 4.0263e-08 0 4.0266e-08 0.0007 4.0269e-08 0 4.0463e-08 0 4.0466e-08 0.0007 4.0469e-08 0 4.0663e-08 0 4.0666e-08 0.0007 4.0669e-08 0 4.0863e-08 0 4.0866e-08 0.0007 4.0869e-08 0 4.1063e-08 0 4.1066e-08 0.0007 4.1069e-08 0 4.1263e-08 0 4.1266e-08 0.0007 4.1269e-08 0 4.1463e-08 0 4.1466e-08 0.0007 4.1469e-08 0 4.1663e-08 0 4.1666e-08 0.0007 4.1669e-08 0 4.1863e-08 0 4.1866e-08 0.0007 4.1869e-08 0 4.2063e-08 0 4.2066e-08 0.0007 4.2069e-08 0 4.2263e-08 0 4.2266e-08 0.0007 4.2269e-08 0 4.2463e-08 0 4.2466e-08 0.0007 4.2469e-08 0 4.2663e-08 0 4.2666e-08 0.0007 4.2669e-08 0 4.2863e-08 0 4.2866e-08 0.0007 4.2869e-08 0 4.3063e-08 0 4.3066e-08 0.0007 4.3069e-08 0 4.3263e-08 0 4.3266e-08 0.0007 4.3269e-08 0 4.3463e-08 0 4.3466e-08 0.0007 4.3469e-08 0 4.3663e-08 0 4.3666e-08 0.0007 4.3669e-08 0 4.3863e-08 0 4.3866e-08 0.0007 4.3869e-08 0 4.4063e-08 0 4.4066e-08 0.0007 4.4069e-08 0 4.4263e-08 0 4.4266e-08 0.0007 4.4269e-08 0 4.4463e-08 0 4.4466e-08 0.0007 4.4469e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.4863e-08 0 4.4866e-08 0.0007 4.4869e-08 0 4.5063e-08 0 4.5066e-08 0.0007 4.5069e-08 0 4.5263e-08 0 4.5266e-08 0.0007 4.5269e-08 0 4.5463e-08 0 4.5466e-08 0.0007 4.5469e-08 0 4.5663e-08 0 4.5666e-08 0.0007 4.5669e-08 0 4.5863e-08 0 4.5866e-08 0.0007 4.5869e-08 0 4.6063e-08 0 4.6066e-08 0.0007 4.6069e-08 0 4.6263e-08 0 4.6266e-08 0.0007 4.6269e-08 0 4.6463e-08 0 4.6466e-08 0.0007 4.6469e-08 0 4.6663e-08 0 4.6666e-08 0.0007 4.6669e-08 0 4.6863e-08 0 4.6866e-08 0.0007 4.6869e-08 0 4.7063e-08 0 4.7066e-08 0.0007 4.7069e-08 0 4.7263e-08 0 4.7266e-08 0.0007 4.7269e-08 0 4.7463e-08 0 4.7466e-08 0.0007 4.7469e-08 0 4.7663e-08 0 4.7666e-08 0.0007 4.7669e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.8063e-08 0 4.8066e-08 0.0007 4.8069e-08 0 4.8263e-08 0 4.8266e-08 0.0007 4.8269e-08 0 4.8463e-08 0 4.8466e-08 0.0007 4.8469e-08 0 4.8663e-08 0 4.8666e-08 0.0007 4.8669e-08 0 4.8863e-08 0 4.8866e-08 0.0007 4.8869e-08 0 4.9063e-08 0 4.9066e-08 0.0007 4.9069e-08 0 4.9263e-08 0 4.9266e-08 0.0007 4.9269e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 4.9663e-08 0 4.9666e-08 0.0007 4.9669e-08 0 4.9863e-08 0 4.9866e-08 0.0007 4.9869e-08 0 5.0063e-08 0 5.0066e-08 0.0007 5.0069e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0463e-08 0 5.0466e-08 0.0007 5.0469e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IA7|H 0 A7_TX  PWL(0 0 2.5663e-08 0 2.5666e-08 0.0007 2.5669e-08 0 2.5863e-08 0 2.5866e-08 0.0007 2.5869e-08 0 2.6063e-08 0 2.6066e-08 0.0007 2.6069e-08 0 2.6263e-08 0 2.6266e-08 0.0007 2.6269e-08 0 2.6463e-08 0 2.6466e-08 0.0007 2.6469e-08 0 2.6663e-08 0 2.6666e-08 0.0007 2.6669e-08 0 2.6863e-08 0 2.6866e-08 0.0007 2.6869e-08 0 2.7063e-08 0 2.7066e-08 0.0007 2.7069e-08 0 2.7263e-08 0 2.7266e-08 0.0007 2.7269e-08 0 2.7463e-08 0 2.7466e-08 0.0007 2.7469e-08 0 2.7663e-08 0 2.7666e-08 0.0007 2.7669e-08 0 2.7863e-08 0 2.7866e-08 0.0007 2.7869e-08 0 2.8063e-08 0 2.8066e-08 0.0007 2.8069e-08 0 2.8263e-08 0 2.8266e-08 0.0007 2.8269e-08 0 2.8463e-08 0 2.8466e-08 0.0007 2.8469e-08 0 2.8663e-08 0 2.8666e-08 0.0007 2.8669e-08 0 2.8863e-08 0 2.8866e-08 0.0007 2.8869e-08 0 2.9063e-08 0 2.9066e-08 0.0007 2.9069e-08 0 2.9263e-08 0 2.9266e-08 0.0007 2.9269e-08 0 2.9463e-08 0 2.9466e-08 0.0007 2.9469e-08 0 2.9663e-08 0 2.9666e-08 0.0007 2.9669e-08 0 2.9863e-08 0 2.9866e-08 0.0007 2.9869e-08 0 3.0063e-08 0 3.0066e-08 0.0007 3.0069e-08 0 3.0263e-08 0 3.0266e-08 0.0007 3.0269e-08 0 3.0463e-08 0 3.0466e-08 0.0007 3.0469e-08 0 3.0663e-08 0 3.0666e-08 0.0007 3.0669e-08 0 3.0863e-08 0 3.0866e-08 0.0007 3.0869e-08 0 3.1063e-08 0 3.1066e-08 0.0007 3.1069e-08 0 3.1263e-08 0 3.1266e-08 0.0007 3.1269e-08 0 3.1463e-08 0 3.1466e-08 0.0007 3.1469e-08 0 3.1663e-08 0 3.1666e-08 0.0007 3.1669e-08 0 3.1863e-08 0 3.1866e-08 0.0007 3.1869e-08 0 3.2063e-08 0 3.2066e-08 0.0007 3.2069e-08 0 3.2263e-08 0 3.2266e-08 0.0007 3.2269e-08 0 3.2463e-08 0 3.2466e-08 0.0007 3.2469e-08 0 3.2663e-08 0 3.2666e-08 0.0007 3.2669e-08 0 3.2863e-08 0 3.2866e-08 0.0007 3.2869e-08 0 3.3063e-08 0 3.3066e-08 0.0007 3.3069e-08 0 3.3263e-08 0 3.3266e-08 0.0007 3.3269e-08 0 3.3463e-08 0 3.3466e-08 0.0007 3.3469e-08 0 3.3663e-08 0 3.3666e-08 0.0007 3.3669e-08 0 3.3863e-08 0 3.3866e-08 0.0007 3.3869e-08 0 3.4063e-08 0 3.4066e-08 0.0007 3.4069e-08 0 3.4263e-08 0 3.4266e-08 0.0007 3.4269e-08 0 3.4463e-08 0 3.4466e-08 0.0007 3.4469e-08 0 3.4663e-08 0 3.4666e-08 0.0007 3.4669e-08 0 3.4863e-08 0 3.4866e-08 0.0007 3.4869e-08 0 3.5063e-08 0 3.5066e-08 0.0007 3.5069e-08 0 3.5263e-08 0 3.5266e-08 0.0007 3.5269e-08 0 3.5463e-08 0 3.5466e-08 0.0007 3.5469e-08 0 3.5663e-08 0 3.5666e-08 0.0007 3.5669e-08 0 3.5863e-08 0 3.5866e-08 0.0007 3.5869e-08 0 3.6063e-08 0 3.6066e-08 0.0007 3.6069e-08 0 3.6263e-08 0 3.6266e-08 0.0007 3.6269e-08 0 3.6463e-08 0 3.6466e-08 0.0007 3.6469e-08 0 3.6663e-08 0 3.6666e-08 0.0007 3.6669e-08 0 3.6863e-08 0 3.6866e-08 0.0007 3.6869e-08 0 3.7063e-08 0 3.7066e-08 0.0007 3.7069e-08 0 3.7263e-08 0 3.7266e-08 0.0007 3.7269e-08 0 3.7463e-08 0 3.7466e-08 0.0007 3.7469e-08 0 3.7663e-08 0 3.7666e-08 0.0007 3.7669e-08 0 3.7863e-08 0 3.7866e-08 0.0007 3.7869e-08 0 3.8063e-08 0 3.8066e-08 0.0007 3.8069e-08 0 3.8263e-08 0 3.8266e-08 0.0007 3.8269e-08 0 3.8463e-08 0 3.8466e-08 0.0007 3.8469e-08 0 3.8663e-08 0 3.8666e-08 0.0007 3.8669e-08 0 3.8863e-08 0 3.8866e-08 0.0007 3.8869e-08 0 3.9063e-08 0 3.9066e-08 0.0007 3.9069e-08 0 3.9263e-08 0 3.9266e-08 0.0007 3.9269e-08 0 3.9463e-08 0 3.9466e-08 0.0007 3.9469e-08 0 3.9663e-08 0 3.9666e-08 0.0007 3.9669e-08 0 3.9863e-08 0 3.9866e-08 0.0007 3.9869e-08 0 4.0063e-08 0 4.0066e-08 0.0007 4.0069e-08 0 4.0263e-08 0 4.0266e-08 0.0007 4.0269e-08 0 4.0463e-08 0 4.0466e-08 0.0007 4.0469e-08 0 4.0663e-08 0 4.0666e-08 0.0007 4.0669e-08 0 4.0863e-08 0 4.0866e-08 0.0007 4.0869e-08 0 4.1063e-08 0 4.1066e-08 0.0007 4.1069e-08 0 4.1263e-08 0 4.1266e-08 0.0007 4.1269e-08 0 4.1463e-08 0 4.1466e-08 0.0007 4.1469e-08 0 4.1663e-08 0 4.1666e-08 0.0007 4.1669e-08 0 4.1863e-08 0 4.1866e-08 0.0007 4.1869e-08 0 4.2063e-08 0 4.2066e-08 0.0007 4.2069e-08 0 4.2263e-08 0 4.2266e-08 0.0007 4.2269e-08 0 4.2463e-08 0 4.2466e-08 0.0007 4.2469e-08 0 4.2663e-08 0 4.2666e-08 0.0007 4.2669e-08 0 4.2863e-08 0 4.2866e-08 0.0007 4.2869e-08 0 4.3063e-08 0 4.3066e-08 0.0007 4.3069e-08 0 4.3263e-08 0 4.3266e-08 0.0007 4.3269e-08 0 4.3463e-08 0 4.3466e-08 0.0007 4.3469e-08 0 4.3663e-08 0 4.3666e-08 0.0007 4.3669e-08 0 4.3863e-08 0 4.3866e-08 0.0007 4.3869e-08 0 4.4063e-08 0 4.4066e-08 0.0007 4.4069e-08 0 4.4263e-08 0 4.4266e-08 0.0007 4.4269e-08 0 4.4463e-08 0 4.4466e-08 0.0007 4.4469e-08 0 4.4663e-08 0 4.4666e-08 0.0007 4.4669e-08 0 4.4863e-08 0 4.4866e-08 0.0007 4.4869e-08 0 4.5063e-08 0 4.5066e-08 0.0007 4.5069e-08 0 4.5263e-08 0 4.5266e-08 0.0007 4.5269e-08 0 4.5463e-08 0 4.5466e-08 0.0007 4.5469e-08 0 4.5663e-08 0 4.5666e-08 0.0007 4.5669e-08 0 4.5863e-08 0 4.5866e-08 0.0007 4.5869e-08 0 4.6063e-08 0 4.6066e-08 0.0007 4.6069e-08 0 4.6263e-08 0 4.6266e-08 0.0007 4.6269e-08 0 4.6463e-08 0 4.6466e-08 0.0007 4.6469e-08 0 4.6663e-08 0 4.6666e-08 0.0007 4.6669e-08 0 4.6863e-08 0 4.6866e-08 0.0007 4.6869e-08 0 4.7063e-08 0 4.7066e-08 0.0007 4.7069e-08 0 4.7263e-08 0 4.7266e-08 0.0007 4.7269e-08 0 4.7463e-08 0 4.7466e-08 0.0007 4.7469e-08 0 4.7663e-08 0 4.7666e-08 0.0007 4.7669e-08 0 4.7863e-08 0 4.7866e-08 0.0007 4.7869e-08 0 4.8063e-08 0 4.8066e-08 0.0007 4.8069e-08 0 4.8263e-08 0 4.8266e-08 0.0007 4.8269e-08 0 4.8463e-08 0 4.8466e-08 0.0007 4.8469e-08 0 4.8663e-08 0 4.8666e-08 0.0007 4.8669e-08 0 4.8863e-08 0 4.8866e-08 0.0007 4.8869e-08 0 4.9063e-08 0 4.9066e-08 0.0007 4.9069e-08 0 4.9263e-08 0 4.9266e-08 0.0007 4.9269e-08 0 4.9463e-08 0 4.9466e-08 0.0007 4.9469e-08 0 4.9663e-08 0 4.9666e-08 0.0007 4.9669e-08 0 4.9863e-08 0 4.9866e-08 0.0007 4.9869e-08 0 5.0063e-08 0 5.0066e-08 0.0007 5.0069e-08 0 5.0263e-08 0 5.0266e-08 0.0007 5.0269e-08 0 5.0463e-08 0 5.0466e-08 0.0007 5.0469e-08 0 5.0663e-08 0 5.0666e-08 0.0007 5.0669e-08 0 5.0863e-08 0 5.0866e-08 0.0007 5.0869e-08 0 5.1063e-08 0 5.1066e-08 0.0007 5.1069e-08 0)
IB0|T 0 B0_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB1|T 0 B1_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB2|T 0 B2_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB3|T 0 B3_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB4|T 0 B4_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB5|T 0 B5_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB6|T 0 B6_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IB7|T 0 B7_TX  PWL(0 0 4.7e-11 0 5e-11 0.0007 5.3e-11 0 2.47e-10 0 2.5e-10 0.0007 2.53e-10 0 4.47e-10 0 4.5e-10 0.0007 4.53e-10 0 6.47e-10 0 6.5e-10 0.0007 6.53e-10 0 8.47e-10 0 8.5e-10 0.0007 8.53e-10 0 1.047e-09 0 1.05e-09 0.0007 1.053e-09 0 1.247e-09 0 1.25e-09 0.0007 1.253e-09 0 1.447e-09 0 1.45e-09 0.0007 1.453e-09 0 1.647e-09 0 1.65e-09 0.0007 1.653e-09 0 1.847e-09 0 1.85e-09 0.0007 1.853e-09 0 2.047e-09 0 2.05e-09 0.0007 2.053e-09 0 2.247e-09 0 2.25e-09 0.0007 2.253e-09 0 2.447e-09 0 2.45e-09 0.0007 2.453e-09 0 2.647e-09 0 2.65e-09 0.0007 2.653e-09 0 2.847e-09 0 2.85e-09 0.0007 2.853e-09 0 3.047e-09 0 3.05e-09 0.0007 3.053e-09 0 3.247e-09 0 3.25e-09 0.0007 3.253e-09 0 3.447e-09 0 3.45e-09 0.0007 3.453e-09 0 3.647e-09 0 3.65e-09 0.0007 3.653e-09 0 3.847e-09 0 3.85e-09 0.0007 3.853e-09 0 4.047e-09 0 4.05e-09 0.0007 4.053e-09 0 4.247e-09 0 4.25e-09 0.0007 4.253e-09 0 4.447e-09 0 4.45e-09 0.0007 4.453e-09 0 4.647e-09 0 4.65e-09 0.0007 4.653e-09 0 4.847e-09 0 4.85e-09 0.0007 4.853e-09 0 5.047e-09 0 5.05e-09 0.0007 5.053e-09 0 5.247e-09 0 5.25e-09 0.0007 5.253e-09 0 5.447e-09 0 5.45e-09 0.0007 5.453e-09 0 5.647e-09 0 5.65e-09 0.0007 5.653e-09 0 5.847e-09 0 5.85e-09 0.0007 5.853e-09 0 6.047e-09 0 6.05e-09 0.0007 6.053e-09 0 6.247e-09 0 6.25e-09 0.0007 6.253e-09 0 6.447e-09 0 6.45e-09 0.0007 6.453e-09 0 6.647e-09 0 6.65e-09 0.0007 6.653e-09 0 6.847e-09 0 6.85e-09 0.0007 6.853e-09 0 7.047e-09 0 7.05e-09 0.0007 7.053e-09 0 7.247e-09 0 7.25e-09 0.0007 7.253e-09 0 7.447e-09 0 7.45e-09 0.0007 7.453e-09 0 7.647e-09 0 7.65e-09 0.0007 7.653e-09 0 7.847e-09 0 7.85e-09 0.0007 7.853e-09 0 8.047e-09 0 8.05e-09 0.0007 8.053e-09 0 8.247e-09 0 8.25e-09 0.0007 8.253e-09 0 8.447e-09 0 8.45e-09 0.0007 8.453e-09 0 8.647e-09 0 8.65e-09 0.0007 8.653e-09 0 8.847e-09 0 8.85e-09 0.0007 8.853e-09 0 9.047e-09 0 9.05e-09 0.0007 9.053e-09 0 9.247e-09 0 9.25e-09 0.0007 9.253e-09 0 9.447e-09 0 9.45e-09 0.0007 9.453e-09 0 9.647e-09 0 9.65e-09 0.0007 9.653e-09 0 9.847e-09 0 9.85e-09 0.0007 9.853e-09 0 1.0047e-08 0 1.005e-08 0.0007 1.0053e-08 0 1.0247e-08 0 1.025e-08 0.0007 1.0253e-08 0 1.0447e-08 0 1.045e-08 0.0007 1.0453e-08 0 1.0647e-08 0 1.065e-08 0.0007 1.0653e-08 0 1.0847e-08 0 1.085e-08 0.0007 1.0853e-08 0 1.1047e-08 0 1.105e-08 0.0007 1.1053e-08 0 1.1247e-08 0 1.125e-08 0.0007 1.1253e-08 0 1.1447e-08 0 1.145e-08 0.0007 1.1453e-08 0 1.1647e-08 0 1.165e-08 0.0007 1.1653e-08 0 1.1847e-08 0 1.185e-08 0.0007 1.1853e-08 0 1.2047e-08 0 1.205e-08 0.0007 1.2053e-08 0 1.2247e-08 0 1.225e-08 0.0007 1.2253e-08 0 1.2447e-08 0 1.245e-08 0.0007 1.2453e-08 0 1.2647e-08 0 1.265e-08 0.0007 1.2653e-08 0 1.2847e-08 0 1.285e-08 0.0007 1.2853e-08 0 1.3047e-08 0 1.305e-08 0.0007 1.3053e-08 0 1.3247e-08 0 1.325e-08 0.0007 1.3253e-08 0 1.3447e-08 0 1.345e-08 0.0007 1.3453e-08 0 1.3647e-08 0 1.365e-08 0.0007 1.3653e-08 0 1.3847e-08 0 1.385e-08 0.0007 1.3853e-08 0 1.4047e-08 0 1.405e-08 0.0007 1.4053e-08 0 1.4247e-08 0 1.425e-08 0.0007 1.4253e-08 0 1.4447e-08 0 1.445e-08 0.0007 1.4453e-08 0 1.4647e-08 0 1.465e-08 0.0007 1.4653e-08 0 1.4847e-08 0 1.485e-08 0.0007 1.4853e-08 0 1.5047e-08 0 1.505e-08 0.0007 1.5053e-08 0 1.5247e-08 0 1.525e-08 0.0007 1.5253e-08 0 1.5447e-08 0 1.545e-08 0.0007 1.5453e-08 0 1.5647e-08 0 1.565e-08 0.0007 1.5653e-08 0 1.5847e-08 0 1.585e-08 0.0007 1.5853e-08 0 1.6047e-08 0 1.605e-08 0.0007 1.6053e-08 0 1.6247e-08 0 1.625e-08 0.0007 1.6253e-08 0 1.6447e-08 0 1.645e-08 0.0007 1.6453e-08 0 1.6647e-08 0 1.665e-08 0.0007 1.6653e-08 0 1.6847e-08 0 1.685e-08 0.0007 1.6853e-08 0 1.7047e-08 0 1.705e-08 0.0007 1.7053e-08 0 1.7247e-08 0 1.725e-08 0.0007 1.7253e-08 0 1.7447e-08 0 1.745e-08 0.0007 1.7453e-08 0 1.7647e-08 0 1.765e-08 0.0007 1.7653e-08 0 1.7847e-08 0 1.785e-08 0.0007 1.7853e-08 0 1.8047e-08 0 1.805e-08 0.0007 1.8053e-08 0 1.8247e-08 0 1.825e-08 0.0007 1.8253e-08 0 1.8447e-08 0 1.845e-08 0.0007 1.8453e-08 0 1.8647e-08 0 1.865e-08 0.0007 1.8653e-08 0 1.8847e-08 0 1.885e-08 0.0007 1.8853e-08 0 1.9047e-08 0 1.905e-08 0.0007 1.9053e-08 0 1.9247e-08 0 1.925e-08 0.0007 1.9253e-08 0 1.9447e-08 0 1.945e-08 0.0007 1.9453e-08 0 1.9647e-08 0 1.965e-08 0.0007 1.9653e-08 0 1.9847e-08 0 1.985e-08 0.0007 1.9853e-08 0 2.0047e-08 0 2.005e-08 0.0007 2.0053e-08 0 2.0247e-08 0 2.025e-08 0.0007 2.0253e-08 0 2.0447e-08 0 2.045e-08 0.0007 2.0453e-08 0 2.0647e-08 0 2.065e-08 0.0007 2.0653e-08 0 2.0847e-08 0 2.085e-08 0.0007 2.0853e-08 0 2.1047e-08 0 2.105e-08 0.0007 2.1053e-08 0 2.1247e-08 0 2.125e-08 0.0007 2.1253e-08 0 2.1447e-08 0 2.145e-08 0.0007 2.1453e-08 0 2.1647e-08 0 2.165e-08 0.0007 2.1653e-08 0 2.1847e-08 0 2.185e-08 0.0007 2.1853e-08 0 2.2047e-08 0 2.205e-08 0.0007 2.2053e-08 0 2.2247e-08 0 2.225e-08 0.0007 2.2253e-08 0 2.2447e-08 0 2.245e-08 0.0007 2.2453e-08 0 2.2647e-08 0 2.265e-08 0.0007 2.2653e-08 0 2.2847e-08 0 2.285e-08 0.0007 2.2853e-08 0 2.3047e-08 0 2.305e-08 0.0007 2.3053e-08 0 2.3247e-08 0 2.325e-08 0.0007 2.3253e-08 0 2.3447e-08 0 2.345e-08 0.0007 2.3453e-08 0 2.3647e-08 0 2.365e-08 0.0007 2.3653e-08 0 2.3847e-08 0 2.385e-08 0.0007 2.3853e-08 0 2.4047e-08 0 2.405e-08 0.0007 2.4053e-08 0 2.4247e-08 0 2.425e-08 0.0007 2.4253e-08 0 2.4447e-08 0 2.445e-08 0.0007 2.4453e-08 0 2.4647e-08 0 2.465e-08 0.0007 2.4653e-08 0 2.4847e-08 0 2.485e-08 0.0007 2.4853e-08 0 2.5047e-08 0 2.505e-08 0.0007 2.5053e-08 0 2.5247e-08 0 2.525e-08 0.0007 2.5253e-08 0 2.5447e-08 0 2.545e-08 0.0007 2.5453e-08 0 2.5647e-08 0 2.565e-08 0.0007 2.5653e-08 0 2.5847e-08 0 2.585e-08 0.0007 2.5853e-08 0 2.6047e-08 0 2.605e-08 0.0007 2.6053e-08 0 2.6247e-08 0 2.625e-08 0.0007 2.6253e-08 0 2.6447e-08 0 2.645e-08 0.0007 2.6453e-08 0 2.6647e-08 0 2.665e-08 0.0007 2.6653e-08 0 2.6847e-08 0 2.685e-08 0.0007 2.6853e-08 0 2.7047e-08 0 2.705e-08 0.0007 2.7053e-08 0 2.7247e-08 0 2.725e-08 0.0007 2.7253e-08 0 2.7447e-08 0 2.745e-08 0.0007 2.7453e-08 0 2.7647e-08 0 2.765e-08 0.0007 2.7653e-08 0 2.7847e-08 0 2.785e-08 0.0007 2.7853e-08 0 2.8047e-08 0 2.805e-08 0.0007 2.8053e-08 0 2.8247e-08 0 2.825e-08 0.0007 2.8253e-08 0 2.8447e-08 0 2.845e-08 0.0007 2.8453e-08 0 2.8647e-08 0 2.865e-08 0.0007 2.8653e-08 0 2.8847e-08 0 2.885e-08 0.0007 2.8853e-08 0 2.9047e-08 0 2.905e-08 0.0007 2.9053e-08 0 2.9247e-08 0 2.925e-08 0.0007 2.9253e-08 0 2.9447e-08 0 2.945e-08 0.0007 2.9453e-08 0 2.9647e-08 0 2.965e-08 0.0007 2.9653e-08 0 2.9847e-08 0 2.985e-08 0.0007 2.9853e-08 0 3.0047e-08 0 3.005e-08 0.0007 3.0053e-08 0 3.0247e-08 0 3.025e-08 0.0007 3.0253e-08 0 3.0447e-08 0 3.045e-08 0.0007 3.0453e-08 0 3.0647e-08 0 3.065e-08 0.0007 3.0653e-08 0 3.0847e-08 0 3.085e-08 0.0007 3.0853e-08 0 3.1047e-08 0 3.105e-08 0.0007 3.1053e-08 0 3.1247e-08 0 3.125e-08 0.0007 3.1253e-08 0 3.1447e-08 0 3.145e-08 0.0007 3.1453e-08 0 3.1647e-08 0 3.165e-08 0.0007 3.1653e-08 0 3.1847e-08 0 3.185e-08 0.0007 3.1853e-08 0 3.2047e-08 0 3.205e-08 0.0007 3.2053e-08 0 3.2247e-08 0 3.225e-08 0.0007 3.2253e-08 0 3.2447e-08 0 3.245e-08 0.0007 3.2453e-08 0 3.2647e-08 0 3.265e-08 0.0007 3.2653e-08 0 3.2847e-08 0 3.285e-08 0.0007 3.2853e-08 0 3.3047e-08 0 3.305e-08 0.0007 3.3053e-08 0 3.3247e-08 0 3.325e-08 0.0007 3.3253e-08 0 3.3447e-08 0 3.345e-08 0.0007 3.3453e-08 0 3.3647e-08 0 3.365e-08 0.0007 3.3653e-08 0 3.3847e-08 0 3.385e-08 0.0007 3.3853e-08 0 3.4047e-08 0 3.405e-08 0.0007 3.4053e-08 0 3.4247e-08 0 3.425e-08 0.0007 3.4253e-08 0 3.4447e-08 0 3.445e-08 0.0007 3.4453e-08 0 3.4647e-08 0 3.465e-08 0.0007 3.4653e-08 0 3.4847e-08 0 3.485e-08 0.0007 3.4853e-08 0 3.5047e-08 0 3.505e-08 0.0007 3.5053e-08 0 3.5247e-08 0 3.525e-08 0.0007 3.5253e-08 0 3.5447e-08 0 3.545e-08 0.0007 3.5453e-08 0 3.5647e-08 0 3.565e-08 0.0007 3.5653e-08 0 3.5847e-08 0 3.585e-08 0.0007 3.5853e-08 0 3.6047e-08 0 3.605e-08 0.0007 3.6053e-08 0 3.6247e-08 0 3.625e-08 0.0007 3.6253e-08 0 3.6447e-08 0 3.645e-08 0.0007 3.6453e-08 0 3.6647e-08 0 3.665e-08 0.0007 3.6653e-08 0 3.6847e-08 0 3.685e-08 0.0007 3.6853e-08 0 3.7047e-08 0 3.705e-08 0.0007 3.7053e-08 0 3.7247e-08 0 3.725e-08 0.0007 3.7253e-08 0 3.7447e-08 0 3.745e-08 0.0007 3.7453e-08 0 3.7647e-08 0 3.765e-08 0.0007 3.7653e-08 0 3.7847e-08 0 3.785e-08 0.0007 3.7853e-08 0 3.8047e-08 0 3.805e-08 0.0007 3.8053e-08 0 3.8247e-08 0 3.825e-08 0.0007 3.8253e-08 0 3.8447e-08 0 3.845e-08 0.0007 3.8453e-08 0 3.8647e-08 0 3.865e-08 0.0007 3.8653e-08 0 3.8847e-08 0 3.885e-08 0.0007 3.8853e-08 0 3.9047e-08 0 3.905e-08 0.0007 3.9053e-08 0 3.9247e-08 0 3.925e-08 0.0007 3.9253e-08 0 3.9447e-08 0 3.945e-08 0.0007 3.9453e-08 0 3.9647e-08 0 3.965e-08 0.0007 3.9653e-08 0 3.9847e-08 0 3.985e-08 0.0007 3.9853e-08 0 4.0047e-08 0 4.005e-08 0.0007 4.0053e-08 0 4.0247e-08 0 4.025e-08 0.0007 4.0253e-08 0 4.0447e-08 0 4.045e-08 0.0007 4.0453e-08 0 4.0647e-08 0 4.065e-08 0.0007 4.0653e-08 0 4.0847e-08 0 4.085e-08 0.0007 4.0853e-08 0 4.1047e-08 0 4.105e-08 0.0007 4.1053e-08 0 4.1247e-08 0 4.125e-08 0.0007 4.1253e-08 0 4.1447e-08 0 4.145e-08 0.0007 4.1453e-08 0 4.1647e-08 0 4.165e-08 0.0007 4.1653e-08 0 4.1847e-08 0 4.185e-08 0.0007 4.1853e-08 0 4.2047e-08 0 4.205e-08 0.0007 4.2053e-08 0 4.2247e-08 0 4.225e-08 0.0007 4.2253e-08 0 4.2447e-08 0 4.245e-08 0.0007 4.2453e-08 0 4.2647e-08 0 4.265e-08 0.0007 4.2653e-08 0 4.2847e-08 0 4.285e-08 0.0007 4.2853e-08 0 4.3047e-08 0 4.305e-08 0.0007 4.3053e-08 0 4.3247e-08 0 4.325e-08 0.0007 4.3253e-08 0 4.3447e-08 0 4.345e-08 0.0007 4.3453e-08 0 4.3647e-08 0 4.365e-08 0.0007 4.3653e-08 0 4.3847e-08 0 4.385e-08 0.0007 4.3853e-08 0 4.4047e-08 0 4.405e-08 0.0007 4.4053e-08 0 4.4247e-08 0 4.425e-08 0.0007 4.4253e-08 0 4.4447e-08 0 4.445e-08 0.0007 4.4453e-08 0 4.4647e-08 0 4.465e-08 0.0007 4.4653e-08 0 4.4847e-08 0 4.485e-08 0.0007 4.4853e-08 0 4.5047e-08 0 4.505e-08 0.0007 4.5053e-08 0 4.5247e-08 0 4.525e-08 0.0007 4.5253e-08 0 4.5447e-08 0 4.545e-08 0.0007 4.5453e-08 0 4.5647e-08 0 4.565e-08 0.0007 4.5653e-08 0 4.5847e-08 0 4.585e-08 0.0007 4.5853e-08 0 4.6047e-08 0 4.605e-08 0.0007 4.6053e-08 0 4.6247e-08 0 4.625e-08 0.0007 4.6253e-08 0 4.6447e-08 0 4.645e-08 0.0007 4.6453e-08 0 4.6647e-08 0 4.665e-08 0.0007 4.6653e-08 0 4.6847e-08 0 4.685e-08 0.0007 4.6853e-08 0 4.7047e-08 0 4.705e-08 0.0007 4.7053e-08 0 4.7247e-08 0 4.725e-08 0.0007 4.7253e-08 0 4.7447e-08 0 4.745e-08 0.0007 4.7453e-08 0 4.7647e-08 0 4.765e-08 0.0007 4.7653e-08 0 4.7847e-08 0 4.785e-08 0.0007 4.7853e-08 0 4.8047e-08 0 4.805e-08 0.0007 4.8053e-08 0 4.8247e-08 0 4.825e-08 0.0007 4.8253e-08 0 4.8447e-08 0 4.845e-08 0.0007 4.8453e-08 0 4.8647e-08 0 4.865e-08 0.0007 4.8653e-08 0 4.8847e-08 0 4.885e-08 0.0007 4.8853e-08 0 4.9047e-08 0 4.905e-08 0.0007 4.9053e-08 0 4.9247e-08 0 4.925e-08 0.0007 4.9253e-08 0 4.9447e-08 0 4.945e-08 0.0007 4.9453e-08 0 4.9647e-08 0 4.965e-08 0.0007 4.9653e-08 0 4.9847e-08 0 4.985e-08 0.0007 4.9853e-08 0 5.0047e-08 0 5.005e-08 0.0007 5.0053e-08 0 5.0247e-08 0 5.025e-08 0.0007 5.0253e-08 0 5.0447e-08 0 5.045e-08 0.0007 5.0453e-08 0 5.0647e-08 0 5.065e-08 0.0007 5.0653e-08 0 5.0847e-08 0 5.085e-08 0.0007 5.0853e-08 0 5.1047e-08 0 5.105e-08 0.0007 5.1053e-08 0 5.1247e-08 0 5.125e-08 0.0007 5.1253e-08 0 5.1447e-08 0 5.145e-08 0.0007 5.1453e-08 0 5.1647e-08 0 5.165e-08 0.0007 5.1653e-08 0 5.1847e-08 0 5.185e-08 0.0007 5.1853e-08 0 5.2047e-08 0 5.205e-08 0.0007 5.2053e-08 0 5.2247e-08 0 5.225e-08 0.0007 5.2253e-08 0 5.2447e-08 0 5.245e-08 0.0007 5.2453e-08 0 5.2647e-08 0 5.265e-08 0.0007 5.2653e-08 0 5.2847e-08 0 5.285e-08 0.0007 5.2853e-08 0 5.3047e-08 0 5.305e-08 0.0007 5.3053e-08 0 5.3247e-08 0 5.325e-08 0.0007 5.3253e-08 0 5.3447e-08 0 5.345e-08 0.0007 5.3453e-08 0 5.3647e-08 0 5.365e-08 0.0007 5.3653e-08 0 5.3847e-08 0 5.385e-08 0.0007 5.3853e-08 0 5.4047e-08 0 5.405e-08 0.0007 5.4053e-08 0 5.4247e-08 0 5.425e-08 0.0007 5.4253e-08 0 5.4447e-08 0 5.445e-08 0.0007 5.4453e-08 0 5.4647e-08 0 5.465e-08 0.0007 5.4653e-08 0 5.4847e-08 0 5.485e-08 0.0007 5.4853e-08 0 5.5047e-08 0 5.505e-08 0.0007 5.5053e-08 0 5.5247e-08 0 5.525e-08 0.0007 5.5253e-08 0 5.5447e-08 0 5.545e-08 0.0007 5.5453e-08 0 5.5647e-08 0 5.565e-08 0.0007 5.5653e-08 0 5.5847e-08 0 5.585e-08 0.0007 5.5853e-08 0 5.6047e-08 0 5.605e-08 0.0007 5.6053e-08 0 5.6247e-08 0 5.625e-08 0.0007 5.6253e-08 0 5.6447e-08 0 5.645e-08 0.0007 5.6453e-08 0 5.6647e-08 0 5.665e-08 0.0007 5.6653e-08 0 5.6847e-08 0 5.685e-08 0.0007 5.6853e-08 0 5.7047e-08 0 5.705e-08 0.0007 5.7053e-08 0 5.7247e-08 0 5.725e-08 0.0007 5.7253e-08 0 5.7447e-08 0 5.745e-08 0.0007 5.7453e-08 0 5.7647e-08 0 5.765e-08 0.0007 5.7653e-08 0 5.7847e-08 0 5.785e-08 0.0007 5.7853e-08 0 5.8047e-08 0 5.805e-08 0.0007 5.8053e-08 0 5.8247e-08 0 5.825e-08 0.0007 5.8253e-08 0 5.8447e-08 0 5.845e-08 0.0007 5.8453e-08 0 5.8647e-08 0 5.865e-08 0.0007 5.8653e-08 0 5.8847e-08 0 5.885e-08 0.0007 5.8853e-08 0 5.9047e-08 0 5.905e-08 0.0007 5.9053e-08 0 5.9247e-08 0 5.925e-08 0.0007 5.9253e-08 0 5.9447e-08 0 5.945e-08 0.0007 5.9453e-08 0 5.9647e-08 0 5.965e-08 0.0007 5.9653e-08 0 5.9847e-08 0 5.985e-08 0.0007 5.9853e-08 0 6.0047e-08 0 6.005e-08 0.0007 6.0053e-08 0 6.0247e-08 0 6.025e-08 0.0007 6.0253e-08 0 6.0447e-08 0 6.045e-08 0.0007 6.0453e-08 0 6.0647e-08 0 6.065e-08 0.0007 6.0653e-08 0 6.0847e-08 0 6.085e-08 0.0007 6.0853e-08 0 6.1047e-08 0 6.105e-08 0.0007 6.1053e-08 0 6.1247e-08 0 6.125e-08 0.0007 6.1253e-08 0 6.1447e-08 0 6.145e-08 0.0007 6.1453e-08 0 6.1647e-08 0 6.165e-08 0.0007 6.1653e-08 0 6.1847e-08 0 6.185e-08 0.0007 6.1853e-08 0 6.2047e-08 0 6.205e-08 0.0007 6.2053e-08 0 6.2247e-08 0 6.225e-08 0.0007 6.2253e-08 0 6.2447e-08 0 6.245e-08 0.0007 6.2453e-08 0 6.2647e-08 0 6.265e-08 0.0007 6.2653e-08 0 6.2847e-08 0 6.285e-08 0.0007 6.2853e-08 0 6.3047e-08 0 6.305e-08 0.0007 6.3053e-08 0 6.3247e-08 0 6.325e-08 0.0007 6.3253e-08 0 6.3447e-08 0 6.345e-08 0.0007 6.3453e-08 0 6.3647e-08 0 6.365e-08 0.0007 6.3653e-08 0 6.3847e-08 0 6.385e-08 0.0007 6.3853e-08 0 6.4047e-08 0 6.405e-08 0.0007 6.4053e-08 0 6.4247e-08 0 6.425e-08 0.0007 6.4253e-08 0 6.4447e-08 0 6.445e-08 0.0007 6.4453e-08 0 6.4647e-08 0 6.465e-08 0.0007 6.4653e-08 0 6.4847e-08 0 6.485e-08 0.0007 6.4853e-08 0 6.5047e-08 0 6.505e-08 0.0007 6.5053e-08 0 6.5247e-08 0 6.525e-08 0.0007 6.5253e-08 0 6.5447e-08 0 6.545e-08 0.0007 6.5453e-08 0 6.5647e-08 0 6.565e-08 0.0007 6.5653e-08 0 6.5847e-08 0 6.585e-08 0.0007 6.5853e-08 0 6.6047e-08 0 6.605e-08 0.0007 6.6053e-08 0 6.6247e-08 0 6.625e-08 0.0007 6.6253e-08 0 6.6447e-08 0 6.645e-08 0.0007 6.6453e-08 0 6.6647e-08 0 6.665e-08 0.0007 6.6653e-08 0 6.6847e-08 0 6.685e-08 0.0007 6.6853e-08 0 6.7047e-08 0 6.705e-08 0.0007 6.7053e-08 0 6.7247e-08 0 6.725e-08 0.0007 6.7253e-08 0 6.7447e-08 0 6.745e-08 0.0007 6.7453e-08 0 6.7647e-08 0 6.765e-08 0.0007 6.7653e-08 0 6.7847e-08 0 6.785e-08 0.0007 6.7853e-08 0 6.8047e-08 0 6.805e-08 0.0007 6.8053e-08 0 6.8247e-08 0 6.825e-08 0.0007 6.8253e-08 0 6.8447e-08 0 6.845e-08 0.0007 6.8453e-08 0 6.8647e-08 0 6.865e-08 0.0007 6.8653e-08 0 6.8847e-08 0 6.885e-08 0.0007 6.8853e-08 0 6.9047e-08 0 6.905e-08 0.0007 6.9053e-08 0 6.9247e-08 0 6.925e-08 0.0007 6.9253e-08 0 6.9447e-08 0 6.945e-08 0.0007 6.9453e-08 0 6.9647e-08 0 6.965e-08 0.0007 6.9653e-08 0 6.9847e-08 0 6.985e-08 0.0007 6.9853e-08 0 7.0047e-08 0 7.005e-08 0.0007 7.0053e-08 0 7.0247e-08 0 7.025e-08 0.0007 7.0253e-08 0 7.0447e-08 0 7.045e-08 0.0007 7.0453e-08 0 7.0647e-08 0 7.065e-08 0.0007 7.0653e-08 0 7.0847e-08 0 7.085e-08 0.0007 7.0853e-08 0 7.1047e-08 0 7.105e-08 0.0007 7.1053e-08 0 7.1247e-08 0 7.125e-08 0.0007 7.1253e-08 0 7.1447e-08 0 7.145e-08 0.0007 7.1453e-08 0 7.1647e-08 0 7.165e-08 0.0007 7.1653e-08 0 7.1847e-08 0 7.185e-08 0.0007 7.1853e-08 0 7.2047e-08 0 7.205e-08 0.0007 7.2053e-08 0 7.2247e-08 0 7.225e-08 0.0007 7.2253e-08 0 7.2447e-08 0 7.245e-08 0.0007 7.2453e-08 0 7.2647e-08 0 7.265e-08 0.0007 7.2653e-08 0 7.2847e-08 0 7.285e-08 0.0007 7.2853e-08 0 7.3047e-08 0 7.305e-08 0.0007 7.3053e-08 0 7.3247e-08 0 7.325e-08 0.0007 7.3253e-08 0 7.3447e-08 0 7.345e-08 0.0007 7.3453e-08 0 7.3647e-08 0 7.365e-08 0.0007 7.3653e-08 0 7.3847e-08 0 7.385e-08 0.0007 7.3853e-08 0 7.4047e-08 0 7.405e-08 0.0007 7.4053e-08 0 7.4247e-08 0 7.425e-08 0.0007 7.4253e-08 0 7.4447e-08 0 7.445e-08 0.0007 7.4453e-08 0 7.4647e-08 0 7.465e-08 0.0007 7.4653e-08 0 7.4847e-08 0 7.485e-08 0.0007 7.4853e-08 0 7.5047e-08 0 7.505e-08 0.0007 7.5053e-08 0 7.5247e-08 0 7.525e-08 0.0007 7.5253e-08 0 7.5447e-08 0 7.545e-08 0.0007 7.5453e-08 0 7.5647e-08 0 7.565e-08 0.0007 7.5653e-08 0 7.5847e-08 0 7.585e-08 0.0007 7.5853e-08 0 7.6047e-08 0 7.605e-08 0.0007 7.6053e-08 0 7.6247e-08 0 7.625e-08 0.0007 7.6253e-08 0 7.6447e-08 0 7.645e-08 0.0007 7.6453e-08 0 7.6647e-08 0 7.665e-08 0.0007 7.6653e-08 0 7.6847e-08 0 7.685e-08 0.0007 7.6853e-08 0 7.7047e-08 0 7.705e-08 0.0007 7.7053e-08 0 7.7247e-08 0 7.725e-08 0.0007 7.7253e-08 0 7.7447e-08 0 7.745e-08 0.0007 7.7453e-08 0 7.7647e-08 0 7.765e-08 0.0007 7.7653e-08 0 7.7847e-08 0 7.785e-08 0.0007 7.7853e-08 0 7.8047e-08 0 7.805e-08 0.0007 7.8053e-08 0 7.8247e-08 0 7.825e-08 0.0007 7.8253e-08 0 7.8447e-08 0 7.845e-08 0.0007 7.8453e-08 0 7.8647e-08 0 7.865e-08 0.0007 7.8653e-08 0 7.8847e-08 0 7.885e-08 0.0007 7.8853e-08 0 7.9047e-08 0 7.905e-08 0.0007 7.9053e-08 0 7.9247e-08 0 7.925e-08 0.0007 7.9253e-08 0 7.9447e-08 0 7.945e-08 0.0007 7.9453e-08 0 7.9647e-08 0 7.965e-08 0.0007 7.9653e-08 0)
IT00|T 0 T00  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT01|T 0 T01  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT02|T 0 T02  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT03|T 0 T03  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT04|T 0 T04  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT05|T 0 T05  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT06|T 0 T06  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT07|T 0 T07  PWL(0 0 3.7e-11 0 4e-11 0.0021 4.3e-11 0 2.37e-10 0 2.4e-10 0.0021 2.43e-10 0 4.37e-10 0 4.4e-10 0.0021 4.43e-10 0 6.37e-10 0 6.4e-10 0.0021 6.43e-10 0 8.37e-10 0 8.4e-10 0.0021 8.43e-10 0 1.037e-09 0 1.04e-09 0.0021 1.043e-09 0 1.237e-09 0 1.24e-09 0.0021 1.243e-09 0 1.437e-09 0 1.44e-09 0.0021 1.443e-09 0 1.637e-09 0 1.64e-09 0.0021 1.643e-09 0 1.837e-09 0 1.84e-09 0.0021 1.843e-09 0 2.037e-09 0 2.04e-09 0.0021 2.043e-09 0 2.237e-09 0 2.24e-09 0.0021 2.243e-09 0 2.437e-09 0 2.44e-09 0.0021 2.443e-09 0 2.637e-09 0 2.64e-09 0.0021 2.643e-09 0 2.837e-09 0 2.84e-09 0.0021 2.843e-09 0 3.037e-09 0 3.04e-09 0.0021 3.043e-09 0 3.237e-09 0 3.24e-09 0.0021 3.243e-09 0 3.437e-09 0 3.44e-09 0.0021 3.443e-09 0 3.637e-09 0 3.64e-09 0.0021 3.643e-09 0 3.837e-09 0 3.84e-09 0.0021 3.843e-09 0 4.037e-09 0 4.04e-09 0.0021 4.043e-09 0 4.237e-09 0 4.24e-09 0.0021 4.243e-09 0 4.437e-09 0 4.44e-09 0.0021 4.443e-09 0 4.637e-09 0 4.64e-09 0.0021 4.643e-09 0 4.837e-09 0 4.84e-09 0.0021 4.843e-09 0 5.037e-09 0 5.04e-09 0.0021 5.043e-09 0 5.237e-09 0 5.24e-09 0.0021 5.243e-09 0 5.437e-09 0 5.44e-09 0.0021 5.443e-09 0 5.637e-09 0 5.64e-09 0.0021 5.643e-09 0 5.837e-09 0 5.84e-09 0.0021 5.843e-09 0 6.037e-09 0 6.04e-09 0.0021 6.043e-09 0 6.237e-09 0 6.24e-09 0.0021 6.243e-09 0 6.437e-09 0 6.44e-09 0.0021 6.443e-09 0 6.637e-09 0 6.64e-09 0.0021 6.643e-09 0 6.837e-09 0 6.84e-09 0.0021 6.843e-09 0 7.037e-09 0 7.04e-09 0.0021 7.043e-09 0 7.237e-09 0 7.24e-09 0.0021 7.243e-09 0 7.437e-09 0 7.44e-09 0.0021 7.443e-09 0 7.637e-09 0 7.64e-09 0.0021 7.643e-09 0 7.837e-09 0 7.84e-09 0.0021 7.843e-09 0 8.037e-09 0 8.04e-09 0.0021 8.043e-09 0 8.237e-09 0 8.24e-09 0.0021 8.243e-09 0 8.437e-09 0 8.44e-09 0.0021 8.443e-09 0 8.637e-09 0 8.64e-09 0.0021 8.643e-09 0 8.837e-09 0 8.84e-09 0.0021 8.843e-09 0 9.037e-09 0 9.04e-09 0.0021 9.043e-09 0 9.237e-09 0 9.24e-09 0.0021 9.243e-09 0 9.437e-09 0 9.44e-09 0.0021 9.443e-09 0 9.637e-09 0 9.64e-09 0.0021 9.643e-09 0 9.837e-09 0 9.84e-09 0.0021 9.843e-09 0 1.0037e-08 0 1.004e-08 0.0021 1.0043e-08 0 1.0237e-08 0 1.024e-08 0.0021 1.0243e-08 0 1.0437e-08 0 1.044e-08 0.0021 1.0443e-08 0 1.0637e-08 0 1.064e-08 0.0021 1.0643e-08 0 1.0837e-08 0 1.084e-08 0.0021 1.0843e-08 0 1.1037e-08 0 1.104e-08 0.0021 1.1043e-08 0 1.1237e-08 0 1.124e-08 0.0021 1.1243e-08 0 1.1437e-08 0 1.144e-08 0.0021 1.1443e-08 0 1.1637e-08 0 1.164e-08 0.0021 1.1643e-08 0 1.1837e-08 0 1.184e-08 0.0021 1.1843e-08 0 1.2037e-08 0 1.204e-08 0.0021 1.2043e-08 0 1.2237e-08 0 1.224e-08 0.0021 1.2243e-08 0 1.2437e-08 0 1.244e-08 0.0021 1.2443e-08 0 1.2637e-08 0 1.264e-08 0.0021 1.2643e-08 0 1.2837e-08 0 1.284e-08 0.0021 1.2843e-08 0 1.3037e-08 0 1.304e-08 0.0021 1.3043e-08 0 1.3237e-08 0 1.324e-08 0.0021 1.3243e-08 0 1.3437e-08 0 1.344e-08 0.0021 1.3443e-08 0 1.3637e-08 0 1.364e-08 0.0021 1.3643e-08 0 1.3837e-08 0 1.384e-08 0.0021 1.3843e-08 0 1.4037e-08 0 1.404e-08 0.0021 1.4043e-08 0 1.4237e-08 0 1.424e-08 0.0021 1.4243e-08 0 1.4437e-08 0 1.444e-08 0.0021 1.4443e-08 0 1.4637e-08 0 1.464e-08 0.0021 1.4643e-08 0 1.4837e-08 0 1.484e-08 0.0021 1.4843e-08 0 1.5037e-08 0 1.504e-08 0.0021 1.5043e-08 0 1.5237e-08 0 1.524e-08 0.0021 1.5243e-08 0 1.5437e-08 0 1.544e-08 0.0021 1.5443e-08 0 1.5637e-08 0 1.564e-08 0.0021 1.5643e-08 0 1.5837e-08 0 1.584e-08 0.0021 1.5843e-08 0 1.6037e-08 0 1.604e-08 0.0021 1.6043e-08 0 1.6237e-08 0 1.624e-08 0.0021 1.6243e-08 0 1.6437e-08 0 1.644e-08 0.0021 1.6443e-08 0 1.6637e-08 0 1.664e-08 0.0021 1.6643e-08 0 1.6837e-08 0 1.684e-08 0.0021 1.6843e-08 0 1.7037e-08 0 1.704e-08 0.0021 1.7043e-08 0 1.7237e-08 0 1.724e-08 0.0021 1.7243e-08 0 1.7437e-08 0 1.744e-08 0.0021 1.7443e-08 0 1.7637e-08 0 1.764e-08 0.0021 1.7643e-08 0 1.7837e-08 0 1.784e-08 0.0021 1.7843e-08 0 1.8037e-08 0 1.804e-08 0.0021 1.8043e-08 0 1.8237e-08 0 1.824e-08 0.0021 1.8243e-08 0 1.8437e-08 0 1.844e-08 0.0021 1.8443e-08 0 1.8637e-08 0 1.864e-08 0.0021 1.8643e-08 0 1.8837e-08 0 1.884e-08 0.0021 1.8843e-08 0 1.9037e-08 0 1.904e-08 0.0021 1.9043e-08 0 1.9237e-08 0 1.924e-08 0.0021 1.9243e-08 0 1.9437e-08 0 1.944e-08 0.0021 1.9443e-08 0 1.9637e-08 0 1.964e-08 0.0021 1.9643e-08 0 1.9837e-08 0 1.984e-08 0.0021 1.9843e-08 0 2.0037e-08 0 2.004e-08 0.0021 2.0043e-08 0 2.0237e-08 0 2.024e-08 0.0021 2.0243e-08 0 2.0437e-08 0 2.044e-08 0.0021 2.0443e-08 0 2.0637e-08 0 2.064e-08 0.0021 2.0643e-08 0 2.0837e-08 0 2.084e-08 0.0021 2.0843e-08 0 2.1037e-08 0 2.104e-08 0.0021 2.1043e-08 0 2.1237e-08 0 2.124e-08 0.0021 2.1243e-08 0 2.1437e-08 0 2.144e-08 0.0021 2.1443e-08 0 2.1637e-08 0 2.164e-08 0.0021 2.1643e-08 0 2.1837e-08 0 2.184e-08 0.0021 2.1843e-08 0 2.2037e-08 0 2.204e-08 0.0021 2.2043e-08 0 2.2237e-08 0 2.224e-08 0.0021 2.2243e-08 0 2.2437e-08 0 2.244e-08 0.0021 2.2443e-08 0 2.2637e-08 0 2.264e-08 0.0021 2.2643e-08 0 2.2837e-08 0 2.284e-08 0.0021 2.2843e-08 0 2.3037e-08 0 2.304e-08 0.0021 2.3043e-08 0 2.3237e-08 0 2.324e-08 0.0021 2.3243e-08 0 2.3437e-08 0 2.344e-08 0.0021 2.3443e-08 0 2.3637e-08 0 2.364e-08 0.0021 2.3643e-08 0 2.3837e-08 0 2.384e-08 0.0021 2.3843e-08 0 2.4037e-08 0 2.404e-08 0.0021 2.4043e-08 0 2.4237e-08 0 2.424e-08 0.0021 2.4243e-08 0 2.4437e-08 0 2.444e-08 0.0021 2.4443e-08 0 2.4637e-08 0 2.464e-08 0.0021 2.4643e-08 0 2.4837e-08 0 2.484e-08 0.0021 2.4843e-08 0 2.5037e-08 0 2.504e-08 0.0021 2.5043e-08 0 2.5237e-08 0 2.524e-08 0.0021 2.5243e-08 0 2.5437e-08 0 2.544e-08 0.0021 2.5443e-08 0 2.5637e-08 0 2.564e-08 0.0021 2.5643e-08 0 2.5837e-08 0 2.584e-08 0.0021 2.5843e-08 0 2.6037e-08 0 2.604e-08 0.0021 2.6043e-08 0 2.6237e-08 0 2.624e-08 0.0021 2.6243e-08 0 2.6437e-08 0 2.644e-08 0.0021 2.6443e-08 0 2.6637e-08 0 2.664e-08 0.0021 2.6643e-08 0 2.6837e-08 0 2.684e-08 0.0021 2.6843e-08 0 2.7037e-08 0 2.704e-08 0.0021 2.7043e-08 0 2.7237e-08 0 2.724e-08 0.0021 2.7243e-08 0 2.7437e-08 0 2.744e-08 0.0021 2.7443e-08 0 2.7637e-08 0 2.764e-08 0.0021 2.7643e-08 0 2.7837e-08 0 2.784e-08 0.0021 2.7843e-08 0 2.8037e-08 0 2.804e-08 0.0021 2.8043e-08 0 2.8237e-08 0 2.824e-08 0.0021 2.8243e-08 0 2.8437e-08 0 2.844e-08 0.0021 2.8443e-08 0 2.8637e-08 0 2.864e-08 0.0021 2.8643e-08 0 2.8837e-08 0 2.884e-08 0.0021 2.8843e-08 0 2.9037e-08 0 2.904e-08 0.0021 2.9043e-08 0 2.9237e-08 0 2.924e-08 0.0021 2.9243e-08 0 2.9437e-08 0 2.944e-08 0.0021 2.9443e-08 0 2.9637e-08 0 2.964e-08 0.0021 2.9643e-08 0 2.9837e-08 0 2.984e-08 0.0021 2.9843e-08 0 3.0037e-08 0 3.004e-08 0.0021 3.0043e-08 0 3.0237e-08 0 3.024e-08 0.0021 3.0243e-08 0 3.0437e-08 0 3.044e-08 0.0021 3.0443e-08 0 3.0637e-08 0 3.064e-08 0.0021 3.0643e-08 0 3.0837e-08 0 3.084e-08 0.0021 3.0843e-08 0 3.1037e-08 0 3.104e-08 0.0021 3.1043e-08 0 3.1237e-08 0 3.124e-08 0.0021 3.1243e-08 0 3.1437e-08 0 3.144e-08 0.0021 3.1443e-08 0 3.1637e-08 0 3.164e-08 0.0021 3.1643e-08 0 3.1837e-08 0 3.184e-08 0.0021 3.1843e-08 0 3.2037e-08 0 3.204e-08 0.0021 3.2043e-08 0 3.2237e-08 0 3.224e-08 0.0021 3.2243e-08 0 3.2437e-08 0 3.244e-08 0.0021 3.2443e-08 0 3.2637e-08 0 3.264e-08 0.0021 3.2643e-08 0 3.2837e-08 0 3.284e-08 0.0021 3.2843e-08 0 3.3037e-08 0 3.304e-08 0.0021 3.3043e-08 0 3.3237e-08 0 3.324e-08 0.0021 3.3243e-08 0 3.3437e-08 0 3.344e-08 0.0021 3.3443e-08 0 3.3637e-08 0 3.364e-08 0.0021 3.3643e-08 0 3.3837e-08 0 3.384e-08 0.0021 3.3843e-08 0 3.4037e-08 0 3.404e-08 0.0021 3.4043e-08 0 3.4237e-08 0 3.424e-08 0.0021 3.4243e-08 0 3.4437e-08 0 3.444e-08 0.0021 3.4443e-08 0 3.4637e-08 0 3.464e-08 0.0021 3.4643e-08 0 3.4837e-08 0 3.484e-08 0.0021 3.4843e-08 0 3.5037e-08 0 3.504e-08 0.0021 3.5043e-08 0 3.5237e-08 0 3.524e-08 0.0021 3.5243e-08 0 3.5437e-08 0 3.544e-08 0.0021 3.5443e-08 0 3.5637e-08 0 3.564e-08 0.0021 3.5643e-08 0 3.5837e-08 0 3.584e-08 0.0021 3.5843e-08 0 3.6037e-08 0 3.604e-08 0.0021 3.6043e-08 0 3.6237e-08 0 3.624e-08 0.0021 3.6243e-08 0 3.6437e-08 0 3.644e-08 0.0021 3.6443e-08 0 3.6637e-08 0 3.664e-08 0.0021 3.6643e-08 0 3.6837e-08 0 3.684e-08 0.0021 3.6843e-08 0 3.7037e-08 0 3.704e-08 0.0021 3.7043e-08 0 3.7237e-08 0 3.724e-08 0.0021 3.7243e-08 0 3.7437e-08 0 3.744e-08 0.0021 3.7443e-08 0 3.7637e-08 0 3.764e-08 0.0021 3.7643e-08 0 3.7837e-08 0 3.784e-08 0.0021 3.7843e-08 0 3.8037e-08 0 3.804e-08 0.0021 3.8043e-08 0 3.8237e-08 0 3.824e-08 0.0021 3.8243e-08 0 3.8437e-08 0 3.844e-08 0.0021 3.8443e-08 0 3.8637e-08 0 3.864e-08 0.0021 3.8643e-08 0 3.8837e-08 0 3.884e-08 0.0021 3.8843e-08 0 3.9037e-08 0 3.904e-08 0.0021 3.9043e-08 0 3.9237e-08 0 3.924e-08 0.0021 3.9243e-08 0 3.9437e-08 0 3.944e-08 0.0021 3.9443e-08 0 3.9637e-08 0 3.964e-08 0.0021 3.9643e-08 0 3.9837e-08 0 3.984e-08 0.0021 3.9843e-08 0 4.0037e-08 0 4.004e-08 0.0021 4.0043e-08 0 4.0237e-08 0 4.024e-08 0.0021 4.0243e-08 0 4.0437e-08 0 4.044e-08 0.0021 4.0443e-08 0 4.0637e-08 0 4.064e-08 0.0021 4.0643e-08 0 4.0837e-08 0 4.084e-08 0.0021 4.0843e-08 0 4.1037e-08 0 4.104e-08 0.0021 4.1043e-08 0 4.1237e-08 0 4.124e-08 0.0021 4.1243e-08 0 4.1437e-08 0 4.144e-08 0.0021 4.1443e-08 0 4.1637e-08 0 4.164e-08 0.0021 4.1643e-08 0 4.1837e-08 0 4.184e-08 0.0021 4.1843e-08 0 4.2037e-08 0 4.204e-08 0.0021 4.2043e-08 0 4.2237e-08 0 4.224e-08 0.0021 4.2243e-08 0 4.2437e-08 0 4.244e-08 0.0021 4.2443e-08 0 4.2637e-08 0 4.264e-08 0.0021 4.2643e-08 0 4.2837e-08 0 4.284e-08 0.0021 4.2843e-08 0 4.3037e-08 0 4.304e-08 0.0021 4.3043e-08 0 4.3237e-08 0 4.324e-08 0.0021 4.3243e-08 0 4.3437e-08 0 4.344e-08 0.0021 4.3443e-08 0 4.3637e-08 0 4.364e-08 0.0021 4.3643e-08 0 4.3837e-08 0 4.384e-08 0.0021 4.3843e-08 0 4.4037e-08 0 4.404e-08 0.0021 4.4043e-08 0 4.4237e-08 0 4.424e-08 0.0021 4.4243e-08 0 4.4437e-08 0 4.444e-08 0.0021 4.4443e-08 0 4.4637e-08 0 4.464e-08 0.0021 4.4643e-08 0 4.4837e-08 0 4.484e-08 0.0021 4.4843e-08 0 4.5037e-08 0 4.504e-08 0.0021 4.5043e-08 0 4.5237e-08 0 4.524e-08 0.0021 4.5243e-08 0 4.5437e-08 0 4.544e-08 0.0021 4.5443e-08 0 4.5637e-08 0 4.564e-08 0.0021 4.5643e-08 0 4.5837e-08 0 4.584e-08 0.0021 4.5843e-08 0 4.6037e-08 0 4.604e-08 0.0021 4.6043e-08 0 4.6237e-08 0 4.624e-08 0.0021 4.6243e-08 0 4.6437e-08 0 4.644e-08 0.0021 4.6443e-08 0 4.6637e-08 0 4.664e-08 0.0021 4.6643e-08 0 4.6837e-08 0 4.684e-08 0.0021 4.6843e-08 0 4.7037e-08 0 4.704e-08 0.0021 4.7043e-08 0 4.7237e-08 0 4.724e-08 0.0021 4.7243e-08 0 4.7437e-08 0 4.744e-08 0.0021 4.7443e-08 0 4.7637e-08 0 4.764e-08 0.0021 4.7643e-08 0 4.7837e-08 0 4.784e-08 0.0021 4.7843e-08 0 4.8037e-08 0 4.804e-08 0.0021 4.8043e-08 0 4.8237e-08 0 4.824e-08 0.0021 4.8243e-08 0 4.8437e-08 0 4.844e-08 0.0021 4.8443e-08 0 4.8637e-08 0 4.864e-08 0.0021 4.8643e-08 0 4.8837e-08 0 4.884e-08 0.0021 4.8843e-08 0 4.9037e-08 0 4.904e-08 0.0021 4.9043e-08 0 4.9237e-08 0 4.924e-08 0.0021 4.9243e-08 0 4.9437e-08 0 4.944e-08 0.0021 4.9443e-08 0 4.9637e-08 0 4.964e-08 0.0021 4.9643e-08 0 4.9837e-08 0 4.984e-08 0.0021 4.9843e-08 0 5.0037e-08 0 5.004e-08 0.0021 5.0043e-08 0 5.0237e-08 0 5.024e-08 0.0021 5.0243e-08 0 5.0437e-08 0 5.044e-08 0.0021 5.0443e-08 0 5.0637e-08 0 5.064e-08 0.0021 5.0643e-08 0 5.0837e-08 0 5.084e-08 0.0021 5.0843e-08 0 5.1037e-08 0 5.104e-08 0.0021 5.1043e-08 0 5.1237e-08 0 5.124e-08 0.0021 5.1243e-08 0 5.1437e-08 0 5.144e-08 0.0021 5.1443e-08 0 5.1637e-08 0 5.164e-08 0.0021 5.1643e-08 0 5.1837e-08 0 5.184e-08 0.0021 5.1843e-08 0 5.2037e-08 0 5.204e-08 0.0021 5.2043e-08 0 5.2237e-08 0 5.224e-08 0.0021 5.2243e-08 0 5.2437e-08 0 5.244e-08 0.0021 5.2443e-08 0 5.2637e-08 0 5.264e-08 0.0021 5.2643e-08 0 5.2837e-08 0 5.284e-08 0.0021 5.2843e-08 0 5.3037e-08 0 5.304e-08 0.0021 5.3043e-08 0 5.3237e-08 0 5.324e-08 0.0021 5.3243e-08 0 5.3437e-08 0 5.344e-08 0.0021 5.3443e-08 0 5.3637e-08 0 5.364e-08 0.0021 5.3643e-08 0 5.3837e-08 0 5.384e-08 0.0021 5.3843e-08 0 5.4037e-08 0 5.404e-08 0.0021 5.4043e-08 0 5.4237e-08 0 5.424e-08 0.0021 5.4243e-08 0 5.4437e-08 0 5.444e-08 0.0021 5.4443e-08 0 5.4637e-08 0 5.464e-08 0.0021 5.4643e-08 0 5.4837e-08 0 5.484e-08 0.0021 5.4843e-08 0 5.5037e-08 0 5.504e-08 0.0021 5.5043e-08 0 5.5237e-08 0 5.524e-08 0.0021 5.5243e-08 0 5.5437e-08 0 5.544e-08 0.0021 5.5443e-08 0 5.5637e-08 0 5.564e-08 0.0021 5.5643e-08 0 5.5837e-08 0 5.584e-08 0.0021 5.5843e-08 0 5.6037e-08 0 5.604e-08 0.0021 5.6043e-08 0 5.6237e-08 0 5.624e-08 0.0021 5.6243e-08 0 5.6437e-08 0 5.644e-08 0.0021 5.6443e-08 0 5.6637e-08 0 5.664e-08 0.0021 5.6643e-08 0 5.6837e-08 0 5.684e-08 0.0021 5.6843e-08 0 5.7037e-08 0 5.704e-08 0.0021 5.7043e-08 0 5.7237e-08 0 5.724e-08 0.0021 5.7243e-08 0 5.7437e-08 0 5.744e-08 0.0021 5.7443e-08 0 5.7637e-08 0 5.764e-08 0.0021 5.7643e-08 0 5.7837e-08 0 5.784e-08 0.0021 5.7843e-08 0 5.8037e-08 0 5.804e-08 0.0021 5.8043e-08 0 5.8237e-08 0 5.824e-08 0.0021 5.8243e-08 0 5.8437e-08 0 5.844e-08 0.0021 5.8443e-08 0 5.8637e-08 0 5.864e-08 0.0021 5.8643e-08 0 5.8837e-08 0 5.884e-08 0.0021 5.8843e-08 0 5.9037e-08 0 5.904e-08 0.0021 5.9043e-08 0 5.9237e-08 0 5.924e-08 0.0021 5.9243e-08 0 5.9437e-08 0 5.944e-08 0.0021 5.9443e-08 0 5.9637e-08 0 5.964e-08 0.0021 5.9643e-08 0 5.9837e-08 0 5.984e-08 0.0021 5.9843e-08 0 6.0037e-08 0 6.004e-08 0.0021 6.0043e-08 0 6.0237e-08 0 6.024e-08 0.0021 6.0243e-08 0 6.0437e-08 0 6.044e-08 0.0021 6.0443e-08 0 6.0637e-08 0 6.064e-08 0.0021 6.0643e-08 0 6.0837e-08 0 6.084e-08 0.0021 6.0843e-08 0 6.1037e-08 0 6.104e-08 0.0021 6.1043e-08 0 6.1237e-08 0 6.124e-08 0.0021 6.1243e-08 0 6.1437e-08 0 6.144e-08 0.0021 6.1443e-08 0 6.1637e-08 0 6.164e-08 0.0021 6.1643e-08 0 6.1837e-08 0 6.184e-08 0.0021 6.1843e-08 0 6.2037e-08 0 6.204e-08 0.0021 6.2043e-08 0 6.2237e-08 0 6.224e-08 0.0021 6.2243e-08 0 6.2437e-08 0 6.244e-08 0.0021 6.2443e-08 0 6.2637e-08 0 6.264e-08 0.0021 6.2643e-08 0 6.2837e-08 0 6.284e-08 0.0021 6.2843e-08 0 6.3037e-08 0 6.304e-08 0.0021 6.3043e-08 0 6.3237e-08 0 6.324e-08 0.0021 6.3243e-08 0 6.3437e-08 0 6.344e-08 0.0021 6.3443e-08 0 6.3637e-08 0 6.364e-08 0.0021 6.3643e-08 0 6.3837e-08 0 6.384e-08 0.0021 6.3843e-08 0 6.4037e-08 0 6.404e-08 0.0021 6.4043e-08 0 6.4237e-08 0 6.424e-08 0.0021 6.4243e-08 0 6.4437e-08 0 6.444e-08 0.0021 6.4443e-08 0 6.4637e-08 0 6.464e-08 0.0021 6.4643e-08 0 6.4837e-08 0 6.484e-08 0.0021 6.4843e-08 0 6.5037e-08 0 6.504e-08 0.0021 6.5043e-08 0 6.5237e-08 0 6.524e-08 0.0021 6.5243e-08 0 6.5437e-08 0 6.544e-08 0.0021 6.5443e-08 0 6.5637e-08 0 6.564e-08 0.0021 6.5643e-08 0 6.5837e-08 0 6.584e-08 0.0021 6.5843e-08 0 6.6037e-08 0 6.604e-08 0.0021 6.6043e-08 0 6.6237e-08 0 6.624e-08 0.0021 6.6243e-08 0 6.6437e-08 0 6.644e-08 0.0021 6.6443e-08 0 6.6637e-08 0 6.664e-08 0.0021 6.6643e-08 0 6.6837e-08 0 6.684e-08 0.0021 6.6843e-08 0 6.7037e-08 0 6.704e-08 0.0021 6.7043e-08 0 6.7237e-08 0 6.724e-08 0.0021 6.7243e-08 0 6.7437e-08 0 6.744e-08 0.0021 6.7443e-08 0 6.7637e-08 0 6.764e-08 0.0021 6.7643e-08 0 6.7837e-08 0 6.784e-08 0.0021 6.7843e-08 0 6.8037e-08 0 6.804e-08 0.0021 6.8043e-08 0 6.8237e-08 0 6.824e-08 0.0021 6.8243e-08 0 6.8437e-08 0 6.844e-08 0.0021 6.8443e-08 0 6.8637e-08 0 6.864e-08 0.0021 6.8643e-08 0 6.8837e-08 0 6.884e-08 0.0021 6.8843e-08 0 6.9037e-08 0 6.904e-08 0.0021 6.9043e-08 0 6.9237e-08 0 6.924e-08 0.0021 6.9243e-08 0 6.9437e-08 0 6.944e-08 0.0021 6.9443e-08 0 6.9637e-08 0 6.964e-08 0.0021 6.9643e-08 0 6.9837e-08 0 6.984e-08 0.0021 6.9843e-08 0 7.0037e-08 0 7.004e-08 0.0021 7.0043e-08 0 7.0237e-08 0 7.024e-08 0.0021 7.0243e-08 0 7.0437e-08 0 7.044e-08 0.0021 7.0443e-08 0 7.0637e-08 0 7.064e-08 0.0021 7.0643e-08 0 7.0837e-08 0 7.084e-08 0.0021 7.0843e-08 0 7.1037e-08 0 7.104e-08 0.0021 7.1043e-08 0 7.1237e-08 0 7.124e-08 0.0021 7.1243e-08 0 7.1437e-08 0 7.144e-08 0.0021 7.1443e-08 0 7.1637e-08 0 7.164e-08 0.0021 7.1643e-08 0 7.1837e-08 0 7.184e-08 0.0021 7.1843e-08 0 7.2037e-08 0 7.204e-08 0.0021 7.2043e-08 0 7.2237e-08 0 7.224e-08 0.0021 7.2243e-08 0 7.2437e-08 0 7.244e-08 0.0021 7.2443e-08 0 7.2637e-08 0 7.264e-08 0.0021 7.2643e-08 0 7.2837e-08 0 7.284e-08 0.0021 7.2843e-08 0 7.3037e-08 0 7.304e-08 0.0021 7.3043e-08 0 7.3237e-08 0 7.324e-08 0.0021 7.3243e-08 0 7.3437e-08 0 7.344e-08 0.0021 7.3443e-08 0 7.3637e-08 0 7.364e-08 0.0021 7.3643e-08 0 7.3837e-08 0 7.384e-08 0.0021 7.3843e-08 0 7.4037e-08 0 7.404e-08 0.0021 7.4043e-08 0 7.4237e-08 0 7.424e-08 0.0021 7.4243e-08 0 7.4437e-08 0 7.444e-08 0.0021 7.4443e-08 0 7.4637e-08 0 7.464e-08 0.0021 7.4643e-08 0 7.4837e-08 0 7.484e-08 0.0021 7.4843e-08 0 7.5037e-08 0 7.504e-08 0.0021 7.5043e-08 0 7.5237e-08 0 7.524e-08 0.0021 7.5243e-08 0 7.5437e-08 0 7.544e-08 0.0021 7.5443e-08 0 7.5637e-08 0 7.564e-08 0.0021 7.5643e-08 0 7.5837e-08 0 7.584e-08 0.0021 7.5843e-08 0 7.6037e-08 0 7.604e-08 0.0021 7.6043e-08 0 7.6237e-08 0 7.624e-08 0.0021 7.6243e-08 0 7.6437e-08 0 7.644e-08 0.0021 7.6443e-08 0 7.6637e-08 0 7.664e-08 0.0021 7.6643e-08 0 7.6837e-08 0 7.684e-08 0.0021 7.6843e-08 0 7.7037e-08 0 7.704e-08 0.0021 7.7043e-08 0 7.7237e-08 0 7.724e-08 0.0021 7.7243e-08 0 7.7437e-08 0 7.744e-08 0.0021 7.7443e-08 0 7.7637e-08 0 7.764e-08 0.0021 7.7643e-08 0 7.7837e-08 0 7.784e-08 0.0021 7.7843e-08 0 7.8037e-08 0 7.804e-08 0.0021 7.8043e-08 0 7.8237e-08 0 7.824e-08 0.0021 7.8243e-08 0 7.8437e-08 0 7.844e-08 0.0021 7.8443e-08 0 7.8637e-08 0 7.864e-08 0.0021 7.8643e-08 0 7.8837e-08 0 7.884e-08 0.0021 7.8843e-08 0 7.9037e-08 0 7.904e-08 0.0021 7.9043e-08 0 7.9237e-08 0 7.924e-08 0.0021 7.9243e-08 0 7.9437e-08 0 7.944e-08 0.0021 7.9443e-08 0 7.9637e-08 0 7.964e-08 0.0021 7.9643e-08 0)
IT10|T 0 T10  PWL(0 0 2.7e-11 0 3e-11 0.0007 3.3e-11 0 2.27e-10 0 2.3e-10 0.0007 2.33e-10 0 4.27e-10 0 4.3e-10 0.0007 4.33e-10 0 6.27e-10 0 6.3e-10 0.0007 6.33e-10 0 8.27e-10 0 8.3e-10 0.0007 8.33e-10 0 1.027e-09 0 1.03e-09 0.0007 1.033e-09 0 1.227e-09 0 1.23e-09 0.0007 1.233e-09 0 1.427e-09 0 1.43e-09 0.0007 1.433e-09 0 1.627e-09 0 1.63e-09 0.0007 1.633e-09 0 1.827e-09 0 1.83e-09 0.0007 1.833e-09 0 2.027e-09 0 2.03e-09 0.0007 2.033e-09 0 2.227e-09 0 2.23e-09 0.0007 2.233e-09 0 2.427e-09 0 2.43e-09 0.0007 2.433e-09 0 2.627e-09 0 2.63e-09 0.0007 2.633e-09 0 2.827e-09 0 2.83e-09 0.0007 2.833e-09 0 3.027e-09 0 3.03e-09 0.0007 3.033e-09 0 3.227e-09 0 3.23e-09 0.0007 3.233e-09 0 3.427e-09 0 3.43e-09 0.0007 3.433e-09 0 3.627e-09 0 3.63e-09 0.0007 3.633e-09 0 3.827e-09 0 3.83e-09 0.0007 3.833e-09 0 4.027e-09 0 4.03e-09 0.0007 4.033e-09 0 4.227e-09 0 4.23e-09 0.0007 4.233e-09 0 4.427e-09 0 4.43e-09 0.0007 4.433e-09 0 4.627e-09 0 4.63e-09 0.0007 4.633e-09 0 4.827e-09 0 4.83e-09 0.0007 4.833e-09 0 5.027e-09 0 5.03e-09 0.0007 5.033e-09 0 5.227e-09 0 5.23e-09 0.0007 5.233e-09 0 5.427e-09 0 5.43e-09 0.0007 5.433e-09 0 5.627e-09 0 5.63e-09 0.0007 5.633e-09 0 5.827e-09 0 5.83e-09 0.0007 5.833e-09 0 6.027e-09 0 6.03e-09 0.0007 6.033e-09 0 6.227e-09 0 6.23e-09 0.0007 6.233e-09 0 6.427e-09 0 6.43e-09 0.0007 6.433e-09 0 6.627e-09 0 6.63e-09 0.0007 6.633e-09 0 6.827e-09 0 6.83e-09 0.0007 6.833e-09 0 7.027e-09 0 7.03e-09 0.0007 7.033e-09 0 7.227e-09 0 7.23e-09 0.0007 7.233e-09 0 7.427e-09 0 7.43e-09 0.0007 7.433e-09 0 7.627e-09 0 7.63e-09 0.0007 7.633e-09 0 7.827e-09 0 7.83e-09 0.0007 7.833e-09 0 8.027e-09 0 8.03e-09 0.0007 8.033e-09 0 8.227e-09 0 8.23e-09 0.0007 8.233e-09 0 8.427e-09 0 8.43e-09 0.0007 8.433e-09 0 8.627e-09 0 8.63e-09 0.0007 8.633e-09 0 8.827e-09 0 8.83e-09 0.0007 8.833e-09 0 9.027e-09 0 9.03e-09 0.0007 9.033e-09 0 9.227e-09 0 9.23e-09 0.0007 9.233e-09 0 9.427e-09 0 9.43e-09 0.0007 9.433e-09 0 9.627e-09 0 9.63e-09 0.0007 9.633e-09 0 9.827e-09 0 9.83e-09 0.0007 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0007 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0007 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0007 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0007 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0007 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0007 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0007 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0007 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0007 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0007 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0007 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0007 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0007 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0007 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0007 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0007 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0007 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0007 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0007 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0007 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0007 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0007 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0007 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0007 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0007 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0007 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0007 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0007 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0007 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0007 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0007 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0007 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0007 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0007 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0007 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0007 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0007 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0007 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0007 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0007 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0007 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0007 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0007 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0007 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0007 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0007 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0007 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0007 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0007 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0007 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0007 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0007 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0007 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0007 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0007 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0007 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0007 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0007 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0007 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0007 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0007 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0007 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0007 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0007 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0007 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0007 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0007 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0007 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0007 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0007 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0007 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0007 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0007 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0007 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0007 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0007 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0007 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0007 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0007 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0007 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0007 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0007 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0007 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0007 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0007 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0007 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0007 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0007 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0007 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0007 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0007 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0007 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0007 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0007 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0007 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0007 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0007 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0007 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0007 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0007 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0007 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0007 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0007 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0007 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0007 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0007 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0007 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0007 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0007 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0007 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0007 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0007 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0007 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0007 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0007 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0007 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0007 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0007 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0007 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0007 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0007 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0007 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0007 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0007 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0007 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0007 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0007 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0007 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0007 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0007 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0007 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0007 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0007 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0007 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0007 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0007 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0007 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0007 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0007 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0007 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0007 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0007 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0007 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0007 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0007 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0007 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0007 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0007 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0007 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0007 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0007 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0007 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0007 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0007 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0007 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0007 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0007 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0007 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0007 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0007 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0007 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0007 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0007 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0007 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0007 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0007 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0007 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0007 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0007 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0007 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0007 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0007 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0007 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0007 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0007 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0007 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0007 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0007 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0007 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0007 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0007 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0007 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0007 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0007 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0007 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0007 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0007 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0007 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0007 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0007 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0007 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0007 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0007 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0007 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0007 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0007 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0007 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0007 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0007 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0007 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0007 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0007 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0007 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0007 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0007 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0007 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0007 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0007 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0007 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0007 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0007 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0007 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0007 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0007 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0007 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0007 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0007 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0007 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0007 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0007 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0007 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0007 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0007 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0007 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0007 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0007 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0007 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0007 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0007 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0007 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0007 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0007 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0007 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0007 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0007 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0007 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0007 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0007 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0007 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0007 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0007 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0007 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0007 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0007 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0007 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0007 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0007 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0007 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0007 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0007 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0007 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0007 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0007 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0007 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0007 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0007 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0007 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0007 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0007 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0007 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0007 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0007 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0007 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0007 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0007 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0007 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0007 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0007 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0007 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0007 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0007 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0007 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0007 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0007 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0007 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0007 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0007 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0007 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0007 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0007 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0007 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0007 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0007 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0007 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0007 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0007 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0007 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0007 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0007 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0007 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0007 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0007 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0007 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0007 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0007 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0007 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0007 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0007 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0007 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0007 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0007 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0007 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0007 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0007 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0007 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0007 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0007 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0007 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0007 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0007 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0007 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0007 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0007 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0007 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0007 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0007 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0007 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0007 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0007 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0007 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0007 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0007 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0007 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0007 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0007 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0007 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0007 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0007 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0007 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0007 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0007 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0007 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0007 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0007 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0007 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0007 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0007 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0007 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0007 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0007 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0007 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0007 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0007 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0007 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0007 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0007 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0007 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0007 7.9633e-08 0)
L_S0_01|1 S0_0 _S0_01|A1  2.067833848e-12
L_S0_01|2 _S0_01|A1 _S0_01|A2  4.135667696e-12
L_S0_01|3 _S0_01|A3 _S0_01|A4  8.271335392e-12
L_S0_01|T T10 _S0_01|T1  2.067833848e-12
L_S0_01|4 _S0_01|T1 _S0_01|T2  4.135667696e-12
L_S0_01|5 _S0_01|A4 _S0_01|Q1  4.135667696e-12
L_S0_01|6 _S0_01|Q1 S0_1_TX  2.067833848e-12
IT11|T 0 T10  PWL(0 0 2.7e-11 0 3e-11 0.0007 3.3e-11 0 2.27e-10 0 2.3e-10 0.0007 2.33e-10 0 4.27e-10 0 4.3e-10 0.0007 4.33e-10 0 6.27e-10 0 6.3e-10 0.0007 6.33e-10 0 8.27e-10 0 8.3e-10 0.0007 8.33e-10 0 1.027e-09 0 1.03e-09 0.0007 1.033e-09 0 1.227e-09 0 1.23e-09 0.0007 1.233e-09 0 1.427e-09 0 1.43e-09 0.0007 1.433e-09 0 1.627e-09 0 1.63e-09 0.0007 1.633e-09 0 1.827e-09 0 1.83e-09 0.0007 1.833e-09 0 2.027e-09 0 2.03e-09 0.0007 2.033e-09 0 2.227e-09 0 2.23e-09 0.0007 2.233e-09 0 2.427e-09 0 2.43e-09 0.0007 2.433e-09 0 2.627e-09 0 2.63e-09 0.0007 2.633e-09 0 2.827e-09 0 2.83e-09 0.0007 2.833e-09 0 3.027e-09 0 3.03e-09 0.0007 3.033e-09 0 3.227e-09 0 3.23e-09 0.0007 3.233e-09 0 3.427e-09 0 3.43e-09 0.0007 3.433e-09 0 3.627e-09 0 3.63e-09 0.0007 3.633e-09 0 3.827e-09 0 3.83e-09 0.0007 3.833e-09 0 4.027e-09 0 4.03e-09 0.0007 4.033e-09 0 4.227e-09 0 4.23e-09 0.0007 4.233e-09 0 4.427e-09 0 4.43e-09 0.0007 4.433e-09 0 4.627e-09 0 4.63e-09 0.0007 4.633e-09 0 4.827e-09 0 4.83e-09 0.0007 4.833e-09 0 5.027e-09 0 5.03e-09 0.0007 5.033e-09 0 5.227e-09 0 5.23e-09 0.0007 5.233e-09 0 5.427e-09 0 5.43e-09 0.0007 5.433e-09 0 5.627e-09 0 5.63e-09 0.0007 5.633e-09 0 5.827e-09 0 5.83e-09 0.0007 5.833e-09 0 6.027e-09 0 6.03e-09 0.0007 6.033e-09 0 6.227e-09 0 6.23e-09 0.0007 6.233e-09 0 6.427e-09 0 6.43e-09 0.0007 6.433e-09 0 6.627e-09 0 6.63e-09 0.0007 6.633e-09 0 6.827e-09 0 6.83e-09 0.0007 6.833e-09 0 7.027e-09 0 7.03e-09 0.0007 7.033e-09 0 7.227e-09 0 7.23e-09 0.0007 7.233e-09 0 7.427e-09 0 7.43e-09 0.0007 7.433e-09 0 7.627e-09 0 7.63e-09 0.0007 7.633e-09 0 7.827e-09 0 7.83e-09 0.0007 7.833e-09 0 8.027e-09 0 8.03e-09 0.0007 8.033e-09 0 8.227e-09 0 8.23e-09 0.0007 8.233e-09 0 8.427e-09 0 8.43e-09 0.0007 8.433e-09 0 8.627e-09 0 8.63e-09 0.0007 8.633e-09 0 8.827e-09 0 8.83e-09 0.0007 8.833e-09 0 9.027e-09 0 9.03e-09 0.0007 9.033e-09 0 9.227e-09 0 9.23e-09 0.0007 9.233e-09 0 9.427e-09 0 9.43e-09 0.0007 9.433e-09 0 9.627e-09 0 9.63e-09 0.0007 9.633e-09 0 9.827e-09 0 9.83e-09 0.0007 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0007 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0007 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0007 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0007 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0007 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0007 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0007 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0007 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0007 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0007 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0007 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0007 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0007 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0007 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0007 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0007 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0007 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0007 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0007 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0007 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0007 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0007 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0007 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0007 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0007 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0007 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0007 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0007 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0007 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0007 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0007 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0007 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0007 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0007 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0007 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0007 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0007 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0007 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0007 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0007 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0007 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0007 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0007 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0007 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0007 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0007 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0007 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0007 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0007 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0007 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0007 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0007 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0007 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0007 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0007 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0007 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0007 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0007 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0007 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0007 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0007 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0007 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0007 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0007 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0007 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0007 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0007 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0007 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0007 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0007 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0007 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0007 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0007 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0007 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0007 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0007 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0007 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0007 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0007 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0007 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0007 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0007 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0007 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0007 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0007 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0007 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0007 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0007 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0007 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0007 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0007 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0007 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0007 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0007 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0007 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0007 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0007 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0007 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0007 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0007 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0007 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0007 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0007 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0007 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0007 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0007 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0007 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0007 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0007 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0007 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0007 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0007 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0007 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0007 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0007 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0007 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0007 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0007 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0007 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0007 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0007 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0007 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0007 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0007 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0007 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0007 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0007 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0007 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0007 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0007 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0007 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0007 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0007 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0007 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0007 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0007 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0007 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0007 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0007 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0007 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0007 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0007 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0007 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0007 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0007 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0007 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0007 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0007 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0007 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0007 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0007 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0007 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0007 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0007 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0007 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0007 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0007 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0007 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0007 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0007 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0007 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0007 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0007 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0007 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0007 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0007 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0007 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0007 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0007 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0007 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0007 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0007 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0007 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0007 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0007 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0007 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0007 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0007 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0007 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0007 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0007 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0007 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0007 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0007 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0007 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0007 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0007 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0007 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0007 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0007 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0007 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0007 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0007 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0007 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0007 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0007 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0007 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0007 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0007 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0007 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0007 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0007 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0007 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0007 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0007 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0007 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0007 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0007 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0007 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0007 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0007 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0007 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0007 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0007 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0007 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0007 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0007 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0007 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0007 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0007 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0007 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0007 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0007 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0007 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0007 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0007 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0007 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0007 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0007 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0007 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0007 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0007 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0007 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0007 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0007 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0007 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0007 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0007 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0007 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0007 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0007 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0007 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0007 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0007 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0007 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0007 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0007 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0007 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0007 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0007 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0007 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0007 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0007 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0007 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0007 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0007 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0007 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0007 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0007 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0007 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0007 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0007 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0007 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0007 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0007 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0007 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0007 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0007 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0007 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0007 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0007 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0007 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0007 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0007 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0007 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0007 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0007 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0007 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0007 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0007 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0007 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0007 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0007 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0007 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0007 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0007 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0007 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0007 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0007 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0007 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0007 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0007 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0007 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0007 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0007 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0007 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0007 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0007 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0007 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0007 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0007 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0007 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0007 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0007 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0007 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0007 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0007 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0007 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0007 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0007 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0007 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0007 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0007 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0007 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0007 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0007 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0007 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0007 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0007 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0007 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0007 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0007 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0007 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0007 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0007 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0007 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0007 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0007 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0007 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0007 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0007 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0007 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0007 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0007 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0007 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0007 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0007 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0007 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0007 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0007 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0007 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0007 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0007 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0007 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0007 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0007 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0007 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0007 7.9633e-08 0)
L_S1_01|A1 IG0_0_TO0 _S1_01|A1  2.067833848e-12
L_S1_01|A2 _S1_01|A1 _S1_01|A2  4.135667696e-12
L_S1_01|A3 _S1_01|A3 _S1_01|AB  8.271335392e-12
L_S1_01|B1 IP1_0_OUT _S1_01|B1  2.067833848e-12
L_S1_01|B2 _S1_01|B1 _S1_01|B2  4.135667696e-12
L_S1_01|B3 _S1_01|B3 _S1_01|AB  8.271335392e-12
L_S1_01|T1 T11 _S1_01|T1  2.067833848e-12
L_S1_01|T2 _S1_01|T1 _S1_01|T2  4.135667696e-12
L_S1_01|Q2 _S1_01|ABTQ _S1_01|Q1  4.135667696e-12
L_S1_01|Q1 _S1_01|Q1 S1_1_TX  2.067833848e-12
IT12|T 0 T12  PWL(0 0 2.7e-11 0 3e-11 0.0028 3.3e-11 0 2.27e-10 0 2.3e-10 0.0028 2.33e-10 0 4.27e-10 0 4.3e-10 0.0028 4.33e-10 0 6.27e-10 0 6.3e-10 0.0028 6.33e-10 0 8.27e-10 0 8.3e-10 0.0028 8.33e-10 0 1.027e-09 0 1.03e-09 0.0028 1.033e-09 0 1.227e-09 0 1.23e-09 0.0028 1.233e-09 0 1.427e-09 0 1.43e-09 0.0028 1.433e-09 0 1.627e-09 0 1.63e-09 0.0028 1.633e-09 0 1.827e-09 0 1.83e-09 0.0028 1.833e-09 0 2.027e-09 0 2.03e-09 0.0028 2.033e-09 0 2.227e-09 0 2.23e-09 0.0028 2.233e-09 0 2.427e-09 0 2.43e-09 0.0028 2.433e-09 0 2.627e-09 0 2.63e-09 0.0028 2.633e-09 0 2.827e-09 0 2.83e-09 0.0028 2.833e-09 0 3.027e-09 0 3.03e-09 0.0028 3.033e-09 0 3.227e-09 0 3.23e-09 0.0028 3.233e-09 0 3.427e-09 0 3.43e-09 0.0028 3.433e-09 0 3.627e-09 0 3.63e-09 0.0028 3.633e-09 0 3.827e-09 0 3.83e-09 0.0028 3.833e-09 0 4.027e-09 0 4.03e-09 0.0028 4.033e-09 0 4.227e-09 0 4.23e-09 0.0028 4.233e-09 0 4.427e-09 0 4.43e-09 0.0028 4.433e-09 0 4.627e-09 0 4.63e-09 0.0028 4.633e-09 0 4.827e-09 0 4.83e-09 0.0028 4.833e-09 0 5.027e-09 0 5.03e-09 0.0028 5.033e-09 0 5.227e-09 0 5.23e-09 0.0028 5.233e-09 0 5.427e-09 0 5.43e-09 0.0028 5.433e-09 0 5.627e-09 0 5.63e-09 0.0028 5.633e-09 0 5.827e-09 0 5.83e-09 0.0028 5.833e-09 0 6.027e-09 0 6.03e-09 0.0028 6.033e-09 0 6.227e-09 0 6.23e-09 0.0028 6.233e-09 0 6.427e-09 0 6.43e-09 0.0028 6.433e-09 0 6.627e-09 0 6.63e-09 0.0028 6.633e-09 0 6.827e-09 0 6.83e-09 0.0028 6.833e-09 0 7.027e-09 0 7.03e-09 0.0028 7.033e-09 0 7.227e-09 0 7.23e-09 0.0028 7.233e-09 0 7.427e-09 0 7.43e-09 0.0028 7.433e-09 0 7.627e-09 0 7.63e-09 0.0028 7.633e-09 0 7.827e-09 0 7.83e-09 0.0028 7.833e-09 0 8.027e-09 0 8.03e-09 0.0028 8.033e-09 0 8.227e-09 0 8.23e-09 0.0028 8.233e-09 0 8.427e-09 0 8.43e-09 0.0028 8.433e-09 0 8.627e-09 0 8.63e-09 0.0028 8.633e-09 0 8.827e-09 0 8.83e-09 0.0028 8.833e-09 0 9.027e-09 0 9.03e-09 0.0028 9.033e-09 0 9.227e-09 0 9.23e-09 0.0028 9.233e-09 0 9.427e-09 0 9.43e-09 0.0028 9.433e-09 0 9.627e-09 0 9.63e-09 0.0028 9.633e-09 0 9.827e-09 0 9.83e-09 0.0028 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0028 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0028 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0028 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0028 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0028 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0028 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0028 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0028 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0028 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0028 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0028 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0028 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0028 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0028 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0028 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0028 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0028 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0028 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0028 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0028 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0028 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0028 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0028 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0028 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0028 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0028 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0028 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0028 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0028 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0028 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0028 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0028 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0028 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0028 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0028 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0028 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0028 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0028 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0028 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0028 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0028 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0028 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0028 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0028 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0028 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0028 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0028 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0028 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0028 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0028 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0028 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0028 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0028 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0028 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0028 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0028 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0028 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0028 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0028 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0028 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0028 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0028 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0028 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0028 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0028 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0028 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0028 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0028 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0028 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0028 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0028 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0028 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0028 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0028 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0028 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0028 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0028 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0028 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0028 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0028 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0028 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0028 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0028 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0028 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0028 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0028 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0028 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0028 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0028 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0028 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0028 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0028 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0028 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0028 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0028 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0028 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0028 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0028 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0028 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0028 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0028 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0028 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0028 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0028 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0028 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0028 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0028 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0028 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0028 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0028 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0028 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0028 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0028 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0028 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0028 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0028 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0028 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0028 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0028 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0028 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0028 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0028 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0028 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0028 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0028 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0028 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0028 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0028 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0028 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0028 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0028 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0028 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0028 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0028 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0028 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0028 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0028 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0028 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0028 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0028 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0028 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0028 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0028 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0028 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0028 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0028 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0028 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0028 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0028 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0028 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0028 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0028 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0028 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0028 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0028 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0028 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0028 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0028 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0028 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0028 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0028 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0028 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0028 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0028 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0028 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0028 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0028 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0028 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0028 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0028 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0028 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0028 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0028 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0028 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0028 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0028 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0028 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0028 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0028 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0028 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0028 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0028 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0028 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0028 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0028 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0028 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0028 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0028 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0028 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0028 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0028 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0028 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0028 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0028 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0028 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0028 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0028 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0028 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0028 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0028 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0028 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0028 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0028 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0028 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0028 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0028 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0028 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0028 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0028 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0028 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0028 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0028 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0028 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0028 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0028 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0028 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0028 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0028 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0028 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0028 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0028 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0028 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0028 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0028 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0028 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0028 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0028 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0028 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0028 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0028 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0028 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0028 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0028 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0028 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0028 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0028 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0028 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0028 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0028 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0028 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0028 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0028 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0028 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0028 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0028 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0028 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0028 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0028 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0028 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0028 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0028 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0028 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0028 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0028 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0028 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0028 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0028 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0028 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0028 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0028 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0028 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0028 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0028 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0028 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0028 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0028 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0028 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0028 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0028 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0028 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0028 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0028 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0028 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0028 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0028 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0028 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0028 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0028 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0028 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0028 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0028 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0028 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0028 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0028 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0028 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0028 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0028 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0028 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0028 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0028 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0028 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0028 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0028 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0028 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0028 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0028 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0028 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0028 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0028 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0028 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0028 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0028 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0028 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0028 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0028 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0028 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0028 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0028 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0028 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0028 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0028 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0028 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0028 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0028 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0028 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0028 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0028 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0028 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0028 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0028 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0028 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0028 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0028 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0028 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0028 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0028 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0028 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0028 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0028 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0028 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0028 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0028 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0028 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0028 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0028 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0028 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0028 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0028 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0028 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0028 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0028 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0028 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0028 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0028 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0028 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0028 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0028 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0028 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0028 7.9633e-08 0)
IT13|T 0 T13  PWL(0 0 2.7e-11 0 3e-11 0.0014 3.3e-11 0 2.27e-10 0 2.3e-10 0.0014 2.33e-10 0 4.27e-10 0 4.3e-10 0.0014 4.33e-10 0 6.27e-10 0 6.3e-10 0.0014 6.33e-10 0 8.27e-10 0 8.3e-10 0.0014 8.33e-10 0 1.027e-09 0 1.03e-09 0.0014 1.033e-09 0 1.227e-09 0 1.23e-09 0.0014 1.233e-09 0 1.427e-09 0 1.43e-09 0.0014 1.433e-09 0 1.627e-09 0 1.63e-09 0.0014 1.633e-09 0 1.827e-09 0 1.83e-09 0.0014 1.833e-09 0 2.027e-09 0 2.03e-09 0.0014 2.033e-09 0 2.227e-09 0 2.23e-09 0.0014 2.233e-09 0 2.427e-09 0 2.43e-09 0.0014 2.433e-09 0 2.627e-09 0 2.63e-09 0.0014 2.633e-09 0 2.827e-09 0 2.83e-09 0.0014 2.833e-09 0 3.027e-09 0 3.03e-09 0.0014 3.033e-09 0 3.227e-09 0 3.23e-09 0.0014 3.233e-09 0 3.427e-09 0 3.43e-09 0.0014 3.433e-09 0 3.627e-09 0 3.63e-09 0.0014 3.633e-09 0 3.827e-09 0 3.83e-09 0.0014 3.833e-09 0 4.027e-09 0 4.03e-09 0.0014 4.033e-09 0 4.227e-09 0 4.23e-09 0.0014 4.233e-09 0 4.427e-09 0 4.43e-09 0.0014 4.433e-09 0 4.627e-09 0 4.63e-09 0.0014 4.633e-09 0 4.827e-09 0 4.83e-09 0.0014 4.833e-09 0 5.027e-09 0 5.03e-09 0.0014 5.033e-09 0 5.227e-09 0 5.23e-09 0.0014 5.233e-09 0 5.427e-09 0 5.43e-09 0.0014 5.433e-09 0 5.627e-09 0 5.63e-09 0.0014 5.633e-09 0 5.827e-09 0 5.83e-09 0.0014 5.833e-09 0 6.027e-09 0 6.03e-09 0.0014 6.033e-09 0 6.227e-09 0 6.23e-09 0.0014 6.233e-09 0 6.427e-09 0 6.43e-09 0.0014 6.433e-09 0 6.627e-09 0 6.63e-09 0.0014 6.633e-09 0 6.827e-09 0 6.83e-09 0.0014 6.833e-09 0 7.027e-09 0 7.03e-09 0.0014 7.033e-09 0 7.227e-09 0 7.23e-09 0.0014 7.233e-09 0 7.427e-09 0 7.43e-09 0.0014 7.433e-09 0 7.627e-09 0 7.63e-09 0.0014 7.633e-09 0 7.827e-09 0 7.83e-09 0.0014 7.833e-09 0 8.027e-09 0 8.03e-09 0.0014 8.033e-09 0 8.227e-09 0 8.23e-09 0.0014 8.233e-09 0 8.427e-09 0 8.43e-09 0.0014 8.433e-09 0 8.627e-09 0 8.63e-09 0.0014 8.633e-09 0 8.827e-09 0 8.83e-09 0.0014 8.833e-09 0 9.027e-09 0 9.03e-09 0.0014 9.033e-09 0 9.227e-09 0 9.23e-09 0.0014 9.233e-09 0 9.427e-09 0 9.43e-09 0.0014 9.433e-09 0 9.627e-09 0 9.63e-09 0.0014 9.633e-09 0 9.827e-09 0 9.83e-09 0.0014 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0014 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0014 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0014 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0014 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0014 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0014 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0014 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0014 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0014 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0014 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0014 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0014 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0014 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0014 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0014 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0014 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0014 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0014 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0014 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0014 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0014 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0014 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0014 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0014 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0014 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0014 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0014 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0014 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0014 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0014 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0014 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0014 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0014 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0014 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0014 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0014 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0014 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0014 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0014 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0014 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0014 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0014 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0014 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0014 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0014 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0014 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0014 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0014 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0014 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0014 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0014 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0014 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0014 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0014 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0014 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0014 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0014 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0014 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0014 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0014 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0014 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0014 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0014 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0014 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0014 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0014 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0014 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0014 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0014 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0014 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0014 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0014 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0014 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0014 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0014 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0014 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0014 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0014 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0014 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0014 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0014 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0014 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0014 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0014 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0014 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0014 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0014 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0014 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0014 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0014 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0014 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0014 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0014 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0014 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0014 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0014 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0014 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0014 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0014 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0014 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0014 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0014 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0014 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0014 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0014 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0014 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0014 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0014 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0014 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0014 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0014 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0014 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0014 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0014 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0014 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0014 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0014 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0014 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0014 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0014 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0014 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0014 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0014 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0014 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0014 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0014 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0014 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0014 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0014 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0014 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0014 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0014 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0014 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0014 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0014 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0014 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0014 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0014 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0014 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0014 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0014 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0014 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0014 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0014 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0014 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0014 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0014 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0014 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0014 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0014 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0014 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0014 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0014 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0014 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0014 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0014 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0014 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0014 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0014 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0014 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0014 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0014 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0014 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0014 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0014 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0014 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0014 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0014 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0014 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0014 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0014 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0014 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0014 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0014 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0014 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0014 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0014 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0014 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0014 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0014 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0014 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0014 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0014 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0014 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0014 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0014 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0014 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0014 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0014 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0014 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0014 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0014 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0014 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0014 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0014 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0014 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0014 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0014 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0014 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0014 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0014 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0014 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0014 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0014 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0014 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0014 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0014 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0014 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0014 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0014 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0014 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0014 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0014 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0014 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0014 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0014 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0014 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0014 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0014 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0014 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0014 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0014 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0014 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0014 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0014 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0014 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0014 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0014 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0014 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0014 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0014 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0014 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0014 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0014 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0014 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0014 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0014 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0014 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0014 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0014 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0014 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0014 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0014 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0014 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0014 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0014 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0014 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0014 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0014 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0014 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0014 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0014 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0014 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0014 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0014 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0014 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0014 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0014 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0014 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0014 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0014 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0014 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0014 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0014 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0014 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0014 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0014 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0014 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0014 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0014 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0014 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0014 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0014 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0014 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0014 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0014 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0014 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0014 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0014 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0014 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0014 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0014 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0014 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0014 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0014 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0014 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0014 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0014 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0014 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0014 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0014 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0014 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0014 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0014 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0014 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0014 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0014 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0014 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0014 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0014 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0014 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0014 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0014 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0014 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0014 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0014 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0014 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0014 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0014 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0014 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0014 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0014 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0014 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0014 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0014 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0014 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0014 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0014 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0014 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0014 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0014 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0014 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0014 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0014 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0014 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0014 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0014 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0014 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0014 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0014 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0014 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0014 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0014 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0014 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0014 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0014 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0014 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0014 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0014 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0014 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0014 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0014 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0014 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0014 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0014 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0014 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0014 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0014 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0014 7.9633e-08 0)
IT14|T 0 T14  PWL(0 0 2.7e-11 0 3e-11 0.0028 3.3e-11 0 2.27e-10 0 2.3e-10 0.0028 2.33e-10 0 4.27e-10 0 4.3e-10 0.0028 4.33e-10 0 6.27e-10 0 6.3e-10 0.0028 6.33e-10 0 8.27e-10 0 8.3e-10 0.0028 8.33e-10 0 1.027e-09 0 1.03e-09 0.0028 1.033e-09 0 1.227e-09 0 1.23e-09 0.0028 1.233e-09 0 1.427e-09 0 1.43e-09 0.0028 1.433e-09 0 1.627e-09 0 1.63e-09 0.0028 1.633e-09 0 1.827e-09 0 1.83e-09 0.0028 1.833e-09 0 2.027e-09 0 2.03e-09 0.0028 2.033e-09 0 2.227e-09 0 2.23e-09 0.0028 2.233e-09 0 2.427e-09 0 2.43e-09 0.0028 2.433e-09 0 2.627e-09 0 2.63e-09 0.0028 2.633e-09 0 2.827e-09 0 2.83e-09 0.0028 2.833e-09 0 3.027e-09 0 3.03e-09 0.0028 3.033e-09 0 3.227e-09 0 3.23e-09 0.0028 3.233e-09 0 3.427e-09 0 3.43e-09 0.0028 3.433e-09 0 3.627e-09 0 3.63e-09 0.0028 3.633e-09 0 3.827e-09 0 3.83e-09 0.0028 3.833e-09 0 4.027e-09 0 4.03e-09 0.0028 4.033e-09 0 4.227e-09 0 4.23e-09 0.0028 4.233e-09 0 4.427e-09 0 4.43e-09 0.0028 4.433e-09 0 4.627e-09 0 4.63e-09 0.0028 4.633e-09 0 4.827e-09 0 4.83e-09 0.0028 4.833e-09 0 5.027e-09 0 5.03e-09 0.0028 5.033e-09 0 5.227e-09 0 5.23e-09 0.0028 5.233e-09 0 5.427e-09 0 5.43e-09 0.0028 5.433e-09 0 5.627e-09 0 5.63e-09 0.0028 5.633e-09 0 5.827e-09 0 5.83e-09 0.0028 5.833e-09 0 6.027e-09 0 6.03e-09 0.0028 6.033e-09 0 6.227e-09 0 6.23e-09 0.0028 6.233e-09 0 6.427e-09 0 6.43e-09 0.0028 6.433e-09 0 6.627e-09 0 6.63e-09 0.0028 6.633e-09 0 6.827e-09 0 6.83e-09 0.0028 6.833e-09 0 7.027e-09 0 7.03e-09 0.0028 7.033e-09 0 7.227e-09 0 7.23e-09 0.0028 7.233e-09 0 7.427e-09 0 7.43e-09 0.0028 7.433e-09 0 7.627e-09 0 7.63e-09 0.0028 7.633e-09 0 7.827e-09 0 7.83e-09 0.0028 7.833e-09 0 8.027e-09 0 8.03e-09 0.0028 8.033e-09 0 8.227e-09 0 8.23e-09 0.0028 8.233e-09 0 8.427e-09 0 8.43e-09 0.0028 8.433e-09 0 8.627e-09 0 8.63e-09 0.0028 8.633e-09 0 8.827e-09 0 8.83e-09 0.0028 8.833e-09 0 9.027e-09 0 9.03e-09 0.0028 9.033e-09 0 9.227e-09 0 9.23e-09 0.0028 9.233e-09 0 9.427e-09 0 9.43e-09 0.0028 9.433e-09 0 9.627e-09 0 9.63e-09 0.0028 9.633e-09 0 9.827e-09 0 9.83e-09 0.0028 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0028 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0028 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0028 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0028 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0028 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0028 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0028 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0028 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0028 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0028 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0028 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0028 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0028 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0028 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0028 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0028 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0028 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0028 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0028 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0028 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0028 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0028 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0028 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0028 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0028 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0028 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0028 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0028 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0028 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0028 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0028 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0028 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0028 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0028 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0028 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0028 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0028 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0028 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0028 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0028 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0028 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0028 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0028 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0028 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0028 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0028 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0028 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0028 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0028 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0028 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0028 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0028 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0028 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0028 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0028 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0028 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0028 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0028 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0028 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0028 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0028 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0028 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0028 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0028 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0028 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0028 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0028 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0028 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0028 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0028 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0028 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0028 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0028 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0028 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0028 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0028 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0028 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0028 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0028 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0028 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0028 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0028 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0028 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0028 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0028 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0028 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0028 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0028 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0028 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0028 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0028 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0028 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0028 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0028 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0028 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0028 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0028 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0028 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0028 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0028 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0028 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0028 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0028 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0028 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0028 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0028 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0028 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0028 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0028 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0028 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0028 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0028 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0028 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0028 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0028 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0028 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0028 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0028 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0028 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0028 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0028 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0028 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0028 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0028 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0028 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0028 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0028 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0028 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0028 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0028 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0028 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0028 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0028 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0028 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0028 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0028 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0028 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0028 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0028 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0028 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0028 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0028 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0028 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0028 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0028 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0028 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0028 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0028 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0028 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0028 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0028 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0028 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0028 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0028 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0028 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0028 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0028 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0028 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0028 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0028 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0028 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0028 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0028 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0028 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0028 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0028 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0028 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0028 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0028 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0028 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0028 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0028 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0028 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0028 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0028 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0028 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0028 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0028 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0028 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0028 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0028 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0028 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0028 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0028 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0028 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0028 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0028 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0028 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0028 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0028 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0028 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0028 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0028 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0028 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0028 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0028 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0028 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0028 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0028 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0028 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0028 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0028 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0028 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0028 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0028 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0028 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0028 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0028 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0028 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0028 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0028 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0028 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0028 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0028 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0028 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0028 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0028 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0028 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0028 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0028 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0028 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0028 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0028 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0028 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0028 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0028 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0028 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0028 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0028 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0028 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0028 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0028 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0028 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0028 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0028 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0028 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0028 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0028 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0028 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0028 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0028 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0028 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0028 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0028 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0028 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0028 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0028 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0028 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0028 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0028 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0028 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0028 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0028 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0028 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0028 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0028 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0028 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0028 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0028 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0028 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0028 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0028 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0028 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0028 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0028 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0028 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0028 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0028 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0028 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0028 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0028 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0028 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0028 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0028 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0028 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0028 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0028 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0028 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0028 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0028 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0028 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0028 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0028 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0028 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0028 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0028 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0028 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0028 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0028 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0028 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0028 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0028 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0028 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0028 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0028 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0028 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0028 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0028 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0028 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0028 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0028 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0028 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0028 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0028 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0028 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0028 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0028 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0028 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0028 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0028 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0028 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0028 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0028 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0028 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0028 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0028 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0028 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0028 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0028 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0028 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0028 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0028 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0028 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0028 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0028 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0028 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0028 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0028 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0028 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0028 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0028 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0028 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0028 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0028 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0028 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0028 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0028 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0028 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0028 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0028 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0028 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0028 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0028 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0028 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0028 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0028 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0028 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0028 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0028 7.9633e-08 0)
IT15|T 0 T15  PWL(0 0 2.7e-11 0 3e-11 0.0007 3.3e-11 0 2.27e-10 0 2.3e-10 0.0007 2.33e-10 0 4.27e-10 0 4.3e-10 0.0007 4.33e-10 0 6.27e-10 0 6.3e-10 0.0007 6.33e-10 0 8.27e-10 0 8.3e-10 0.0007 8.33e-10 0 1.027e-09 0 1.03e-09 0.0007 1.033e-09 0 1.227e-09 0 1.23e-09 0.0007 1.233e-09 0 1.427e-09 0 1.43e-09 0.0007 1.433e-09 0 1.627e-09 0 1.63e-09 0.0007 1.633e-09 0 1.827e-09 0 1.83e-09 0.0007 1.833e-09 0 2.027e-09 0 2.03e-09 0.0007 2.033e-09 0 2.227e-09 0 2.23e-09 0.0007 2.233e-09 0 2.427e-09 0 2.43e-09 0.0007 2.433e-09 0 2.627e-09 0 2.63e-09 0.0007 2.633e-09 0 2.827e-09 0 2.83e-09 0.0007 2.833e-09 0 3.027e-09 0 3.03e-09 0.0007 3.033e-09 0 3.227e-09 0 3.23e-09 0.0007 3.233e-09 0 3.427e-09 0 3.43e-09 0.0007 3.433e-09 0 3.627e-09 0 3.63e-09 0.0007 3.633e-09 0 3.827e-09 0 3.83e-09 0.0007 3.833e-09 0 4.027e-09 0 4.03e-09 0.0007 4.033e-09 0 4.227e-09 0 4.23e-09 0.0007 4.233e-09 0 4.427e-09 0 4.43e-09 0.0007 4.433e-09 0 4.627e-09 0 4.63e-09 0.0007 4.633e-09 0 4.827e-09 0 4.83e-09 0.0007 4.833e-09 0 5.027e-09 0 5.03e-09 0.0007 5.033e-09 0 5.227e-09 0 5.23e-09 0.0007 5.233e-09 0 5.427e-09 0 5.43e-09 0.0007 5.433e-09 0 5.627e-09 0 5.63e-09 0.0007 5.633e-09 0 5.827e-09 0 5.83e-09 0.0007 5.833e-09 0 6.027e-09 0 6.03e-09 0.0007 6.033e-09 0 6.227e-09 0 6.23e-09 0.0007 6.233e-09 0 6.427e-09 0 6.43e-09 0.0007 6.433e-09 0 6.627e-09 0 6.63e-09 0.0007 6.633e-09 0 6.827e-09 0 6.83e-09 0.0007 6.833e-09 0 7.027e-09 0 7.03e-09 0.0007 7.033e-09 0 7.227e-09 0 7.23e-09 0.0007 7.233e-09 0 7.427e-09 0 7.43e-09 0.0007 7.433e-09 0 7.627e-09 0 7.63e-09 0.0007 7.633e-09 0 7.827e-09 0 7.83e-09 0.0007 7.833e-09 0 8.027e-09 0 8.03e-09 0.0007 8.033e-09 0 8.227e-09 0 8.23e-09 0.0007 8.233e-09 0 8.427e-09 0 8.43e-09 0.0007 8.433e-09 0 8.627e-09 0 8.63e-09 0.0007 8.633e-09 0 8.827e-09 0 8.83e-09 0.0007 8.833e-09 0 9.027e-09 0 9.03e-09 0.0007 9.033e-09 0 9.227e-09 0 9.23e-09 0.0007 9.233e-09 0 9.427e-09 0 9.43e-09 0.0007 9.433e-09 0 9.627e-09 0 9.63e-09 0.0007 9.633e-09 0 9.827e-09 0 9.83e-09 0.0007 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0007 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0007 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0007 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0007 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0007 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0007 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0007 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0007 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0007 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0007 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0007 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0007 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0007 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0007 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0007 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0007 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0007 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0007 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0007 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0007 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0007 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0007 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0007 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0007 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0007 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0007 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0007 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0007 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0007 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0007 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0007 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0007 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0007 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0007 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0007 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0007 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0007 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0007 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0007 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0007 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0007 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0007 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0007 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0007 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0007 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0007 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0007 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0007 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0007 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0007 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0007 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0007 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0007 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0007 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0007 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0007 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0007 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0007 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0007 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0007 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0007 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0007 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0007 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0007 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0007 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0007 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0007 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0007 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0007 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0007 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0007 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0007 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0007 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0007 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0007 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0007 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0007 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0007 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0007 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0007 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0007 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0007 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0007 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0007 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0007 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0007 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0007 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0007 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0007 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0007 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0007 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0007 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0007 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0007 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0007 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0007 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0007 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0007 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0007 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0007 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0007 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0007 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0007 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0007 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0007 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0007 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0007 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0007 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0007 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0007 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0007 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0007 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0007 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0007 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0007 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0007 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0007 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0007 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0007 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0007 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0007 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0007 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0007 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0007 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0007 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0007 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0007 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0007 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0007 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0007 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0007 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0007 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0007 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0007 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0007 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0007 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0007 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0007 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0007 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0007 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0007 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0007 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0007 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0007 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0007 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0007 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0007 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0007 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0007 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0007 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0007 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0007 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0007 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0007 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0007 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0007 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0007 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0007 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0007 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0007 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0007 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0007 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0007 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0007 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0007 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0007 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0007 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0007 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0007 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0007 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0007 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0007 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0007 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0007 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0007 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0007 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0007 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0007 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0007 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0007 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0007 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0007 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0007 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0007 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0007 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0007 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0007 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0007 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0007 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0007 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0007 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0007 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0007 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0007 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0007 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0007 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0007 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0007 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0007 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0007 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0007 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0007 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0007 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0007 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0007 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0007 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0007 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0007 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0007 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0007 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0007 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0007 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0007 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0007 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0007 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0007 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0007 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0007 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0007 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0007 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0007 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0007 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0007 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0007 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0007 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0007 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0007 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0007 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0007 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0007 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0007 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0007 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0007 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0007 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0007 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0007 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0007 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0007 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0007 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0007 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0007 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0007 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0007 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0007 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0007 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0007 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0007 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0007 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0007 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0007 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0007 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0007 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0007 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0007 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0007 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0007 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0007 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0007 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0007 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0007 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0007 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0007 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0007 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0007 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0007 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0007 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0007 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0007 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0007 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0007 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0007 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0007 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0007 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0007 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0007 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0007 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0007 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0007 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0007 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0007 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0007 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0007 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0007 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0007 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0007 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0007 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0007 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0007 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0007 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0007 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0007 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0007 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0007 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0007 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0007 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0007 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0007 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0007 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0007 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0007 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0007 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0007 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0007 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0007 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0007 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0007 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0007 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0007 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0007 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0007 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0007 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0007 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0007 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0007 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0007 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0007 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0007 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0007 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0007 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0007 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0007 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0007 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0007 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0007 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0007 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0007 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0007 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0007 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0007 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0007 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0007 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0007 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0007 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0007 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0007 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0007 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0007 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0007 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0007 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0007 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0007 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0007 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0007 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0007 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0007 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0007 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0007 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0007 7.9633e-08 0)
L_IP3_OUT|1 IP3_0_OUT _IP3_OUT|A1  2.067833848e-12
L_IP3_OUT|2 _IP3_OUT|A1 _IP3_OUT|A2  4.135667696e-12
L_IP3_OUT|3 _IP3_OUT|A3 _IP3_OUT|A4  8.271335392e-12
L_IP3_OUT|T T15 _IP3_OUT|T1  2.067833848e-12
L_IP3_OUT|4 _IP3_OUT|T1 _IP3_OUT|T2  4.135667696e-12
L_IP3_OUT|5 _IP3_OUT|A4 _IP3_OUT|Q1  4.135667696e-12
L_IP3_OUT|6 _IP3_OUT|Q1 IP3_1_OUT_TX  2.067833848e-12
IT16|T 0 T16  PWL(0 0 2.7e-11 0 3e-11 0.0014 3.3e-11 0 2.27e-10 0 2.3e-10 0.0014 2.33e-10 0 4.27e-10 0 4.3e-10 0.0014 4.33e-10 0 6.27e-10 0 6.3e-10 0.0014 6.33e-10 0 8.27e-10 0 8.3e-10 0.0014 8.33e-10 0 1.027e-09 0 1.03e-09 0.0014 1.033e-09 0 1.227e-09 0 1.23e-09 0.0014 1.233e-09 0 1.427e-09 0 1.43e-09 0.0014 1.433e-09 0 1.627e-09 0 1.63e-09 0.0014 1.633e-09 0 1.827e-09 0 1.83e-09 0.0014 1.833e-09 0 2.027e-09 0 2.03e-09 0.0014 2.033e-09 0 2.227e-09 0 2.23e-09 0.0014 2.233e-09 0 2.427e-09 0 2.43e-09 0.0014 2.433e-09 0 2.627e-09 0 2.63e-09 0.0014 2.633e-09 0 2.827e-09 0 2.83e-09 0.0014 2.833e-09 0 3.027e-09 0 3.03e-09 0.0014 3.033e-09 0 3.227e-09 0 3.23e-09 0.0014 3.233e-09 0 3.427e-09 0 3.43e-09 0.0014 3.433e-09 0 3.627e-09 0 3.63e-09 0.0014 3.633e-09 0 3.827e-09 0 3.83e-09 0.0014 3.833e-09 0 4.027e-09 0 4.03e-09 0.0014 4.033e-09 0 4.227e-09 0 4.23e-09 0.0014 4.233e-09 0 4.427e-09 0 4.43e-09 0.0014 4.433e-09 0 4.627e-09 0 4.63e-09 0.0014 4.633e-09 0 4.827e-09 0 4.83e-09 0.0014 4.833e-09 0 5.027e-09 0 5.03e-09 0.0014 5.033e-09 0 5.227e-09 0 5.23e-09 0.0014 5.233e-09 0 5.427e-09 0 5.43e-09 0.0014 5.433e-09 0 5.627e-09 0 5.63e-09 0.0014 5.633e-09 0 5.827e-09 0 5.83e-09 0.0014 5.833e-09 0 6.027e-09 0 6.03e-09 0.0014 6.033e-09 0 6.227e-09 0 6.23e-09 0.0014 6.233e-09 0 6.427e-09 0 6.43e-09 0.0014 6.433e-09 0 6.627e-09 0 6.63e-09 0.0014 6.633e-09 0 6.827e-09 0 6.83e-09 0.0014 6.833e-09 0 7.027e-09 0 7.03e-09 0.0014 7.033e-09 0 7.227e-09 0 7.23e-09 0.0014 7.233e-09 0 7.427e-09 0 7.43e-09 0.0014 7.433e-09 0 7.627e-09 0 7.63e-09 0.0014 7.633e-09 0 7.827e-09 0 7.83e-09 0.0014 7.833e-09 0 8.027e-09 0 8.03e-09 0.0014 8.033e-09 0 8.227e-09 0 8.23e-09 0.0014 8.233e-09 0 8.427e-09 0 8.43e-09 0.0014 8.433e-09 0 8.627e-09 0 8.63e-09 0.0014 8.633e-09 0 8.827e-09 0 8.83e-09 0.0014 8.833e-09 0 9.027e-09 0 9.03e-09 0.0014 9.033e-09 0 9.227e-09 0 9.23e-09 0.0014 9.233e-09 0 9.427e-09 0 9.43e-09 0.0014 9.433e-09 0 9.627e-09 0 9.63e-09 0.0014 9.633e-09 0 9.827e-09 0 9.83e-09 0.0014 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0014 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0014 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0014 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0014 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0014 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0014 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0014 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0014 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0014 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0014 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0014 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0014 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0014 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0014 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0014 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0014 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0014 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0014 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0014 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0014 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0014 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0014 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0014 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0014 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0014 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0014 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0014 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0014 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0014 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0014 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0014 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0014 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0014 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0014 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0014 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0014 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0014 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0014 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0014 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0014 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0014 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0014 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0014 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0014 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0014 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0014 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0014 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0014 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0014 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0014 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0014 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0014 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0014 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0014 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0014 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0014 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0014 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0014 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0014 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0014 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0014 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0014 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0014 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0014 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0014 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0014 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0014 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0014 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0014 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0014 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0014 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0014 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0014 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0014 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0014 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0014 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0014 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0014 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0014 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0014 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0014 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0014 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0014 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0014 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0014 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0014 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0014 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0014 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0014 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0014 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0014 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0014 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0014 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0014 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0014 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0014 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0014 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0014 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0014 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0014 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0014 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0014 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0014 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0014 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0014 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0014 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0014 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0014 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0014 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0014 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0014 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0014 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0014 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0014 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0014 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0014 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0014 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0014 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0014 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0014 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0014 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0014 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0014 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0014 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0014 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0014 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0014 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0014 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0014 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0014 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0014 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0014 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0014 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0014 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0014 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0014 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0014 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0014 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0014 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0014 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0014 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0014 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0014 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0014 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0014 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0014 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0014 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0014 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0014 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0014 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0014 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0014 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0014 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0014 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0014 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0014 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0014 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0014 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0014 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0014 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0014 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0014 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0014 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0014 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0014 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0014 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0014 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0014 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0014 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0014 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0014 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0014 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0014 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0014 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0014 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0014 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0014 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0014 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0014 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0014 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0014 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0014 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0014 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0014 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0014 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0014 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0014 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0014 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0014 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0014 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0014 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0014 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0014 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0014 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0014 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0014 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0014 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0014 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0014 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0014 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0014 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0014 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0014 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0014 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0014 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0014 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0014 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0014 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0014 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0014 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0014 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0014 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0014 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0014 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0014 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0014 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0014 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0014 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0014 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0014 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0014 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0014 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0014 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0014 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0014 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0014 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0014 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0014 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0014 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0014 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0014 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0014 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0014 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0014 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0014 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0014 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0014 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0014 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0014 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0014 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0014 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0014 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0014 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0014 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0014 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0014 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0014 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0014 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0014 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0014 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0014 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0014 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0014 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0014 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0014 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0014 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0014 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0014 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0014 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0014 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0014 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0014 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0014 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0014 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0014 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0014 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0014 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0014 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0014 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0014 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0014 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0014 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0014 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0014 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0014 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0014 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0014 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0014 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0014 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0014 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0014 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0014 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0014 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0014 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0014 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0014 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0014 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0014 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0014 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0014 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0014 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0014 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0014 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0014 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0014 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0014 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0014 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0014 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0014 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0014 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0014 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0014 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0014 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0014 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0014 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0014 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0014 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0014 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0014 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0014 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0014 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0014 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0014 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0014 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0014 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0014 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0014 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0014 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0014 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0014 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0014 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0014 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0014 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0014 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0014 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0014 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0014 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0014 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0014 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0014 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0014 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0014 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0014 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0014 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0014 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0014 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0014 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0014 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0014 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0014 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0014 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0014 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0014 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0014 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0014 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0014 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0014 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0014 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0014 7.9633e-08 0)
IT17|T 0 T17  PWL(0 0 2.7e-11 0 3e-11 0.0028 3.3e-11 0 2.27e-10 0 2.3e-10 0.0028 2.33e-10 0 4.27e-10 0 4.3e-10 0.0028 4.33e-10 0 6.27e-10 0 6.3e-10 0.0028 6.33e-10 0 8.27e-10 0 8.3e-10 0.0028 8.33e-10 0 1.027e-09 0 1.03e-09 0.0028 1.033e-09 0 1.227e-09 0 1.23e-09 0.0028 1.233e-09 0 1.427e-09 0 1.43e-09 0.0028 1.433e-09 0 1.627e-09 0 1.63e-09 0.0028 1.633e-09 0 1.827e-09 0 1.83e-09 0.0028 1.833e-09 0 2.027e-09 0 2.03e-09 0.0028 2.033e-09 0 2.227e-09 0 2.23e-09 0.0028 2.233e-09 0 2.427e-09 0 2.43e-09 0.0028 2.433e-09 0 2.627e-09 0 2.63e-09 0.0028 2.633e-09 0 2.827e-09 0 2.83e-09 0.0028 2.833e-09 0 3.027e-09 0 3.03e-09 0.0028 3.033e-09 0 3.227e-09 0 3.23e-09 0.0028 3.233e-09 0 3.427e-09 0 3.43e-09 0.0028 3.433e-09 0 3.627e-09 0 3.63e-09 0.0028 3.633e-09 0 3.827e-09 0 3.83e-09 0.0028 3.833e-09 0 4.027e-09 0 4.03e-09 0.0028 4.033e-09 0 4.227e-09 0 4.23e-09 0.0028 4.233e-09 0 4.427e-09 0 4.43e-09 0.0028 4.433e-09 0 4.627e-09 0 4.63e-09 0.0028 4.633e-09 0 4.827e-09 0 4.83e-09 0.0028 4.833e-09 0 5.027e-09 0 5.03e-09 0.0028 5.033e-09 0 5.227e-09 0 5.23e-09 0.0028 5.233e-09 0 5.427e-09 0 5.43e-09 0.0028 5.433e-09 0 5.627e-09 0 5.63e-09 0.0028 5.633e-09 0 5.827e-09 0 5.83e-09 0.0028 5.833e-09 0 6.027e-09 0 6.03e-09 0.0028 6.033e-09 0 6.227e-09 0 6.23e-09 0.0028 6.233e-09 0 6.427e-09 0 6.43e-09 0.0028 6.433e-09 0 6.627e-09 0 6.63e-09 0.0028 6.633e-09 0 6.827e-09 0 6.83e-09 0.0028 6.833e-09 0 7.027e-09 0 7.03e-09 0.0028 7.033e-09 0 7.227e-09 0 7.23e-09 0.0028 7.233e-09 0 7.427e-09 0 7.43e-09 0.0028 7.433e-09 0 7.627e-09 0 7.63e-09 0.0028 7.633e-09 0 7.827e-09 0 7.83e-09 0.0028 7.833e-09 0 8.027e-09 0 8.03e-09 0.0028 8.033e-09 0 8.227e-09 0 8.23e-09 0.0028 8.233e-09 0 8.427e-09 0 8.43e-09 0.0028 8.433e-09 0 8.627e-09 0 8.63e-09 0.0028 8.633e-09 0 8.827e-09 0 8.83e-09 0.0028 8.833e-09 0 9.027e-09 0 9.03e-09 0.0028 9.033e-09 0 9.227e-09 0 9.23e-09 0.0028 9.233e-09 0 9.427e-09 0 9.43e-09 0.0028 9.433e-09 0 9.627e-09 0 9.63e-09 0.0028 9.633e-09 0 9.827e-09 0 9.83e-09 0.0028 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0028 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0028 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0028 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0028 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0028 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0028 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0028 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0028 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0028 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0028 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0028 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0028 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0028 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0028 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0028 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0028 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0028 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0028 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0028 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0028 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0028 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0028 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0028 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0028 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0028 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0028 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0028 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0028 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0028 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0028 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0028 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0028 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0028 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0028 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0028 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0028 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0028 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0028 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0028 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0028 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0028 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0028 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0028 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0028 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0028 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0028 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0028 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0028 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0028 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0028 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0028 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0028 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0028 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0028 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0028 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0028 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0028 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0028 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0028 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0028 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0028 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0028 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0028 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0028 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0028 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0028 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0028 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0028 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0028 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0028 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0028 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0028 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0028 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0028 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0028 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0028 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0028 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0028 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0028 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0028 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0028 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0028 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0028 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0028 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0028 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0028 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0028 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0028 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0028 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0028 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0028 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0028 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0028 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0028 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0028 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0028 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0028 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0028 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0028 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0028 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0028 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0028 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0028 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0028 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0028 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0028 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0028 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0028 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0028 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0028 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0028 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0028 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0028 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0028 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0028 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0028 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0028 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0028 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0028 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0028 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0028 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0028 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0028 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0028 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0028 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0028 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0028 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0028 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0028 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0028 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0028 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0028 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0028 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0028 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0028 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0028 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0028 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0028 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0028 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0028 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0028 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0028 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0028 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0028 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0028 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0028 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0028 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0028 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0028 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0028 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0028 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0028 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0028 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0028 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0028 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0028 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0028 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0028 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0028 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0028 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0028 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0028 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0028 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0028 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0028 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0028 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0028 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0028 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0028 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0028 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0028 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0028 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0028 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0028 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0028 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0028 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0028 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0028 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0028 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0028 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0028 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0028 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0028 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0028 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0028 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0028 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0028 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0028 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0028 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0028 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0028 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0028 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0028 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0028 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0028 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0028 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0028 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0028 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0028 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0028 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0028 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0028 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0028 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0028 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0028 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0028 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0028 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0028 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0028 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0028 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0028 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0028 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0028 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0028 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0028 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0028 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0028 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0028 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0028 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0028 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0028 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0028 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0028 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0028 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0028 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0028 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0028 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0028 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0028 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0028 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0028 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0028 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0028 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0028 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0028 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0028 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0028 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0028 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0028 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0028 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0028 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0028 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0028 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0028 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0028 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0028 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0028 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0028 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0028 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0028 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0028 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0028 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0028 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0028 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0028 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0028 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0028 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0028 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0028 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0028 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0028 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0028 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0028 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0028 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0028 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0028 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0028 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0028 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0028 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0028 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0028 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0028 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0028 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0028 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0028 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0028 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0028 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0028 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0028 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0028 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0028 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0028 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0028 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0028 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0028 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0028 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0028 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0028 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0028 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0028 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0028 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0028 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0028 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0028 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0028 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0028 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0028 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0028 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0028 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0028 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0028 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0028 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0028 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0028 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0028 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0028 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0028 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0028 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0028 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0028 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0028 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0028 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0028 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0028 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0028 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0028 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0028 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0028 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0028 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0028 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0028 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0028 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0028 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0028 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0028 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0028 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0028 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0028 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0028 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0028 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0028 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0028 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0028 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0028 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0028 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0028 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0028 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0028 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0028 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0028 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0028 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0028 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0028 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0028 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0028 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0028 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0028 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0028 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0028 7.9633e-08 0)
IT18|T 0 T18  PWL(0 0 2.7e-11 0 3e-11 0.0007 3.3e-11 0 2.27e-10 0 2.3e-10 0.0007 2.33e-10 0 4.27e-10 0 4.3e-10 0.0007 4.33e-10 0 6.27e-10 0 6.3e-10 0.0007 6.33e-10 0 8.27e-10 0 8.3e-10 0.0007 8.33e-10 0 1.027e-09 0 1.03e-09 0.0007 1.033e-09 0 1.227e-09 0 1.23e-09 0.0007 1.233e-09 0 1.427e-09 0 1.43e-09 0.0007 1.433e-09 0 1.627e-09 0 1.63e-09 0.0007 1.633e-09 0 1.827e-09 0 1.83e-09 0.0007 1.833e-09 0 2.027e-09 0 2.03e-09 0.0007 2.033e-09 0 2.227e-09 0 2.23e-09 0.0007 2.233e-09 0 2.427e-09 0 2.43e-09 0.0007 2.433e-09 0 2.627e-09 0 2.63e-09 0.0007 2.633e-09 0 2.827e-09 0 2.83e-09 0.0007 2.833e-09 0 3.027e-09 0 3.03e-09 0.0007 3.033e-09 0 3.227e-09 0 3.23e-09 0.0007 3.233e-09 0 3.427e-09 0 3.43e-09 0.0007 3.433e-09 0 3.627e-09 0 3.63e-09 0.0007 3.633e-09 0 3.827e-09 0 3.83e-09 0.0007 3.833e-09 0 4.027e-09 0 4.03e-09 0.0007 4.033e-09 0 4.227e-09 0 4.23e-09 0.0007 4.233e-09 0 4.427e-09 0 4.43e-09 0.0007 4.433e-09 0 4.627e-09 0 4.63e-09 0.0007 4.633e-09 0 4.827e-09 0 4.83e-09 0.0007 4.833e-09 0 5.027e-09 0 5.03e-09 0.0007 5.033e-09 0 5.227e-09 0 5.23e-09 0.0007 5.233e-09 0 5.427e-09 0 5.43e-09 0.0007 5.433e-09 0 5.627e-09 0 5.63e-09 0.0007 5.633e-09 0 5.827e-09 0 5.83e-09 0.0007 5.833e-09 0 6.027e-09 0 6.03e-09 0.0007 6.033e-09 0 6.227e-09 0 6.23e-09 0.0007 6.233e-09 0 6.427e-09 0 6.43e-09 0.0007 6.433e-09 0 6.627e-09 0 6.63e-09 0.0007 6.633e-09 0 6.827e-09 0 6.83e-09 0.0007 6.833e-09 0 7.027e-09 0 7.03e-09 0.0007 7.033e-09 0 7.227e-09 0 7.23e-09 0.0007 7.233e-09 0 7.427e-09 0 7.43e-09 0.0007 7.433e-09 0 7.627e-09 0 7.63e-09 0.0007 7.633e-09 0 7.827e-09 0 7.83e-09 0.0007 7.833e-09 0 8.027e-09 0 8.03e-09 0.0007 8.033e-09 0 8.227e-09 0 8.23e-09 0.0007 8.233e-09 0 8.427e-09 0 8.43e-09 0.0007 8.433e-09 0 8.627e-09 0 8.63e-09 0.0007 8.633e-09 0 8.827e-09 0 8.83e-09 0.0007 8.833e-09 0 9.027e-09 0 9.03e-09 0.0007 9.033e-09 0 9.227e-09 0 9.23e-09 0.0007 9.233e-09 0 9.427e-09 0 9.43e-09 0.0007 9.433e-09 0 9.627e-09 0 9.63e-09 0.0007 9.633e-09 0 9.827e-09 0 9.83e-09 0.0007 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0007 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0007 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0007 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0007 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0007 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0007 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0007 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0007 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0007 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0007 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0007 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0007 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0007 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0007 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0007 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0007 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0007 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0007 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0007 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0007 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0007 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0007 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0007 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0007 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0007 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0007 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0007 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0007 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0007 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0007 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0007 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0007 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0007 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0007 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0007 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0007 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0007 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0007 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0007 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0007 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0007 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0007 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0007 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0007 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0007 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0007 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0007 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0007 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0007 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0007 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0007 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0007 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0007 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0007 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0007 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0007 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0007 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0007 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0007 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0007 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0007 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0007 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0007 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0007 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0007 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0007 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0007 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0007 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0007 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0007 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0007 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0007 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0007 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0007 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0007 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0007 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0007 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0007 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0007 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0007 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0007 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0007 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0007 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0007 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0007 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0007 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0007 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0007 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0007 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0007 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0007 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0007 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0007 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0007 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0007 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0007 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0007 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0007 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0007 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0007 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0007 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0007 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0007 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0007 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0007 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0007 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0007 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0007 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0007 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0007 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0007 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0007 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0007 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0007 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0007 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0007 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0007 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0007 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0007 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0007 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0007 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0007 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0007 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0007 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0007 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0007 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0007 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0007 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0007 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0007 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0007 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0007 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0007 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0007 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0007 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0007 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0007 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0007 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0007 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0007 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0007 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0007 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0007 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0007 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0007 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0007 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0007 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0007 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0007 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0007 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0007 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0007 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0007 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0007 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0007 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0007 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0007 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0007 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0007 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0007 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0007 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0007 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0007 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0007 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0007 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0007 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0007 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0007 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0007 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0007 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0007 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0007 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0007 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0007 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0007 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0007 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0007 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0007 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0007 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0007 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0007 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0007 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0007 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0007 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0007 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0007 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0007 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0007 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0007 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0007 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0007 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0007 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0007 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0007 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0007 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0007 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0007 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0007 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0007 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0007 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0007 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0007 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0007 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0007 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0007 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0007 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0007 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0007 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0007 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0007 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0007 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0007 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0007 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0007 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0007 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0007 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0007 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0007 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0007 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0007 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0007 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0007 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0007 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0007 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0007 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0007 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0007 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0007 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0007 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0007 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0007 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0007 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0007 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0007 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0007 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0007 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0007 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0007 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0007 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0007 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0007 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0007 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0007 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0007 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0007 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0007 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0007 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0007 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0007 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0007 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0007 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0007 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0007 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0007 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0007 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0007 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0007 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0007 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0007 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0007 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0007 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0007 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0007 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0007 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0007 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0007 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0007 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0007 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0007 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0007 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0007 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0007 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0007 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0007 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0007 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0007 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0007 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0007 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0007 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0007 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0007 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0007 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0007 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0007 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0007 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0007 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0007 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0007 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0007 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0007 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0007 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0007 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0007 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0007 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0007 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0007 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0007 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0007 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0007 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0007 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0007 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0007 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0007 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0007 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0007 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0007 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0007 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0007 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0007 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0007 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0007 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0007 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0007 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0007 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0007 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0007 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0007 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0007 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0007 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0007 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0007 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0007 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0007 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0007 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0007 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0007 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0007 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0007 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0007 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0007 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0007 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0007 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0007 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0007 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0007 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0007 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0007 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0007 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0007 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0007 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0007 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0007 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0007 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0007 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0007 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0007 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0007 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0007 7.9633e-08 0)
L_IP5_OUT|1 IP5_0_OUT _IP5_OUT|A1  2.067833848e-12
L_IP5_OUT|2 _IP5_OUT|A1 _IP5_OUT|A2  4.135667696e-12
L_IP5_OUT|3 _IP5_OUT|A3 _IP5_OUT|A4  8.271335392e-12
L_IP5_OUT|T T18 _IP5_OUT|T1  2.067833848e-12
L_IP5_OUT|4 _IP5_OUT|T1 _IP5_OUT|T2  4.135667696e-12
L_IP5_OUT|5 _IP5_OUT|A4 _IP5_OUT|Q1  4.135667696e-12
L_IP5_OUT|6 _IP5_OUT|Q1 IP5_1_OUT_TX  2.067833848e-12
IT19|T 0 T19  PWL(0 0 2.7e-11 0 3e-11 0.0014 3.3e-11 0 2.27e-10 0 2.3e-10 0.0014 2.33e-10 0 4.27e-10 0 4.3e-10 0.0014 4.33e-10 0 6.27e-10 0 6.3e-10 0.0014 6.33e-10 0 8.27e-10 0 8.3e-10 0.0014 8.33e-10 0 1.027e-09 0 1.03e-09 0.0014 1.033e-09 0 1.227e-09 0 1.23e-09 0.0014 1.233e-09 0 1.427e-09 0 1.43e-09 0.0014 1.433e-09 0 1.627e-09 0 1.63e-09 0.0014 1.633e-09 0 1.827e-09 0 1.83e-09 0.0014 1.833e-09 0 2.027e-09 0 2.03e-09 0.0014 2.033e-09 0 2.227e-09 0 2.23e-09 0.0014 2.233e-09 0 2.427e-09 0 2.43e-09 0.0014 2.433e-09 0 2.627e-09 0 2.63e-09 0.0014 2.633e-09 0 2.827e-09 0 2.83e-09 0.0014 2.833e-09 0 3.027e-09 0 3.03e-09 0.0014 3.033e-09 0 3.227e-09 0 3.23e-09 0.0014 3.233e-09 0 3.427e-09 0 3.43e-09 0.0014 3.433e-09 0 3.627e-09 0 3.63e-09 0.0014 3.633e-09 0 3.827e-09 0 3.83e-09 0.0014 3.833e-09 0 4.027e-09 0 4.03e-09 0.0014 4.033e-09 0 4.227e-09 0 4.23e-09 0.0014 4.233e-09 0 4.427e-09 0 4.43e-09 0.0014 4.433e-09 0 4.627e-09 0 4.63e-09 0.0014 4.633e-09 0 4.827e-09 0 4.83e-09 0.0014 4.833e-09 0 5.027e-09 0 5.03e-09 0.0014 5.033e-09 0 5.227e-09 0 5.23e-09 0.0014 5.233e-09 0 5.427e-09 0 5.43e-09 0.0014 5.433e-09 0 5.627e-09 0 5.63e-09 0.0014 5.633e-09 0 5.827e-09 0 5.83e-09 0.0014 5.833e-09 0 6.027e-09 0 6.03e-09 0.0014 6.033e-09 0 6.227e-09 0 6.23e-09 0.0014 6.233e-09 0 6.427e-09 0 6.43e-09 0.0014 6.433e-09 0 6.627e-09 0 6.63e-09 0.0014 6.633e-09 0 6.827e-09 0 6.83e-09 0.0014 6.833e-09 0 7.027e-09 0 7.03e-09 0.0014 7.033e-09 0 7.227e-09 0 7.23e-09 0.0014 7.233e-09 0 7.427e-09 0 7.43e-09 0.0014 7.433e-09 0 7.627e-09 0 7.63e-09 0.0014 7.633e-09 0 7.827e-09 0 7.83e-09 0.0014 7.833e-09 0 8.027e-09 0 8.03e-09 0.0014 8.033e-09 0 8.227e-09 0 8.23e-09 0.0014 8.233e-09 0 8.427e-09 0 8.43e-09 0.0014 8.433e-09 0 8.627e-09 0 8.63e-09 0.0014 8.633e-09 0 8.827e-09 0 8.83e-09 0.0014 8.833e-09 0 9.027e-09 0 9.03e-09 0.0014 9.033e-09 0 9.227e-09 0 9.23e-09 0.0014 9.233e-09 0 9.427e-09 0 9.43e-09 0.0014 9.433e-09 0 9.627e-09 0 9.63e-09 0.0014 9.633e-09 0 9.827e-09 0 9.83e-09 0.0014 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0014 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0014 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0014 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0014 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0014 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0014 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0014 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0014 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0014 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0014 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0014 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0014 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0014 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0014 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0014 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0014 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0014 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0014 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0014 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0014 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0014 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0014 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0014 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0014 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0014 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0014 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0014 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0014 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0014 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0014 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0014 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0014 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0014 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0014 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0014 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0014 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0014 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0014 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0014 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0014 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0014 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0014 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0014 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0014 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0014 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0014 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0014 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0014 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0014 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0014 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0014 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0014 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0014 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0014 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0014 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0014 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0014 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0014 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0014 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0014 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0014 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0014 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0014 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0014 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0014 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0014 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0014 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0014 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0014 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0014 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0014 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0014 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0014 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0014 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0014 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0014 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0014 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0014 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0014 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0014 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0014 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0014 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0014 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0014 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0014 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0014 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0014 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0014 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0014 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0014 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0014 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0014 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0014 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0014 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0014 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0014 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0014 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0014 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0014 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0014 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0014 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0014 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0014 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0014 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0014 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0014 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0014 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0014 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0014 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0014 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0014 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0014 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0014 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0014 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0014 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0014 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0014 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0014 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0014 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0014 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0014 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0014 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0014 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0014 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0014 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0014 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0014 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0014 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0014 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0014 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0014 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0014 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0014 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0014 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0014 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0014 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0014 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0014 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0014 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0014 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0014 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0014 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0014 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0014 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0014 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0014 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0014 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0014 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0014 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0014 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0014 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0014 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0014 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0014 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0014 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0014 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0014 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0014 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0014 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0014 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0014 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0014 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0014 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0014 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0014 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0014 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0014 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0014 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0014 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0014 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0014 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0014 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0014 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0014 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0014 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0014 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0014 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0014 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0014 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0014 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0014 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0014 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0014 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0014 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0014 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0014 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0014 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0014 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0014 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0014 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0014 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0014 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0014 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0014 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0014 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0014 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0014 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0014 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0014 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0014 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0014 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0014 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0014 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0014 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0014 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0014 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0014 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0014 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0014 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0014 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0014 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0014 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0014 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0014 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0014 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0014 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0014 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0014 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0014 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0014 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0014 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0014 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0014 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0014 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0014 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0014 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0014 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0014 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0014 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0014 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0014 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0014 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0014 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0014 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0014 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0014 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0014 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0014 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0014 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0014 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0014 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0014 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0014 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0014 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0014 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0014 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0014 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0014 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0014 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0014 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0014 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0014 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0014 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0014 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0014 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0014 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0014 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0014 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0014 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0014 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0014 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0014 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0014 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0014 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0014 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0014 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0014 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0014 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0014 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0014 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0014 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0014 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0014 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0014 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0014 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0014 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0014 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0014 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0014 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0014 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0014 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0014 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0014 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0014 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0014 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0014 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0014 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0014 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0014 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0014 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0014 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0014 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0014 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0014 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0014 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0014 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0014 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0014 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0014 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0014 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0014 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0014 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0014 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0014 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0014 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0014 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0014 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0014 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0014 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0014 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0014 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0014 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0014 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0014 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0014 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0014 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0014 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0014 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0014 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0014 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0014 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0014 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0014 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0014 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0014 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0014 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0014 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0014 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0014 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0014 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0014 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0014 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0014 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0014 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0014 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0014 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0014 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0014 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0014 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0014 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0014 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0014 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0014 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0014 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0014 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0014 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0014 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0014 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0014 7.9633e-08 0)
IT1A|T 0 T1A  PWL(0 0 2.7e-11 0 3e-11 0.0028 3.3e-11 0 2.27e-10 0 2.3e-10 0.0028 2.33e-10 0 4.27e-10 0 4.3e-10 0.0028 4.33e-10 0 6.27e-10 0 6.3e-10 0.0028 6.33e-10 0 8.27e-10 0 8.3e-10 0.0028 8.33e-10 0 1.027e-09 0 1.03e-09 0.0028 1.033e-09 0 1.227e-09 0 1.23e-09 0.0028 1.233e-09 0 1.427e-09 0 1.43e-09 0.0028 1.433e-09 0 1.627e-09 0 1.63e-09 0.0028 1.633e-09 0 1.827e-09 0 1.83e-09 0.0028 1.833e-09 0 2.027e-09 0 2.03e-09 0.0028 2.033e-09 0 2.227e-09 0 2.23e-09 0.0028 2.233e-09 0 2.427e-09 0 2.43e-09 0.0028 2.433e-09 0 2.627e-09 0 2.63e-09 0.0028 2.633e-09 0 2.827e-09 0 2.83e-09 0.0028 2.833e-09 0 3.027e-09 0 3.03e-09 0.0028 3.033e-09 0 3.227e-09 0 3.23e-09 0.0028 3.233e-09 0 3.427e-09 0 3.43e-09 0.0028 3.433e-09 0 3.627e-09 0 3.63e-09 0.0028 3.633e-09 0 3.827e-09 0 3.83e-09 0.0028 3.833e-09 0 4.027e-09 0 4.03e-09 0.0028 4.033e-09 0 4.227e-09 0 4.23e-09 0.0028 4.233e-09 0 4.427e-09 0 4.43e-09 0.0028 4.433e-09 0 4.627e-09 0 4.63e-09 0.0028 4.633e-09 0 4.827e-09 0 4.83e-09 0.0028 4.833e-09 0 5.027e-09 0 5.03e-09 0.0028 5.033e-09 0 5.227e-09 0 5.23e-09 0.0028 5.233e-09 0 5.427e-09 0 5.43e-09 0.0028 5.433e-09 0 5.627e-09 0 5.63e-09 0.0028 5.633e-09 0 5.827e-09 0 5.83e-09 0.0028 5.833e-09 0 6.027e-09 0 6.03e-09 0.0028 6.033e-09 0 6.227e-09 0 6.23e-09 0.0028 6.233e-09 0 6.427e-09 0 6.43e-09 0.0028 6.433e-09 0 6.627e-09 0 6.63e-09 0.0028 6.633e-09 0 6.827e-09 0 6.83e-09 0.0028 6.833e-09 0 7.027e-09 0 7.03e-09 0.0028 7.033e-09 0 7.227e-09 0 7.23e-09 0.0028 7.233e-09 0 7.427e-09 0 7.43e-09 0.0028 7.433e-09 0 7.627e-09 0 7.63e-09 0.0028 7.633e-09 0 7.827e-09 0 7.83e-09 0.0028 7.833e-09 0 8.027e-09 0 8.03e-09 0.0028 8.033e-09 0 8.227e-09 0 8.23e-09 0.0028 8.233e-09 0 8.427e-09 0 8.43e-09 0.0028 8.433e-09 0 8.627e-09 0 8.63e-09 0.0028 8.633e-09 0 8.827e-09 0 8.83e-09 0.0028 8.833e-09 0 9.027e-09 0 9.03e-09 0.0028 9.033e-09 0 9.227e-09 0 9.23e-09 0.0028 9.233e-09 0 9.427e-09 0 9.43e-09 0.0028 9.433e-09 0 9.627e-09 0 9.63e-09 0.0028 9.633e-09 0 9.827e-09 0 9.83e-09 0.0028 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0028 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0028 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0028 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0028 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0028 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0028 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0028 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0028 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0028 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0028 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0028 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0028 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0028 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0028 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0028 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0028 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0028 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0028 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0028 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0028 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0028 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0028 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0028 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0028 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0028 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0028 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0028 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0028 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0028 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0028 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0028 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0028 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0028 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0028 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0028 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0028 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0028 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0028 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0028 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0028 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0028 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0028 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0028 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0028 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0028 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0028 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0028 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0028 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0028 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0028 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0028 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0028 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0028 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0028 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0028 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0028 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0028 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0028 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0028 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0028 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0028 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0028 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0028 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0028 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0028 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0028 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0028 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0028 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0028 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0028 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0028 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0028 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0028 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0028 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0028 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0028 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0028 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0028 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0028 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0028 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0028 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0028 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0028 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0028 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0028 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0028 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0028 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0028 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0028 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0028 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0028 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0028 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0028 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0028 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0028 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0028 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0028 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0028 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0028 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0028 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0028 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0028 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0028 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0028 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0028 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0028 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0028 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0028 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0028 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0028 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0028 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0028 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0028 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0028 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0028 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0028 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0028 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0028 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0028 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0028 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0028 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0028 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0028 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0028 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0028 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0028 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0028 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0028 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0028 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0028 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0028 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0028 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0028 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0028 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0028 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0028 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0028 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0028 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0028 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0028 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0028 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0028 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0028 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0028 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0028 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0028 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0028 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0028 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0028 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0028 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0028 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0028 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0028 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0028 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0028 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0028 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0028 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0028 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0028 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0028 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0028 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0028 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0028 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0028 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0028 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0028 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0028 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0028 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0028 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0028 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0028 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0028 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0028 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0028 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0028 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0028 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0028 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0028 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0028 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0028 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0028 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0028 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0028 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0028 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0028 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0028 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0028 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0028 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0028 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0028 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0028 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0028 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0028 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0028 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0028 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0028 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0028 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0028 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0028 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0028 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0028 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0028 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0028 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0028 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0028 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0028 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0028 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0028 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0028 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0028 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0028 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0028 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0028 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0028 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0028 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0028 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0028 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0028 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0028 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0028 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0028 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0028 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0028 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0028 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0028 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0028 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0028 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0028 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0028 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0028 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0028 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0028 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0028 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0028 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0028 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0028 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0028 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0028 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0028 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0028 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0028 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0028 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0028 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0028 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0028 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0028 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0028 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0028 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0028 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0028 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0028 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0028 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0028 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0028 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0028 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0028 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0028 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0028 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0028 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0028 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0028 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0028 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0028 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0028 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0028 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0028 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0028 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0028 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0028 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0028 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0028 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0028 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0028 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0028 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0028 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0028 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0028 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0028 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0028 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0028 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0028 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0028 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0028 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0028 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0028 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0028 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0028 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0028 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0028 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0028 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0028 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0028 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0028 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0028 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0028 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0028 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0028 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0028 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0028 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0028 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0028 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0028 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0028 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0028 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0028 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0028 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0028 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0028 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0028 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0028 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0028 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0028 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0028 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0028 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0028 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0028 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0028 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0028 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0028 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0028 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0028 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0028 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0028 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0028 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0028 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0028 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0028 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0028 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0028 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0028 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0028 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0028 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0028 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0028 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0028 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0028 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0028 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0028 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0028 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0028 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0028 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0028 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0028 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0028 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0028 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0028 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0028 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0028 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0028 7.9633e-08 0)
IT1B|T 0 T21  PWL(0 0 2.7e-11 0 3e-11 0.0007 3.3e-11 0 2.27e-10 0 2.3e-10 0.0007 2.33e-10 0 4.27e-10 0 4.3e-10 0.0007 4.33e-10 0 6.27e-10 0 6.3e-10 0.0007 6.33e-10 0 8.27e-10 0 8.3e-10 0.0007 8.33e-10 0 1.027e-09 0 1.03e-09 0.0007 1.033e-09 0 1.227e-09 0 1.23e-09 0.0007 1.233e-09 0 1.427e-09 0 1.43e-09 0.0007 1.433e-09 0 1.627e-09 0 1.63e-09 0.0007 1.633e-09 0 1.827e-09 0 1.83e-09 0.0007 1.833e-09 0 2.027e-09 0 2.03e-09 0.0007 2.033e-09 0 2.227e-09 0 2.23e-09 0.0007 2.233e-09 0 2.427e-09 0 2.43e-09 0.0007 2.433e-09 0 2.627e-09 0 2.63e-09 0.0007 2.633e-09 0 2.827e-09 0 2.83e-09 0.0007 2.833e-09 0 3.027e-09 0 3.03e-09 0.0007 3.033e-09 0 3.227e-09 0 3.23e-09 0.0007 3.233e-09 0 3.427e-09 0 3.43e-09 0.0007 3.433e-09 0 3.627e-09 0 3.63e-09 0.0007 3.633e-09 0 3.827e-09 0 3.83e-09 0.0007 3.833e-09 0 4.027e-09 0 4.03e-09 0.0007 4.033e-09 0 4.227e-09 0 4.23e-09 0.0007 4.233e-09 0 4.427e-09 0 4.43e-09 0.0007 4.433e-09 0 4.627e-09 0 4.63e-09 0.0007 4.633e-09 0 4.827e-09 0 4.83e-09 0.0007 4.833e-09 0 5.027e-09 0 5.03e-09 0.0007 5.033e-09 0 5.227e-09 0 5.23e-09 0.0007 5.233e-09 0 5.427e-09 0 5.43e-09 0.0007 5.433e-09 0 5.627e-09 0 5.63e-09 0.0007 5.633e-09 0 5.827e-09 0 5.83e-09 0.0007 5.833e-09 0 6.027e-09 0 6.03e-09 0.0007 6.033e-09 0 6.227e-09 0 6.23e-09 0.0007 6.233e-09 0 6.427e-09 0 6.43e-09 0.0007 6.433e-09 0 6.627e-09 0 6.63e-09 0.0007 6.633e-09 0 6.827e-09 0 6.83e-09 0.0007 6.833e-09 0 7.027e-09 0 7.03e-09 0.0007 7.033e-09 0 7.227e-09 0 7.23e-09 0.0007 7.233e-09 0 7.427e-09 0 7.43e-09 0.0007 7.433e-09 0 7.627e-09 0 7.63e-09 0.0007 7.633e-09 0 7.827e-09 0 7.83e-09 0.0007 7.833e-09 0 8.027e-09 0 8.03e-09 0.0007 8.033e-09 0 8.227e-09 0 8.23e-09 0.0007 8.233e-09 0 8.427e-09 0 8.43e-09 0.0007 8.433e-09 0 8.627e-09 0 8.63e-09 0.0007 8.633e-09 0 8.827e-09 0 8.83e-09 0.0007 8.833e-09 0 9.027e-09 0 9.03e-09 0.0007 9.033e-09 0 9.227e-09 0 9.23e-09 0.0007 9.233e-09 0 9.427e-09 0 9.43e-09 0.0007 9.433e-09 0 9.627e-09 0 9.63e-09 0.0007 9.633e-09 0 9.827e-09 0 9.83e-09 0.0007 9.833e-09 0 1.0027e-08 0 1.003e-08 0.0007 1.0033e-08 0 1.0227e-08 0 1.023e-08 0.0007 1.0233e-08 0 1.0427e-08 0 1.043e-08 0.0007 1.0433e-08 0 1.0627e-08 0 1.063e-08 0.0007 1.0633e-08 0 1.0827e-08 0 1.083e-08 0.0007 1.0833e-08 0 1.1027e-08 0 1.103e-08 0.0007 1.1033e-08 0 1.1227e-08 0 1.123e-08 0.0007 1.1233e-08 0 1.1427e-08 0 1.143e-08 0.0007 1.1433e-08 0 1.1627e-08 0 1.163e-08 0.0007 1.1633e-08 0 1.1827e-08 0 1.183e-08 0.0007 1.1833e-08 0 1.2027e-08 0 1.203e-08 0.0007 1.2033e-08 0 1.2227e-08 0 1.223e-08 0.0007 1.2233e-08 0 1.2427e-08 0 1.243e-08 0.0007 1.2433e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2827e-08 0 1.283e-08 0.0007 1.2833e-08 0 1.3027e-08 0 1.303e-08 0.0007 1.3033e-08 0 1.3227e-08 0 1.323e-08 0.0007 1.3233e-08 0 1.3427e-08 0 1.343e-08 0.0007 1.3433e-08 0 1.3627e-08 0 1.363e-08 0.0007 1.3633e-08 0 1.3827e-08 0 1.383e-08 0.0007 1.3833e-08 0 1.4027e-08 0 1.403e-08 0.0007 1.4033e-08 0 1.4227e-08 0 1.423e-08 0.0007 1.4233e-08 0 1.4427e-08 0 1.443e-08 0.0007 1.4433e-08 0 1.4627e-08 0 1.463e-08 0.0007 1.4633e-08 0 1.4827e-08 0 1.483e-08 0.0007 1.4833e-08 0 1.5027e-08 0 1.503e-08 0.0007 1.5033e-08 0 1.5227e-08 0 1.523e-08 0.0007 1.5233e-08 0 1.5427e-08 0 1.543e-08 0.0007 1.5433e-08 0 1.5627e-08 0 1.563e-08 0.0007 1.5633e-08 0 1.5827e-08 0 1.583e-08 0.0007 1.5833e-08 0 1.6027e-08 0 1.603e-08 0.0007 1.6033e-08 0 1.6227e-08 0 1.623e-08 0.0007 1.6233e-08 0 1.6427e-08 0 1.643e-08 0.0007 1.6433e-08 0 1.6627e-08 0 1.663e-08 0.0007 1.6633e-08 0 1.6827e-08 0 1.683e-08 0.0007 1.6833e-08 0 1.7027e-08 0 1.703e-08 0.0007 1.7033e-08 0 1.7227e-08 0 1.723e-08 0.0007 1.7233e-08 0 1.7427e-08 0 1.743e-08 0.0007 1.7433e-08 0 1.7627e-08 0 1.763e-08 0.0007 1.7633e-08 0 1.7827e-08 0 1.783e-08 0.0007 1.7833e-08 0 1.8027e-08 0 1.803e-08 0.0007 1.8033e-08 0 1.8227e-08 0 1.823e-08 0.0007 1.8233e-08 0 1.8427e-08 0 1.843e-08 0.0007 1.8433e-08 0 1.8627e-08 0 1.863e-08 0.0007 1.8633e-08 0 1.8827e-08 0 1.883e-08 0.0007 1.8833e-08 0 1.9027e-08 0 1.903e-08 0.0007 1.9033e-08 0 1.9227e-08 0 1.923e-08 0.0007 1.9233e-08 0 1.9427e-08 0 1.943e-08 0.0007 1.9433e-08 0 1.9627e-08 0 1.963e-08 0.0007 1.9633e-08 0 1.9827e-08 0 1.983e-08 0.0007 1.9833e-08 0 2.0027e-08 0 2.003e-08 0.0007 2.0033e-08 0 2.0227e-08 0 2.023e-08 0.0007 2.0233e-08 0 2.0427e-08 0 2.043e-08 0.0007 2.0433e-08 0 2.0627e-08 0 2.063e-08 0.0007 2.0633e-08 0 2.0827e-08 0 2.083e-08 0.0007 2.0833e-08 0 2.1027e-08 0 2.103e-08 0.0007 2.1033e-08 0 2.1227e-08 0 2.123e-08 0.0007 2.1233e-08 0 2.1427e-08 0 2.143e-08 0.0007 2.1433e-08 0 2.1627e-08 0 2.163e-08 0.0007 2.1633e-08 0 2.1827e-08 0 2.183e-08 0.0007 2.1833e-08 0 2.2027e-08 0 2.203e-08 0.0007 2.2033e-08 0 2.2227e-08 0 2.223e-08 0.0007 2.2233e-08 0 2.2427e-08 0 2.243e-08 0.0007 2.2433e-08 0 2.2627e-08 0 2.263e-08 0.0007 2.2633e-08 0 2.2827e-08 0 2.283e-08 0.0007 2.2833e-08 0 2.3027e-08 0 2.303e-08 0.0007 2.3033e-08 0 2.3227e-08 0 2.323e-08 0.0007 2.3233e-08 0 2.3427e-08 0 2.343e-08 0.0007 2.3433e-08 0 2.3627e-08 0 2.363e-08 0.0007 2.3633e-08 0 2.3827e-08 0 2.383e-08 0.0007 2.3833e-08 0 2.4027e-08 0 2.403e-08 0.0007 2.4033e-08 0 2.4227e-08 0 2.423e-08 0.0007 2.4233e-08 0 2.4427e-08 0 2.443e-08 0.0007 2.4433e-08 0 2.4627e-08 0 2.463e-08 0.0007 2.4633e-08 0 2.4827e-08 0 2.483e-08 0.0007 2.4833e-08 0 2.5027e-08 0 2.503e-08 0.0007 2.5033e-08 0 2.5227e-08 0 2.523e-08 0.0007 2.5233e-08 0 2.5427e-08 0 2.543e-08 0.0007 2.5433e-08 0 2.5627e-08 0 2.563e-08 0.0007 2.5633e-08 0 2.5827e-08 0 2.583e-08 0.0007 2.5833e-08 0 2.6027e-08 0 2.603e-08 0.0007 2.6033e-08 0 2.6227e-08 0 2.623e-08 0.0007 2.6233e-08 0 2.6427e-08 0 2.643e-08 0.0007 2.6433e-08 0 2.6627e-08 0 2.663e-08 0.0007 2.6633e-08 0 2.6827e-08 0 2.683e-08 0.0007 2.6833e-08 0 2.7027e-08 0 2.703e-08 0.0007 2.7033e-08 0 2.7227e-08 0 2.723e-08 0.0007 2.7233e-08 0 2.7427e-08 0 2.743e-08 0.0007 2.7433e-08 0 2.7627e-08 0 2.763e-08 0.0007 2.7633e-08 0 2.7827e-08 0 2.783e-08 0.0007 2.7833e-08 0 2.8027e-08 0 2.803e-08 0.0007 2.8033e-08 0 2.8227e-08 0 2.823e-08 0.0007 2.8233e-08 0 2.8427e-08 0 2.843e-08 0.0007 2.8433e-08 0 2.8627e-08 0 2.863e-08 0.0007 2.8633e-08 0 2.8827e-08 0 2.883e-08 0.0007 2.8833e-08 0 2.9027e-08 0 2.903e-08 0.0007 2.9033e-08 0 2.9227e-08 0 2.923e-08 0.0007 2.9233e-08 0 2.9427e-08 0 2.943e-08 0.0007 2.9433e-08 0 2.9627e-08 0 2.963e-08 0.0007 2.9633e-08 0 2.9827e-08 0 2.983e-08 0.0007 2.9833e-08 0 3.0027e-08 0 3.003e-08 0.0007 3.0033e-08 0 3.0227e-08 0 3.023e-08 0.0007 3.0233e-08 0 3.0427e-08 0 3.043e-08 0.0007 3.0433e-08 0 3.0627e-08 0 3.063e-08 0.0007 3.0633e-08 0 3.0827e-08 0 3.083e-08 0.0007 3.0833e-08 0 3.1027e-08 0 3.103e-08 0.0007 3.1033e-08 0 3.1227e-08 0 3.123e-08 0.0007 3.1233e-08 0 3.1427e-08 0 3.143e-08 0.0007 3.1433e-08 0 3.1627e-08 0 3.163e-08 0.0007 3.1633e-08 0 3.1827e-08 0 3.183e-08 0.0007 3.1833e-08 0 3.2027e-08 0 3.203e-08 0.0007 3.2033e-08 0 3.2227e-08 0 3.223e-08 0.0007 3.2233e-08 0 3.2427e-08 0 3.243e-08 0.0007 3.2433e-08 0 3.2627e-08 0 3.263e-08 0.0007 3.2633e-08 0 3.2827e-08 0 3.283e-08 0.0007 3.2833e-08 0 3.3027e-08 0 3.303e-08 0.0007 3.3033e-08 0 3.3227e-08 0 3.323e-08 0.0007 3.3233e-08 0 3.3427e-08 0 3.343e-08 0.0007 3.3433e-08 0 3.3627e-08 0 3.363e-08 0.0007 3.3633e-08 0 3.3827e-08 0 3.383e-08 0.0007 3.3833e-08 0 3.4027e-08 0 3.403e-08 0.0007 3.4033e-08 0 3.4227e-08 0 3.423e-08 0.0007 3.4233e-08 0 3.4427e-08 0 3.443e-08 0.0007 3.4433e-08 0 3.4627e-08 0 3.463e-08 0.0007 3.4633e-08 0 3.4827e-08 0 3.483e-08 0.0007 3.4833e-08 0 3.5027e-08 0 3.503e-08 0.0007 3.5033e-08 0 3.5227e-08 0 3.523e-08 0.0007 3.5233e-08 0 3.5427e-08 0 3.543e-08 0.0007 3.5433e-08 0 3.5627e-08 0 3.563e-08 0.0007 3.5633e-08 0 3.5827e-08 0 3.583e-08 0.0007 3.5833e-08 0 3.6027e-08 0 3.603e-08 0.0007 3.6033e-08 0 3.6227e-08 0 3.623e-08 0.0007 3.6233e-08 0 3.6427e-08 0 3.643e-08 0.0007 3.6433e-08 0 3.6627e-08 0 3.663e-08 0.0007 3.6633e-08 0 3.6827e-08 0 3.683e-08 0.0007 3.6833e-08 0 3.7027e-08 0 3.703e-08 0.0007 3.7033e-08 0 3.7227e-08 0 3.723e-08 0.0007 3.7233e-08 0 3.7427e-08 0 3.743e-08 0.0007 3.7433e-08 0 3.7627e-08 0 3.763e-08 0.0007 3.7633e-08 0 3.7827e-08 0 3.783e-08 0.0007 3.7833e-08 0 3.8027e-08 0 3.803e-08 0.0007 3.8033e-08 0 3.8227e-08 0 3.823e-08 0.0007 3.8233e-08 0 3.8427e-08 0 3.843e-08 0.0007 3.8433e-08 0 3.8627e-08 0 3.863e-08 0.0007 3.8633e-08 0 3.8827e-08 0 3.883e-08 0.0007 3.8833e-08 0 3.9027e-08 0 3.903e-08 0.0007 3.9033e-08 0 3.9227e-08 0 3.923e-08 0.0007 3.9233e-08 0 3.9427e-08 0 3.943e-08 0.0007 3.9433e-08 0 3.9627e-08 0 3.963e-08 0.0007 3.9633e-08 0 3.9827e-08 0 3.983e-08 0.0007 3.9833e-08 0 4.0027e-08 0 4.003e-08 0.0007 4.0033e-08 0 4.0227e-08 0 4.023e-08 0.0007 4.0233e-08 0 4.0427e-08 0 4.043e-08 0.0007 4.0433e-08 0 4.0627e-08 0 4.063e-08 0.0007 4.0633e-08 0 4.0827e-08 0 4.083e-08 0.0007 4.0833e-08 0 4.1027e-08 0 4.103e-08 0.0007 4.1033e-08 0 4.1227e-08 0 4.123e-08 0.0007 4.1233e-08 0 4.1427e-08 0 4.143e-08 0.0007 4.1433e-08 0 4.1627e-08 0 4.163e-08 0.0007 4.1633e-08 0 4.1827e-08 0 4.183e-08 0.0007 4.1833e-08 0 4.2027e-08 0 4.203e-08 0.0007 4.2033e-08 0 4.2227e-08 0 4.223e-08 0.0007 4.2233e-08 0 4.2427e-08 0 4.243e-08 0.0007 4.2433e-08 0 4.2627e-08 0 4.263e-08 0.0007 4.2633e-08 0 4.2827e-08 0 4.283e-08 0.0007 4.2833e-08 0 4.3027e-08 0 4.303e-08 0.0007 4.3033e-08 0 4.3227e-08 0 4.323e-08 0.0007 4.3233e-08 0 4.3427e-08 0 4.343e-08 0.0007 4.3433e-08 0 4.3627e-08 0 4.363e-08 0.0007 4.3633e-08 0 4.3827e-08 0 4.383e-08 0.0007 4.3833e-08 0 4.4027e-08 0 4.403e-08 0.0007 4.4033e-08 0 4.4227e-08 0 4.423e-08 0.0007 4.4233e-08 0 4.4427e-08 0 4.443e-08 0.0007 4.4433e-08 0 4.4627e-08 0 4.463e-08 0.0007 4.4633e-08 0 4.4827e-08 0 4.483e-08 0.0007 4.4833e-08 0 4.5027e-08 0 4.503e-08 0.0007 4.5033e-08 0 4.5227e-08 0 4.523e-08 0.0007 4.5233e-08 0 4.5427e-08 0 4.543e-08 0.0007 4.5433e-08 0 4.5627e-08 0 4.563e-08 0.0007 4.5633e-08 0 4.5827e-08 0 4.583e-08 0.0007 4.5833e-08 0 4.6027e-08 0 4.603e-08 0.0007 4.6033e-08 0 4.6227e-08 0 4.623e-08 0.0007 4.6233e-08 0 4.6427e-08 0 4.643e-08 0.0007 4.6433e-08 0 4.6627e-08 0 4.663e-08 0.0007 4.6633e-08 0 4.6827e-08 0 4.683e-08 0.0007 4.6833e-08 0 4.7027e-08 0 4.703e-08 0.0007 4.7033e-08 0 4.7227e-08 0 4.723e-08 0.0007 4.7233e-08 0 4.7427e-08 0 4.743e-08 0.0007 4.7433e-08 0 4.7627e-08 0 4.763e-08 0.0007 4.7633e-08 0 4.7827e-08 0 4.783e-08 0.0007 4.7833e-08 0 4.8027e-08 0 4.803e-08 0.0007 4.8033e-08 0 4.8227e-08 0 4.823e-08 0.0007 4.8233e-08 0 4.8427e-08 0 4.843e-08 0.0007 4.8433e-08 0 4.8627e-08 0 4.863e-08 0.0007 4.8633e-08 0 4.8827e-08 0 4.883e-08 0.0007 4.8833e-08 0 4.9027e-08 0 4.903e-08 0.0007 4.9033e-08 0 4.9227e-08 0 4.923e-08 0.0007 4.9233e-08 0 4.9427e-08 0 4.943e-08 0.0007 4.9433e-08 0 4.9627e-08 0 4.963e-08 0.0007 4.9633e-08 0 4.9827e-08 0 4.983e-08 0.0007 4.9833e-08 0 5.0027e-08 0 5.003e-08 0.0007 5.0033e-08 0 5.0227e-08 0 5.023e-08 0.0007 5.0233e-08 0 5.0427e-08 0 5.043e-08 0.0007 5.0433e-08 0 5.0627e-08 0 5.063e-08 0.0007 5.0633e-08 0 5.0827e-08 0 5.083e-08 0.0007 5.0833e-08 0 5.1027e-08 0 5.103e-08 0.0007 5.1033e-08 0 5.1227e-08 0 5.123e-08 0.0007 5.1233e-08 0 5.1427e-08 0 5.143e-08 0.0007 5.1433e-08 0 5.1627e-08 0 5.163e-08 0.0007 5.1633e-08 0 5.1827e-08 0 5.183e-08 0.0007 5.1833e-08 0 5.2027e-08 0 5.203e-08 0.0007 5.2033e-08 0 5.2227e-08 0 5.223e-08 0.0007 5.2233e-08 0 5.2427e-08 0 5.243e-08 0.0007 5.2433e-08 0 5.2627e-08 0 5.263e-08 0.0007 5.2633e-08 0 5.2827e-08 0 5.283e-08 0.0007 5.2833e-08 0 5.3027e-08 0 5.303e-08 0.0007 5.3033e-08 0 5.3227e-08 0 5.323e-08 0.0007 5.3233e-08 0 5.3427e-08 0 5.343e-08 0.0007 5.3433e-08 0 5.3627e-08 0 5.363e-08 0.0007 5.3633e-08 0 5.3827e-08 0 5.383e-08 0.0007 5.3833e-08 0 5.4027e-08 0 5.403e-08 0.0007 5.4033e-08 0 5.4227e-08 0 5.423e-08 0.0007 5.4233e-08 0 5.4427e-08 0 5.443e-08 0.0007 5.4433e-08 0 5.4627e-08 0 5.463e-08 0.0007 5.4633e-08 0 5.4827e-08 0 5.483e-08 0.0007 5.4833e-08 0 5.5027e-08 0 5.503e-08 0.0007 5.5033e-08 0 5.5227e-08 0 5.523e-08 0.0007 5.5233e-08 0 5.5427e-08 0 5.543e-08 0.0007 5.5433e-08 0 5.5627e-08 0 5.563e-08 0.0007 5.5633e-08 0 5.5827e-08 0 5.583e-08 0.0007 5.5833e-08 0 5.6027e-08 0 5.603e-08 0.0007 5.6033e-08 0 5.6227e-08 0 5.623e-08 0.0007 5.6233e-08 0 5.6427e-08 0 5.643e-08 0.0007 5.6433e-08 0 5.6627e-08 0 5.663e-08 0.0007 5.6633e-08 0 5.6827e-08 0 5.683e-08 0.0007 5.6833e-08 0 5.7027e-08 0 5.703e-08 0.0007 5.7033e-08 0 5.7227e-08 0 5.723e-08 0.0007 5.7233e-08 0 5.7427e-08 0 5.743e-08 0.0007 5.7433e-08 0 5.7627e-08 0 5.763e-08 0.0007 5.7633e-08 0 5.7827e-08 0 5.783e-08 0.0007 5.7833e-08 0 5.8027e-08 0 5.803e-08 0.0007 5.8033e-08 0 5.8227e-08 0 5.823e-08 0.0007 5.8233e-08 0 5.8427e-08 0 5.843e-08 0.0007 5.8433e-08 0 5.8627e-08 0 5.863e-08 0.0007 5.8633e-08 0 5.8827e-08 0 5.883e-08 0.0007 5.8833e-08 0 5.9027e-08 0 5.903e-08 0.0007 5.9033e-08 0 5.9227e-08 0 5.923e-08 0.0007 5.9233e-08 0 5.9427e-08 0 5.943e-08 0.0007 5.9433e-08 0 5.9627e-08 0 5.963e-08 0.0007 5.9633e-08 0 5.9827e-08 0 5.983e-08 0.0007 5.9833e-08 0 6.0027e-08 0 6.003e-08 0.0007 6.0033e-08 0 6.0227e-08 0 6.023e-08 0.0007 6.0233e-08 0 6.0427e-08 0 6.043e-08 0.0007 6.0433e-08 0 6.0627e-08 0 6.063e-08 0.0007 6.0633e-08 0 6.0827e-08 0 6.083e-08 0.0007 6.0833e-08 0 6.1027e-08 0 6.103e-08 0.0007 6.1033e-08 0 6.1227e-08 0 6.123e-08 0.0007 6.1233e-08 0 6.1427e-08 0 6.143e-08 0.0007 6.1433e-08 0 6.1627e-08 0 6.163e-08 0.0007 6.1633e-08 0 6.1827e-08 0 6.183e-08 0.0007 6.1833e-08 0 6.2027e-08 0 6.203e-08 0.0007 6.2033e-08 0 6.2227e-08 0 6.223e-08 0.0007 6.2233e-08 0 6.2427e-08 0 6.243e-08 0.0007 6.2433e-08 0 6.2627e-08 0 6.263e-08 0.0007 6.2633e-08 0 6.2827e-08 0 6.283e-08 0.0007 6.2833e-08 0 6.3027e-08 0 6.303e-08 0.0007 6.3033e-08 0 6.3227e-08 0 6.323e-08 0.0007 6.3233e-08 0 6.3427e-08 0 6.343e-08 0.0007 6.3433e-08 0 6.3627e-08 0 6.363e-08 0.0007 6.3633e-08 0 6.3827e-08 0 6.383e-08 0.0007 6.3833e-08 0 6.4027e-08 0 6.403e-08 0.0007 6.4033e-08 0 6.4227e-08 0 6.423e-08 0.0007 6.4233e-08 0 6.4427e-08 0 6.443e-08 0.0007 6.4433e-08 0 6.4627e-08 0 6.463e-08 0.0007 6.4633e-08 0 6.4827e-08 0 6.483e-08 0.0007 6.4833e-08 0 6.5027e-08 0 6.503e-08 0.0007 6.5033e-08 0 6.5227e-08 0 6.523e-08 0.0007 6.5233e-08 0 6.5427e-08 0 6.543e-08 0.0007 6.5433e-08 0 6.5627e-08 0 6.563e-08 0.0007 6.5633e-08 0 6.5827e-08 0 6.583e-08 0.0007 6.5833e-08 0 6.6027e-08 0 6.603e-08 0.0007 6.6033e-08 0 6.6227e-08 0 6.623e-08 0.0007 6.6233e-08 0 6.6427e-08 0 6.643e-08 0.0007 6.6433e-08 0 6.6627e-08 0 6.663e-08 0.0007 6.6633e-08 0 6.6827e-08 0 6.683e-08 0.0007 6.6833e-08 0 6.7027e-08 0 6.703e-08 0.0007 6.7033e-08 0 6.7227e-08 0 6.723e-08 0.0007 6.7233e-08 0 6.7427e-08 0 6.743e-08 0.0007 6.7433e-08 0 6.7627e-08 0 6.763e-08 0.0007 6.7633e-08 0 6.7827e-08 0 6.783e-08 0.0007 6.7833e-08 0 6.8027e-08 0 6.803e-08 0.0007 6.8033e-08 0 6.8227e-08 0 6.823e-08 0.0007 6.8233e-08 0 6.8427e-08 0 6.843e-08 0.0007 6.8433e-08 0 6.8627e-08 0 6.863e-08 0.0007 6.8633e-08 0 6.8827e-08 0 6.883e-08 0.0007 6.8833e-08 0 6.9027e-08 0 6.903e-08 0.0007 6.9033e-08 0 6.9227e-08 0 6.923e-08 0.0007 6.9233e-08 0 6.9427e-08 0 6.943e-08 0.0007 6.9433e-08 0 6.9627e-08 0 6.963e-08 0.0007 6.9633e-08 0 6.9827e-08 0 6.983e-08 0.0007 6.9833e-08 0 7.0027e-08 0 7.003e-08 0.0007 7.0033e-08 0 7.0227e-08 0 7.023e-08 0.0007 7.0233e-08 0 7.0427e-08 0 7.043e-08 0.0007 7.0433e-08 0 7.0627e-08 0 7.063e-08 0.0007 7.0633e-08 0 7.0827e-08 0 7.083e-08 0.0007 7.0833e-08 0 7.1027e-08 0 7.103e-08 0.0007 7.1033e-08 0 7.1227e-08 0 7.123e-08 0.0007 7.1233e-08 0 7.1427e-08 0 7.143e-08 0.0007 7.1433e-08 0 7.1627e-08 0 7.163e-08 0.0007 7.1633e-08 0 7.1827e-08 0 7.183e-08 0.0007 7.1833e-08 0 7.2027e-08 0 7.203e-08 0.0007 7.2033e-08 0 7.2227e-08 0 7.223e-08 0.0007 7.2233e-08 0 7.2427e-08 0 7.243e-08 0.0007 7.2433e-08 0 7.2627e-08 0 7.263e-08 0.0007 7.2633e-08 0 7.2827e-08 0 7.283e-08 0.0007 7.2833e-08 0 7.3027e-08 0 7.303e-08 0.0007 7.3033e-08 0 7.3227e-08 0 7.323e-08 0.0007 7.3233e-08 0 7.3427e-08 0 7.343e-08 0.0007 7.3433e-08 0 7.3627e-08 0 7.363e-08 0.0007 7.3633e-08 0 7.3827e-08 0 7.383e-08 0.0007 7.3833e-08 0 7.4027e-08 0 7.403e-08 0.0007 7.4033e-08 0 7.4227e-08 0 7.423e-08 0.0007 7.4233e-08 0 7.4427e-08 0 7.443e-08 0.0007 7.4433e-08 0 7.4627e-08 0 7.463e-08 0.0007 7.4633e-08 0 7.4827e-08 0 7.483e-08 0.0007 7.4833e-08 0 7.5027e-08 0 7.503e-08 0.0007 7.5033e-08 0 7.5227e-08 0 7.523e-08 0.0007 7.5233e-08 0 7.5427e-08 0 7.543e-08 0.0007 7.5433e-08 0 7.5627e-08 0 7.563e-08 0.0007 7.5633e-08 0 7.5827e-08 0 7.583e-08 0.0007 7.5833e-08 0 7.6027e-08 0 7.603e-08 0.0007 7.6033e-08 0 7.6227e-08 0 7.623e-08 0.0007 7.6233e-08 0 7.6427e-08 0 7.643e-08 0.0007 7.6433e-08 0 7.6627e-08 0 7.663e-08 0.0007 7.6633e-08 0 7.6827e-08 0 7.683e-08 0.0007 7.6833e-08 0 7.7027e-08 0 7.703e-08 0.0007 7.7033e-08 0 7.7227e-08 0 7.723e-08 0.0007 7.7233e-08 0 7.7427e-08 0 7.743e-08 0.0007 7.7433e-08 0 7.7627e-08 0 7.763e-08 0.0007 7.7633e-08 0 7.7827e-08 0 7.783e-08 0.0007 7.7833e-08 0 7.8027e-08 0 7.803e-08 0.0007 7.8033e-08 0 7.8227e-08 0 7.823e-08 0.0007 7.8233e-08 0 7.8427e-08 0 7.843e-08 0.0007 7.8433e-08 0 7.8627e-08 0 7.863e-08 0.0007 7.8633e-08 0 7.8827e-08 0 7.883e-08 0.0007 7.8833e-08 0 7.9027e-08 0 7.903e-08 0.0007 7.9033e-08 0 7.9227e-08 0 7.923e-08 0.0007 7.9233e-08 0 7.9427e-08 0 7.943e-08 0.0007 7.9433e-08 0 7.9627e-08 0 7.963e-08 0.0007 7.9633e-08 0)
L_IP7_OUT|1 IP7_0_OUT _IP7_OUT|A1  2.067833848e-12
L_IP7_OUT|2 _IP7_OUT|A1 _IP7_OUT|A2  4.135667696e-12
L_IP7_OUT|3 _IP7_OUT|A3 _IP7_OUT|A4  8.271335392e-12
L_IP7_OUT|T T1B _IP7_OUT|T1  2.067833848e-12
L_IP7_OUT|4 _IP7_OUT|T1 _IP7_OUT|T2  4.135667696e-12
L_IP7_OUT|5 _IP7_OUT|A4 _IP7_OUT|Q1  4.135667696e-12
L_IP7_OUT|6 _IP7_OUT|Q1 IP7_1_OUT_TX  2.067833848e-12
IT20|T 0 T20  PWL(0 0 1.7e-11 0 2e-11 0.0007 2.3e-11 0 2.17e-10 0 2.2e-10 0.0007 2.23e-10 0 4.17e-10 0 4.2e-10 0.0007 4.23e-10 0 6.17e-10 0 6.2e-10 0.0007 6.23e-10 0 8.17e-10 0 8.2e-10 0.0007 8.23e-10 0 1.017e-09 0 1.02e-09 0.0007 1.023e-09 0 1.217e-09 0 1.22e-09 0.0007 1.223e-09 0 1.417e-09 0 1.42e-09 0.0007 1.423e-09 0 1.617e-09 0 1.62e-09 0.0007 1.623e-09 0 1.817e-09 0 1.82e-09 0.0007 1.823e-09 0 2.017e-09 0 2.02e-09 0.0007 2.023e-09 0 2.217e-09 0 2.22e-09 0.0007 2.223e-09 0 2.417e-09 0 2.42e-09 0.0007 2.423e-09 0 2.617e-09 0 2.62e-09 0.0007 2.623e-09 0 2.817e-09 0 2.82e-09 0.0007 2.823e-09 0 3.017e-09 0 3.02e-09 0.0007 3.023e-09 0 3.217e-09 0 3.22e-09 0.0007 3.223e-09 0 3.417e-09 0 3.42e-09 0.0007 3.423e-09 0 3.617e-09 0 3.62e-09 0.0007 3.623e-09 0 3.817e-09 0 3.82e-09 0.0007 3.823e-09 0 4.017e-09 0 4.02e-09 0.0007 4.023e-09 0 4.217e-09 0 4.22e-09 0.0007 4.223e-09 0 4.417e-09 0 4.42e-09 0.0007 4.423e-09 0 4.617e-09 0 4.62e-09 0.0007 4.623e-09 0 4.817e-09 0 4.82e-09 0.0007 4.823e-09 0 5.017e-09 0 5.02e-09 0.0007 5.023e-09 0 5.217e-09 0 5.22e-09 0.0007 5.223e-09 0 5.417e-09 0 5.42e-09 0.0007 5.423e-09 0 5.617e-09 0 5.62e-09 0.0007 5.623e-09 0 5.817e-09 0 5.82e-09 0.0007 5.823e-09 0 6.017e-09 0 6.02e-09 0.0007 6.023e-09 0 6.217e-09 0 6.22e-09 0.0007 6.223e-09 0 6.417e-09 0 6.42e-09 0.0007 6.423e-09 0 6.617e-09 0 6.62e-09 0.0007 6.623e-09 0 6.817e-09 0 6.82e-09 0.0007 6.823e-09 0 7.017e-09 0 7.02e-09 0.0007 7.023e-09 0 7.217e-09 0 7.22e-09 0.0007 7.223e-09 0 7.417e-09 0 7.42e-09 0.0007 7.423e-09 0 7.617e-09 0 7.62e-09 0.0007 7.623e-09 0 7.817e-09 0 7.82e-09 0.0007 7.823e-09 0 8.017e-09 0 8.02e-09 0.0007 8.023e-09 0 8.217e-09 0 8.22e-09 0.0007 8.223e-09 0 8.417e-09 0 8.42e-09 0.0007 8.423e-09 0 8.617e-09 0 8.62e-09 0.0007 8.623e-09 0 8.817e-09 0 8.82e-09 0.0007 8.823e-09 0 9.017e-09 0 9.02e-09 0.0007 9.023e-09 0 9.217e-09 0 9.22e-09 0.0007 9.223e-09 0 9.417e-09 0 9.42e-09 0.0007 9.423e-09 0 9.617e-09 0 9.62e-09 0.0007 9.623e-09 0 9.817e-09 0 9.82e-09 0.0007 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0007 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0007 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0007 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0007 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0007 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0007 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0007 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0007 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0007 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0007 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0007 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0007 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0007 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0007 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0007 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0007 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0007 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0007 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0007 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0007 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0007 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0007 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0007 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0007 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0007 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0007 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0007 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0007 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0007 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0007 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0007 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0007 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0007 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0007 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0007 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0007 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0007 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0007 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0007 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0007 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0007 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0007 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0007 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0007 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0007 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0007 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0007 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0007 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0007 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0007 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0007 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0007 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0007 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0007 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0007 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0007 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0007 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0007 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0007 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0007 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0007 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0007 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0007 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0007 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0007 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0007 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0007 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0007 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0007 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0007 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0007 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0007 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0007 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0007 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0007 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0007 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0007 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0007 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0007 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0007 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0007 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0007 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0007 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0007 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0007 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0007 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0007 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0007 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0007 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0007 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0007 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0007 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0007 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0007 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0007 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0007 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0007 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0007 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0007 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0007 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0007 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0007 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0007 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0007 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0007 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0007 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0007 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0007 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0007 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0007 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0007 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0007 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0007 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0007 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0007 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0007 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0007 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0007 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0007 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0007 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0007 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0007 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0007 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0007 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0007 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0007 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0007 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0007 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0007 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0007 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0007 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0007 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0007 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0007 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0007 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0007 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0007 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0007 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0007 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0007 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0007 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0007 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0007 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0007 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0007 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0007 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0007 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0007 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0007 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0007 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0007 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0007 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0007 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0007 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0007 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0007 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0007 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0007 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0007 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0007 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0007 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0007 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0007 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0007 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0007 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0007 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0007 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0007 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0007 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0007 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0007 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0007 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0007 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0007 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0007 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0007 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0007 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0007 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0007 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0007 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0007 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0007 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0007 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0007 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0007 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0007 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0007 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0007 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0007 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0007 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0007 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0007 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0007 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0007 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0007 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0007 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0007 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0007 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0007 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0007 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0007 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0007 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0007 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0007 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0007 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0007 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0007 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0007 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0007 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0007 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0007 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0007 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0007 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0007 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0007 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0007 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0007 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0007 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0007 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0007 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0007 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0007 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0007 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0007 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0007 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0007 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0007 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0007 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0007 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0007 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0007 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0007 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0007 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0007 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0007 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0007 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0007 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0007 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0007 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0007 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0007 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0007 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0007 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0007 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0007 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0007 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0007 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0007 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0007 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0007 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0007 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0007 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0007 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0007 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0007 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0007 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0007 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0007 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0007 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0007 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0007 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0007 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0007 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0007 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0007 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0007 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0007 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0007 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0007 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0007 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0007 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0007 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0007 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0007 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0007 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0007 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0007 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0007 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0007 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0007 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0007 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0007 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0007 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0007 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0007 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0007 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0007 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0007 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0007 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0007 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0007 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0007 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0007 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0007 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0007 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0007 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0007 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0007 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0007 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0007 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0007 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0007 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0007 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0007 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0007 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0007 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0007 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0007 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0007 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0007 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0007 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0007 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0007 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0007 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0007 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0007 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0007 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0007 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0007 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0007 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0007 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0007 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0007 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0007 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0007 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0007 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0007 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0007 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0007 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0007 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0007 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0007 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0007 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0007 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0007 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0007 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0007 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0007 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0007 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0007 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0007 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0007 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0007 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0007 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0007 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0007 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0007 7.9623e-08 0)
L_S0_12|1 S0_1 _S0_12|A1  2.067833848e-12
L_S0_12|2 _S0_12|A1 _S0_12|A2  4.135667696e-12
L_S0_12|3 _S0_12|A3 _S0_12|A4  8.271335392e-12
L_S0_12|T T20 _S0_12|T1  2.067833848e-12
L_S0_12|4 _S0_12|T1 _S0_12|T2  4.135667696e-12
L_S0_12|5 _S0_12|A4 _S0_12|Q1  4.135667696e-12
L_S0_12|6 _S0_12|Q1 S0_2_TX  2.067833848e-12
IT21|T 0 T21  PWL(0 0 1.7e-11 0 2e-11 0.0007 2.3e-11 0 2.17e-10 0 2.2e-10 0.0007 2.23e-10 0 4.17e-10 0 4.2e-10 0.0007 4.23e-10 0 6.17e-10 0 6.2e-10 0.0007 6.23e-10 0 8.17e-10 0 8.2e-10 0.0007 8.23e-10 0 1.017e-09 0 1.02e-09 0.0007 1.023e-09 0 1.217e-09 0 1.22e-09 0.0007 1.223e-09 0 1.417e-09 0 1.42e-09 0.0007 1.423e-09 0 1.617e-09 0 1.62e-09 0.0007 1.623e-09 0 1.817e-09 0 1.82e-09 0.0007 1.823e-09 0 2.017e-09 0 2.02e-09 0.0007 2.023e-09 0 2.217e-09 0 2.22e-09 0.0007 2.223e-09 0 2.417e-09 0 2.42e-09 0.0007 2.423e-09 0 2.617e-09 0 2.62e-09 0.0007 2.623e-09 0 2.817e-09 0 2.82e-09 0.0007 2.823e-09 0 3.017e-09 0 3.02e-09 0.0007 3.023e-09 0 3.217e-09 0 3.22e-09 0.0007 3.223e-09 0 3.417e-09 0 3.42e-09 0.0007 3.423e-09 0 3.617e-09 0 3.62e-09 0.0007 3.623e-09 0 3.817e-09 0 3.82e-09 0.0007 3.823e-09 0 4.017e-09 0 4.02e-09 0.0007 4.023e-09 0 4.217e-09 0 4.22e-09 0.0007 4.223e-09 0 4.417e-09 0 4.42e-09 0.0007 4.423e-09 0 4.617e-09 0 4.62e-09 0.0007 4.623e-09 0 4.817e-09 0 4.82e-09 0.0007 4.823e-09 0 5.017e-09 0 5.02e-09 0.0007 5.023e-09 0 5.217e-09 0 5.22e-09 0.0007 5.223e-09 0 5.417e-09 0 5.42e-09 0.0007 5.423e-09 0 5.617e-09 0 5.62e-09 0.0007 5.623e-09 0 5.817e-09 0 5.82e-09 0.0007 5.823e-09 0 6.017e-09 0 6.02e-09 0.0007 6.023e-09 0 6.217e-09 0 6.22e-09 0.0007 6.223e-09 0 6.417e-09 0 6.42e-09 0.0007 6.423e-09 0 6.617e-09 0 6.62e-09 0.0007 6.623e-09 0 6.817e-09 0 6.82e-09 0.0007 6.823e-09 0 7.017e-09 0 7.02e-09 0.0007 7.023e-09 0 7.217e-09 0 7.22e-09 0.0007 7.223e-09 0 7.417e-09 0 7.42e-09 0.0007 7.423e-09 0 7.617e-09 0 7.62e-09 0.0007 7.623e-09 0 7.817e-09 0 7.82e-09 0.0007 7.823e-09 0 8.017e-09 0 8.02e-09 0.0007 8.023e-09 0 8.217e-09 0 8.22e-09 0.0007 8.223e-09 0 8.417e-09 0 8.42e-09 0.0007 8.423e-09 0 8.617e-09 0 8.62e-09 0.0007 8.623e-09 0 8.817e-09 0 8.82e-09 0.0007 8.823e-09 0 9.017e-09 0 9.02e-09 0.0007 9.023e-09 0 9.217e-09 0 9.22e-09 0.0007 9.223e-09 0 9.417e-09 0 9.42e-09 0.0007 9.423e-09 0 9.617e-09 0 9.62e-09 0.0007 9.623e-09 0 9.817e-09 0 9.82e-09 0.0007 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0007 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0007 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0007 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0007 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0007 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0007 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0007 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0007 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0007 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0007 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0007 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0007 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0007 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0007 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0007 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0007 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0007 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0007 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0007 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0007 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0007 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0007 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0007 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0007 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0007 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0007 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0007 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0007 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0007 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0007 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0007 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0007 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0007 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0007 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0007 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0007 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0007 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0007 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0007 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0007 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0007 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0007 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0007 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0007 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0007 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0007 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0007 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0007 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0007 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0007 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0007 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0007 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0007 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0007 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0007 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0007 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0007 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0007 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0007 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0007 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0007 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0007 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0007 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0007 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0007 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0007 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0007 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0007 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0007 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0007 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0007 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0007 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0007 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0007 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0007 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0007 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0007 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0007 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0007 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0007 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0007 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0007 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0007 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0007 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0007 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0007 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0007 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0007 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0007 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0007 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0007 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0007 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0007 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0007 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0007 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0007 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0007 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0007 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0007 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0007 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0007 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0007 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0007 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0007 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0007 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0007 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0007 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0007 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0007 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0007 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0007 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0007 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0007 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0007 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0007 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0007 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0007 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0007 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0007 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0007 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0007 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0007 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0007 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0007 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0007 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0007 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0007 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0007 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0007 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0007 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0007 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0007 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0007 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0007 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0007 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0007 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0007 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0007 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0007 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0007 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0007 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0007 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0007 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0007 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0007 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0007 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0007 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0007 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0007 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0007 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0007 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0007 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0007 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0007 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0007 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0007 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0007 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0007 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0007 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0007 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0007 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0007 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0007 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0007 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0007 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0007 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0007 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0007 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0007 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0007 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0007 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0007 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0007 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0007 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0007 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0007 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0007 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0007 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0007 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0007 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0007 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0007 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0007 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0007 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0007 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0007 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0007 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0007 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0007 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0007 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0007 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0007 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0007 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0007 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0007 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0007 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0007 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0007 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0007 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0007 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0007 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0007 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0007 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0007 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0007 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0007 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0007 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0007 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0007 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0007 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0007 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0007 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0007 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0007 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0007 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0007 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0007 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0007 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0007 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0007 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0007 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0007 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0007 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0007 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0007 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0007 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0007 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0007 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0007 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0007 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0007 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0007 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0007 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0007 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0007 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0007 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0007 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0007 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0007 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0007 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0007 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0007 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0007 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0007 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0007 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0007 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0007 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0007 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0007 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0007 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0007 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0007 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0007 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0007 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0007 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0007 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0007 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0007 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0007 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0007 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0007 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0007 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0007 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0007 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0007 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0007 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0007 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0007 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0007 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0007 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0007 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0007 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0007 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0007 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0007 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0007 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0007 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0007 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0007 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0007 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0007 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0007 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0007 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0007 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0007 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0007 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0007 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0007 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0007 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0007 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0007 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0007 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0007 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0007 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0007 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0007 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0007 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0007 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0007 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0007 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0007 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0007 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0007 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0007 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0007 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0007 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0007 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0007 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0007 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0007 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0007 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0007 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0007 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0007 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0007 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0007 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0007 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0007 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0007 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0007 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0007 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0007 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0007 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0007 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0007 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0007 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0007 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0007 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0007 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0007 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0007 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0007 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0007 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0007 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0007 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0007 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0007 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0007 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0007 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0007 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0007 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0007 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0007 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0007 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0007 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0007 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0007 7.9623e-08 0)
L_S1_12|1 S1_1 _S1_12|A1  2.067833848e-12
L_S1_12|2 _S1_12|A1 _S1_12|A2  4.135667696e-12
L_S1_12|3 _S1_12|A3 _S1_12|A4  8.271335392e-12
L_S1_12|T T21 _S1_12|T1  2.067833848e-12
L_S1_12|4 _S1_12|T1 _S1_12|T2  4.135667696e-12
L_S1_12|5 _S1_12|A4 _S1_12|Q1  4.135667696e-12
L_S1_12|6 _S1_12|Q1 S1_2_TX  2.067833848e-12
IT22|T 0 T22  PWL(0 0 1.7e-11 0 2e-11 0.0007 2.3e-11 0 2.17e-10 0 2.2e-10 0.0007 2.23e-10 0 4.17e-10 0 4.2e-10 0.0007 4.23e-10 0 6.17e-10 0 6.2e-10 0.0007 6.23e-10 0 8.17e-10 0 8.2e-10 0.0007 8.23e-10 0 1.017e-09 0 1.02e-09 0.0007 1.023e-09 0 1.217e-09 0 1.22e-09 0.0007 1.223e-09 0 1.417e-09 0 1.42e-09 0.0007 1.423e-09 0 1.617e-09 0 1.62e-09 0.0007 1.623e-09 0 1.817e-09 0 1.82e-09 0.0007 1.823e-09 0 2.017e-09 0 2.02e-09 0.0007 2.023e-09 0 2.217e-09 0 2.22e-09 0.0007 2.223e-09 0 2.417e-09 0 2.42e-09 0.0007 2.423e-09 0 2.617e-09 0 2.62e-09 0.0007 2.623e-09 0 2.817e-09 0 2.82e-09 0.0007 2.823e-09 0 3.017e-09 0 3.02e-09 0.0007 3.023e-09 0 3.217e-09 0 3.22e-09 0.0007 3.223e-09 0 3.417e-09 0 3.42e-09 0.0007 3.423e-09 0 3.617e-09 0 3.62e-09 0.0007 3.623e-09 0 3.817e-09 0 3.82e-09 0.0007 3.823e-09 0 4.017e-09 0 4.02e-09 0.0007 4.023e-09 0 4.217e-09 0 4.22e-09 0.0007 4.223e-09 0 4.417e-09 0 4.42e-09 0.0007 4.423e-09 0 4.617e-09 0 4.62e-09 0.0007 4.623e-09 0 4.817e-09 0 4.82e-09 0.0007 4.823e-09 0 5.017e-09 0 5.02e-09 0.0007 5.023e-09 0 5.217e-09 0 5.22e-09 0.0007 5.223e-09 0 5.417e-09 0 5.42e-09 0.0007 5.423e-09 0 5.617e-09 0 5.62e-09 0.0007 5.623e-09 0 5.817e-09 0 5.82e-09 0.0007 5.823e-09 0 6.017e-09 0 6.02e-09 0.0007 6.023e-09 0 6.217e-09 0 6.22e-09 0.0007 6.223e-09 0 6.417e-09 0 6.42e-09 0.0007 6.423e-09 0 6.617e-09 0 6.62e-09 0.0007 6.623e-09 0 6.817e-09 0 6.82e-09 0.0007 6.823e-09 0 7.017e-09 0 7.02e-09 0.0007 7.023e-09 0 7.217e-09 0 7.22e-09 0.0007 7.223e-09 0 7.417e-09 0 7.42e-09 0.0007 7.423e-09 0 7.617e-09 0 7.62e-09 0.0007 7.623e-09 0 7.817e-09 0 7.82e-09 0.0007 7.823e-09 0 8.017e-09 0 8.02e-09 0.0007 8.023e-09 0 8.217e-09 0 8.22e-09 0.0007 8.223e-09 0 8.417e-09 0 8.42e-09 0.0007 8.423e-09 0 8.617e-09 0 8.62e-09 0.0007 8.623e-09 0 8.817e-09 0 8.82e-09 0.0007 8.823e-09 0 9.017e-09 0 9.02e-09 0.0007 9.023e-09 0 9.217e-09 0 9.22e-09 0.0007 9.223e-09 0 9.417e-09 0 9.42e-09 0.0007 9.423e-09 0 9.617e-09 0 9.62e-09 0.0007 9.623e-09 0 9.817e-09 0 9.82e-09 0.0007 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0007 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0007 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0007 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0007 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0007 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0007 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0007 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0007 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0007 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0007 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0007 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0007 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0007 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0007 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0007 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0007 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0007 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0007 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0007 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0007 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0007 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0007 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0007 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0007 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0007 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0007 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0007 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0007 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0007 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0007 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0007 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0007 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0007 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0007 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0007 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0007 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0007 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0007 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0007 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0007 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0007 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0007 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0007 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0007 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0007 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0007 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0007 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0007 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0007 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0007 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0007 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0007 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0007 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0007 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0007 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0007 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0007 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0007 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0007 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0007 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0007 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0007 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0007 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0007 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0007 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0007 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0007 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0007 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0007 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0007 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0007 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0007 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0007 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0007 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0007 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0007 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0007 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0007 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0007 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0007 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0007 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0007 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0007 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0007 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0007 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0007 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0007 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0007 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0007 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0007 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0007 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0007 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0007 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0007 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0007 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0007 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0007 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0007 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0007 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0007 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0007 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0007 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0007 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0007 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0007 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0007 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0007 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0007 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0007 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0007 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0007 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0007 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0007 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0007 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0007 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0007 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0007 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0007 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0007 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0007 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0007 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0007 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0007 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0007 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0007 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0007 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0007 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0007 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0007 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0007 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0007 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0007 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0007 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0007 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0007 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0007 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0007 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0007 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0007 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0007 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0007 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0007 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0007 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0007 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0007 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0007 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0007 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0007 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0007 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0007 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0007 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0007 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0007 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0007 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0007 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0007 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0007 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0007 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0007 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0007 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0007 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0007 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0007 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0007 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0007 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0007 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0007 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0007 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0007 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0007 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0007 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0007 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0007 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0007 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0007 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0007 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0007 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0007 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0007 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0007 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0007 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0007 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0007 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0007 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0007 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0007 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0007 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0007 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0007 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0007 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0007 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0007 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0007 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0007 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0007 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0007 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0007 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0007 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0007 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0007 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0007 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0007 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0007 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0007 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0007 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0007 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0007 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0007 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0007 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0007 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0007 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0007 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0007 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0007 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0007 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0007 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0007 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0007 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0007 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0007 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0007 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0007 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0007 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0007 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0007 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0007 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0007 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0007 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0007 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0007 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0007 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0007 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0007 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0007 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0007 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0007 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0007 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0007 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0007 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0007 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0007 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0007 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0007 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0007 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0007 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0007 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0007 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0007 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0007 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0007 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0007 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0007 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0007 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0007 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0007 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0007 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0007 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0007 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0007 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0007 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0007 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0007 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0007 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0007 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0007 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0007 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0007 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0007 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0007 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0007 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0007 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0007 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0007 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0007 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0007 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0007 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0007 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0007 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0007 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0007 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0007 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0007 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0007 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0007 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0007 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0007 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0007 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0007 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0007 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0007 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0007 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0007 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0007 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0007 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0007 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0007 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0007 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0007 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0007 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0007 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0007 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0007 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0007 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0007 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0007 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0007 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0007 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0007 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0007 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0007 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0007 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0007 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0007 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0007 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0007 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0007 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0007 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0007 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0007 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0007 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0007 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0007 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0007 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0007 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0007 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0007 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0007 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0007 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0007 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0007 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0007 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0007 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0007 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0007 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0007 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0007 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0007 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0007 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0007 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0007 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0007 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0007 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0007 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0007 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0007 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0007 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0007 7.9623e-08 0)
L_S2_12|A1 G1_1_OUT _S2_12|A1  2.067833848e-12
L_S2_12|A2 _S2_12|A1 _S2_12|A2  4.135667696e-12
L_S2_12|A3 _S2_12|A3 _S2_12|AB  8.271335392e-12
L_S2_12|B1 P2_1_OUT _S2_12|B1  2.067833848e-12
L_S2_12|B2 _S2_12|B1 _S2_12|B2  4.135667696e-12
L_S2_12|B3 _S2_12|B3 _S2_12|AB  8.271335392e-12
L_S2_12|T1 T22 _S2_12|T1  2.067833848e-12
L_S2_12|T2 _S2_12|T1 _S2_12|T2  4.135667696e-12
L_S2_12|Q2 _S2_12|ABTQ _S2_12|Q1  4.135667696e-12
L_S2_12|Q1 _S2_12|Q1 S2_2_TX  2.067833848e-12
IT23|T 0 T23  PWL(0 0 1.7e-11 0 2e-11 0.0028 2.3e-11 0 2.17e-10 0 2.2e-10 0.0028 2.23e-10 0 4.17e-10 0 4.2e-10 0.0028 4.23e-10 0 6.17e-10 0 6.2e-10 0.0028 6.23e-10 0 8.17e-10 0 8.2e-10 0.0028 8.23e-10 0 1.017e-09 0 1.02e-09 0.0028 1.023e-09 0 1.217e-09 0 1.22e-09 0.0028 1.223e-09 0 1.417e-09 0 1.42e-09 0.0028 1.423e-09 0 1.617e-09 0 1.62e-09 0.0028 1.623e-09 0 1.817e-09 0 1.82e-09 0.0028 1.823e-09 0 2.017e-09 0 2.02e-09 0.0028 2.023e-09 0 2.217e-09 0 2.22e-09 0.0028 2.223e-09 0 2.417e-09 0 2.42e-09 0.0028 2.423e-09 0 2.617e-09 0 2.62e-09 0.0028 2.623e-09 0 2.817e-09 0 2.82e-09 0.0028 2.823e-09 0 3.017e-09 0 3.02e-09 0.0028 3.023e-09 0 3.217e-09 0 3.22e-09 0.0028 3.223e-09 0 3.417e-09 0 3.42e-09 0.0028 3.423e-09 0 3.617e-09 0 3.62e-09 0.0028 3.623e-09 0 3.817e-09 0 3.82e-09 0.0028 3.823e-09 0 4.017e-09 0 4.02e-09 0.0028 4.023e-09 0 4.217e-09 0 4.22e-09 0.0028 4.223e-09 0 4.417e-09 0 4.42e-09 0.0028 4.423e-09 0 4.617e-09 0 4.62e-09 0.0028 4.623e-09 0 4.817e-09 0 4.82e-09 0.0028 4.823e-09 0 5.017e-09 0 5.02e-09 0.0028 5.023e-09 0 5.217e-09 0 5.22e-09 0.0028 5.223e-09 0 5.417e-09 0 5.42e-09 0.0028 5.423e-09 0 5.617e-09 0 5.62e-09 0.0028 5.623e-09 0 5.817e-09 0 5.82e-09 0.0028 5.823e-09 0 6.017e-09 0 6.02e-09 0.0028 6.023e-09 0 6.217e-09 0 6.22e-09 0.0028 6.223e-09 0 6.417e-09 0 6.42e-09 0.0028 6.423e-09 0 6.617e-09 0 6.62e-09 0.0028 6.623e-09 0 6.817e-09 0 6.82e-09 0.0028 6.823e-09 0 7.017e-09 0 7.02e-09 0.0028 7.023e-09 0 7.217e-09 0 7.22e-09 0.0028 7.223e-09 0 7.417e-09 0 7.42e-09 0.0028 7.423e-09 0 7.617e-09 0 7.62e-09 0.0028 7.623e-09 0 7.817e-09 0 7.82e-09 0.0028 7.823e-09 0 8.017e-09 0 8.02e-09 0.0028 8.023e-09 0 8.217e-09 0 8.22e-09 0.0028 8.223e-09 0 8.417e-09 0 8.42e-09 0.0028 8.423e-09 0 8.617e-09 0 8.62e-09 0.0028 8.623e-09 0 8.817e-09 0 8.82e-09 0.0028 8.823e-09 0 9.017e-09 0 9.02e-09 0.0028 9.023e-09 0 9.217e-09 0 9.22e-09 0.0028 9.223e-09 0 9.417e-09 0 9.42e-09 0.0028 9.423e-09 0 9.617e-09 0 9.62e-09 0.0028 9.623e-09 0 9.817e-09 0 9.82e-09 0.0028 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0028 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0028 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0028 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0028 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0028 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0028 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0028 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0028 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0028 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0028 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0028 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0028 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0028 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0028 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0028 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0028 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0028 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0028 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0028 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0028 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0028 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0028 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0028 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0028 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0028 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0028 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0028 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0028 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0028 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0028 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0028 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0028 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0028 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0028 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0028 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0028 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0028 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0028 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0028 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0028 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0028 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0028 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0028 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0028 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0028 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0028 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0028 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0028 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0028 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0028 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0028 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0028 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0028 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0028 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0028 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0028 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0028 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0028 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0028 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0028 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0028 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0028 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0028 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0028 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0028 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0028 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0028 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0028 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0028 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0028 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0028 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0028 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0028 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0028 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0028 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0028 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0028 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0028 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0028 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0028 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0028 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0028 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0028 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0028 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0028 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0028 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0028 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0028 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0028 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0028 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0028 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0028 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0028 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0028 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0028 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0028 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0028 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0028 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0028 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0028 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0028 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0028 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0028 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0028 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0028 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0028 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0028 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0028 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0028 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0028 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0028 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0028 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0028 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0028 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0028 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0028 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0028 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0028 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0028 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0028 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0028 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0028 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0028 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0028 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0028 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0028 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0028 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0028 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0028 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0028 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0028 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0028 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0028 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0028 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0028 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0028 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0028 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0028 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0028 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0028 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0028 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0028 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0028 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0028 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0028 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0028 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0028 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0028 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0028 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0028 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0028 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0028 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0028 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0028 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0028 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0028 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0028 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0028 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0028 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0028 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0028 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0028 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0028 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0028 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0028 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0028 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0028 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0028 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0028 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0028 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0028 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0028 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0028 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0028 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0028 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0028 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0028 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0028 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0028 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0028 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0028 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0028 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0028 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0028 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0028 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0028 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0028 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0028 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0028 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0028 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0028 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0028 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0028 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0028 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0028 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0028 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0028 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0028 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0028 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0028 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0028 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0028 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0028 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0028 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0028 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0028 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0028 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0028 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0028 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0028 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0028 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0028 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0028 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0028 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0028 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0028 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0028 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0028 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0028 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0028 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0028 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0028 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0028 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0028 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0028 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0028 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0028 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0028 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0028 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0028 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0028 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0028 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0028 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0028 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0028 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0028 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0028 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0028 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0028 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0028 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0028 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0028 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0028 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0028 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0028 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0028 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0028 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0028 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0028 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0028 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0028 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0028 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0028 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0028 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0028 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0028 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0028 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0028 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0028 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0028 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0028 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0028 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0028 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0028 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0028 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0028 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0028 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0028 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0028 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0028 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0028 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0028 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0028 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0028 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0028 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0028 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0028 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0028 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0028 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0028 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0028 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0028 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0028 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0028 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0028 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0028 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0028 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0028 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0028 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0028 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0028 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0028 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0028 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0028 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0028 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0028 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0028 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0028 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0028 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0028 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0028 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0028 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0028 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0028 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0028 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0028 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0028 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0028 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0028 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0028 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0028 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0028 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0028 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0028 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0028 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0028 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0028 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0028 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0028 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0028 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0028 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0028 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0028 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0028 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0028 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0028 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0028 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0028 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0028 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0028 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0028 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0028 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0028 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0028 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0028 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0028 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0028 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0028 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0028 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0028 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0028 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0028 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0028 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0028 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0028 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0028 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0028 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0028 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0028 7.9623e-08 0)
IT24|T 0 T24  PWL(0 0 1.7e-11 0 2e-11 0.0028 2.3e-11 0 2.17e-10 0 2.2e-10 0.0028 2.23e-10 0 4.17e-10 0 4.2e-10 0.0028 4.23e-10 0 6.17e-10 0 6.2e-10 0.0028 6.23e-10 0 8.17e-10 0 8.2e-10 0.0028 8.23e-10 0 1.017e-09 0 1.02e-09 0.0028 1.023e-09 0 1.217e-09 0 1.22e-09 0.0028 1.223e-09 0 1.417e-09 0 1.42e-09 0.0028 1.423e-09 0 1.617e-09 0 1.62e-09 0.0028 1.623e-09 0 1.817e-09 0 1.82e-09 0.0028 1.823e-09 0 2.017e-09 0 2.02e-09 0.0028 2.023e-09 0 2.217e-09 0 2.22e-09 0.0028 2.223e-09 0 2.417e-09 0 2.42e-09 0.0028 2.423e-09 0 2.617e-09 0 2.62e-09 0.0028 2.623e-09 0 2.817e-09 0 2.82e-09 0.0028 2.823e-09 0 3.017e-09 0 3.02e-09 0.0028 3.023e-09 0 3.217e-09 0 3.22e-09 0.0028 3.223e-09 0 3.417e-09 0 3.42e-09 0.0028 3.423e-09 0 3.617e-09 0 3.62e-09 0.0028 3.623e-09 0 3.817e-09 0 3.82e-09 0.0028 3.823e-09 0 4.017e-09 0 4.02e-09 0.0028 4.023e-09 0 4.217e-09 0 4.22e-09 0.0028 4.223e-09 0 4.417e-09 0 4.42e-09 0.0028 4.423e-09 0 4.617e-09 0 4.62e-09 0.0028 4.623e-09 0 4.817e-09 0 4.82e-09 0.0028 4.823e-09 0 5.017e-09 0 5.02e-09 0.0028 5.023e-09 0 5.217e-09 0 5.22e-09 0.0028 5.223e-09 0 5.417e-09 0 5.42e-09 0.0028 5.423e-09 0 5.617e-09 0 5.62e-09 0.0028 5.623e-09 0 5.817e-09 0 5.82e-09 0.0028 5.823e-09 0 6.017e-09 0 6.02e-09 0.0028 6.023e-09 0 6.217e-09 0 6.22e-09 0.0028 6.223e-09 0 6.417e-09 0 6.42e-09 0.0028 6.423e-09 0 6.617e-09 0 6.62e-09 0.0028 6.623e-09 0 6.817e-09 0 6.82e-09 0.0028 6.823e-09 0 7.017e-09 0 7.02e-09 0.0028 7.023e-09 0 7.217e-09 0 7.22e-09 0.0028 7.223e-09 0 7.417e-09 0 7.42e-09 0.0028 7.423e-09 0 7.617e-09 0 7.62e-09 0.0028 7.623e-09 0 7.817e-09 0 7.82e-09 0.0028 7.823e-09 0 8.017e-09 0 8.02e-09 0.0028 8.023e-09 0 8.217e-09 0 8.22e-09 0.0028 8.223e-09 0 8.417e-09 0 8.42e-09 0.0028 8.423e-09 0 8.617e-09 0 8.62e-09 0.0028 8.623e-09 0 8.817e-09 0 8.82e-09 0.0028 8.823e-09 0 9.017e-09 0 9.02e-09 0.0028 9.023e-09 0 9.217e-09 0 9.22e-09 0.0028 9.223e-09 0 9.417e-09 0 9.42e-09 0.0028 9.423e-09 0 9.617e-09 0 9.62e-09 0.0028 9.623e-09 0 9.817e-09 0 9.82e-09 0.0028 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0028 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0028 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0028 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0028 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0028 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0028 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0028 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0028 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0028 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0028 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0028 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0028 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0028 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0028 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0028 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0028 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0028 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0028 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0028 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0028 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0028 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0028 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0028 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0028 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0028 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0028 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0028 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0028 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0028 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0028 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0028 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0028 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0028 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0028 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0028 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0028 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0028 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0028 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0028 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0028 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0028 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0028 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0028 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0028 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0028 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0028 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0028 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0028 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0028 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0028 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0028 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0028 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0028 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0028 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0028 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0028 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0028 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0028 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0028 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0028 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0028 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0028 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0028 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0028 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0028 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0028 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0028 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0028 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0028 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0028 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0028 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0028 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0028 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0028 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0028 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0028 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0028 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0028 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0028 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0028 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0028 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0028 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0028 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0028 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0028 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0028 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0028 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0028 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0028 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0028 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0028 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0028 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0028 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0028 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0028 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0028 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0028 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0028 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0028 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0028 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0028 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0028 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0028 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0028 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0028 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0028 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0028 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0028 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0028 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0028 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0028 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0028 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0028 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0028 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0028 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0028 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0028 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0028 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0028 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0028 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0028 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0028 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0028 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0028 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0028 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0028 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0028 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0028 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0028 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0028 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0028 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0028 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0028 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0028 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0028 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0028 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0028 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0028 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0028 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0028 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0028 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0028 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0028 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0028 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0028 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0028 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0028 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0028 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0028 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0028 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0028 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0028 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0028 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0028 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0028 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0028 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0028 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0028 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0028 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0028 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0028 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0028 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0028 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0028 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0028 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0028 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0028 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0028 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0028 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0028 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0028 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0028 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0028 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0028 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0028 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0028 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0028 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0028 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0028 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0028 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0028 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0028 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0028 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0028 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0028 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0028 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0028 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0028 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0028 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0028 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0028 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0028 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0028 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0028 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0028 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0028 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0028 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0028 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0028 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0028 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0028 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0028 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0028 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0028 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0028 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0028 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0028 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0028 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0028 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0028 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0028 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0028 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0028 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0028 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0028 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0028 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0028 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0028 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0028 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0028 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0028 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0028 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0028 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0028 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0028 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0028 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0028 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0028 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0028 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0028 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0028 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0028 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0028 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0028 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0028 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0028 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0028 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0028 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0028 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0028 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0028 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0028 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0028 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0028 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0028 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0028 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0028 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0028 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0028 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0028 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0028 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0028 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0028 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0028 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0028 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0028 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0028 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0028 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0028 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0028 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0028 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0028 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0028 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0028 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0028 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0028 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0028 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0028 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0028 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0028 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0028 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0028 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0028 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0028 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0028 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0028 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0028 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0028 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0028 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0028 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0028 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0028 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0028 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0028 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0028 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0028 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0028 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0028 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0028 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0028 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0028 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0028 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0028 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0028 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0028 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0028 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0028 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0028 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0028 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0028 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0028 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0028 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0028 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0028 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0028 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0028 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0028 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0028 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0028 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0028 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0028 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0028 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0028 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0028 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0028 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0028 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0028 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0028 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0028 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0028 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0028 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0028 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0028 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0028 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0028 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0028 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0028 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0028 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0028 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0028 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0028 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0028 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0028 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0028 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0028 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0028 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0028 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0028 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0028 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0028 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0028 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0028 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0028 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0028 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0028 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0028 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0028 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0028 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0028 7.9623e-08 0)
IT25|T 0 T25  PWL(0 0 1.7e-11 0 2e-11 0.0014 2.3e-11 0 2.17e-10 0 2.2e-10 0.0014 2.23e-10 0 4.17e-10 0 4.2e-10 0.0014 4.23e-10 0 6.17e-10 0 6.2e-10 0.0014 6.23e-10 0 8.17e-10 0 8.2e-10 0.0014 8.23e-10 0 1.017e-09 0 1.02e-09 0.0014 1.023e-09 0 1.217e-09 0 1.22e-09 0.0014 1.223e-09 0 1.417e-09 0 1.42e-09 0.0014 1.423e-09 0 1.617e-09 0 1.62e-09 0.0014 1.623e-09 0 1.817e-09 0 1.82e-09 0.0014 1.823e-09 0 2.017e-09 0 2.02e-09 0.0014 2.023e-09 0 2.217e-09 0 2.22e-09 0.0014 2.223e-09 0 2.417e-09 0 2.42e-09 0.0014 2.423e-09 0 2.617e-09 0 2.62e-09 0.0014 2.623e-09 0 2.817e-09 0 2.82e-09 0.0014 2.823e-09 0 3.017e-09 0 3.02e-09 0.0014 3.023e-09 0 3.217e-09 0 3.22e-09 0.0014 3.223e-09 0 3.417e-09 0 3.42e-09 0.0014 3.423e-09 0 3.617e-09 0 3.62e-09 0.0014 3.623e-09 0 3.817e-09 0 3.82e-09 0.0014 3.823e-09 0 4.017e-09 0 4.02e-09 0.0014 4.023e-09 0 4.217e-09 0 4.22e-09 0.0014 4.223e-09 0 4.417e-09 0 4.42e-09 0.0014 4.423e-09 0 4.617e-09 0 4.62e-09 0.0014 4.623e-09 0 4.817e-09 0 4.82e-09 0.0014 4.823e-09 0 5.017e-09 0 5.02e-09 0.0014 5.023e-09 0 5.217e-09 0 5.22e-09 0.0014 5.223e-09 0 5.417e-09 0 5.42e-09 0.0014 5.423e-09 0 5.617e-09 0 5.62e-09 0.0014 5.623e-09 0 5.817e-09 0 5.82e-09 0.0014 5.823e-09 0 6.017e-09 0 6.02e-09 0.0014 6.023e-09 0 6.217e-09 0 6.22e-09 0.0014 6.223e-09 0 6.417e-09 0 6.42e-09 0.0014 6.423e-09 0 6.617e-09 0 6.62e-09 0.0014 6.623e-09 0 6.817e-09 0 6.82e-09 0.0014 6.823e-09 0 7.017e-09 0 7.02e-09 0.0014 7.023e-09 0 7.217e-09 0 7.22e-09 0.0014 7.223e-09 0 7.417e-09 0 7.42e-09 0.0014 7.423e-09 0 7.617e-09 0 7.62e-09 0.0014 7.623e-09 0 7.817e-09 0 7.82e-09 0.0014 7.823e-09 0 8.017e-09 0 8.02e-09 0.0014 8.023e-09 0 8.217e-09 0 8.22e-09 0.0014 8.223e-09 0 8.417e-09 0 8.42e-09 0.0014 8.423e-09 0 8.617e-09 0 8.62e-09 0.0014 8.623e-09 0 8.817e-09 0 8.82e-09 0.0014 8.823e-09 0 9.017e-09 0 9.02e-09 0.0014 9.023e-09 0 9.217e-09 0 9.22e-09 0.0014 9.223e-09 0 9.417e-09 0 9.42e-09 0.0014 9.423e-09 0 9.617e-09 0 9.62e-09 0.0014 9.623e-09 0 9.817e-09 0 9.82e-09 0.0014 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0014 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0014 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0014 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0014 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0014 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0014 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0014 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0014 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0014 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0014 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0014 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0014 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0014 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0014 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0014 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0014 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0014 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0014 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0014 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0014 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0014 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0014 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0014 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0014 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0014 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0014 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0014 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0014 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0014 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0014 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0014 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0014 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0014 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0014 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0014 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0014 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0014 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0014 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0014 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0014 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0014 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0014 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0014 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0014 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0014 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0014 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0014 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0014 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0014 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0014 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0014 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0014 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0014 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0014 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0014 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0014 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0014 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0014 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0014 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0014 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0014 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0014 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0014 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0014 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0014 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0014 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0014 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0014 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0014 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0014 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0014 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0014 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0014 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0014 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0014 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0014 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0014 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0014 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0014 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0014 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0014 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0014 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0014 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0014 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0014 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0014 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0014 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0014 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0014 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0014 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0014 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0014 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0014 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0014 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0014 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0014 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0014 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0014 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0014 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0014 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0014 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0014 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0014 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0014 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0014 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0014 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0014 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0014 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0014 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0014 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0014 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0014 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0014 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0014 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0014 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0014 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0014 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0014 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0014 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0014 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0014 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0014 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0014 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0014 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0014 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0014 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0014 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0014 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0014 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0014 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0014 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0014 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0014 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0014 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0014 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0014 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0014 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0014 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0014 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0014 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0014 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0014 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0014 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0014 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0014 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0014 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0014 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0014 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0014 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0014 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0014 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0014 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0014 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0014 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0014 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0014 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0014 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0014 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0014 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0014 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0014 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0014 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0014 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0014 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0014 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0014 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0014 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0014 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0014 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0014 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0014 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0014 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0014 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0014 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0014 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0014 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0014 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0014 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0014 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0014 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0014 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0014 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0014 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0014 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0014 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0014 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0014 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0014 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0014 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0014 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0014 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0014 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0014 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0014 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0014 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0014 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0014 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0014 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0014 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0014 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0014 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0014 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0014 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0014 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0014 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0014 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0014 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0014 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0014 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0014 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0014 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0014 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0014 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0014 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0014 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0014 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0014 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0014 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0014 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0014 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0014 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0014 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0014 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0014 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0014 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0014 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0014 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0014 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0014 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0014 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0014 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0014 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0014 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0014 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0014 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0014 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0014 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0014 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0014 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0014 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0014 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0014 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0014 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0014 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0014 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0014 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0014 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0014 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0014 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0014 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0014 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0014 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0014 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0014 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0014 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0014 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0014 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0014 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0014 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0014 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0014 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0014 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0014 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0014 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0014 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0014 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0014 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0014 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0014 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0014 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0014 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0014 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0014 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0014 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0014 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0014 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0014 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0014 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0014 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0014 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0014 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0014 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0014 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0014 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0014 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0014 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0014 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0014 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0014 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0014 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0014 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0014 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0014 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0014 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0014 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0014 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0014 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0014 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0014 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0014 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0014 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0014 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0014 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0014 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0014 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0014 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0014 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0014 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0014 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0014 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0014 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0014 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0014 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0014 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0014 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0014 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0014 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0014 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0014 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0014 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0014 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0014 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0014 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0014 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0014 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0014 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0014 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0014 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0014 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0014 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0014 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0014 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0014 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0014 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0014 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0014 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0014 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0014 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0014 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0014 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0014 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0014 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0014 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0014 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0014 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0014 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0014 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0014 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0014 7.9623e-08 0)
IT26|T 0 T26  PWL(0 0 1.7e-11 0 2e-11 0.0014 2.3e-11 0 2.17e-10 0 2.2e-10 0.0014 2.23e-10 0 4.17e-10 0 4.2e-10 0.0014 4.23e-10 0 6.17e-10 0 6.2e-10 0.0014 6.23e-10 0 8.17e-10 0 8.2e-10 0.0014 8.23e-10 0 1.017e-09 0 1.02e-09 0.0014 1.023e-09 0 1.217e-09 0 1.22e-09 0.0014 1.223e-09 0 1.417e-09 0 1.42e-09 0.0014 1.423e-09 0 1.617e-09 0 1.62e-09 0.0014 1.623e-09 0 1.817e-09 0 1.82e-09 0.0014 1.823e-09 0 2.017e-09 0 2.02e-09 0.0014 2.023e-09 0 2.217e-09 0 2.22e-09 0.0014 2.223e-09 0 2.417e-09 0 2.42e-09 0.0014 2.423e-09 0 2.617e-09 0 2.62e-09 0.0014 2.623e-09 0 2.817e-09 0 2.82e-09 0.0014 2.823e-09 0 3.017e-09 0 3.02e-09 0.0014 3.023e-09 0 3.217e-09 0 3.22e-09 0.0014 3.223e-09 0 3.417e-09 0 3.42e-09 0.0014 3.423e-09 0 3.617e-09 0 3.62e-09 0.0014 3.623e-09 0 3.817e-09 0 3.82e-09 0.0014 3.823e-09 0 4.017e-09 0 4.02e-09 0.0014 4.023e-09 0 4.217e-09 0 4.22e-09 0.0014 4.223e-09 0 4.417e-09 0 4.42e-09 0.0014 4.423e-09 0 4.617e-09 0 4.62e-09 0.0014 4.623e-09 0 4.817e-09 0 4.82e-09 0.0014 4.823e-09 0 5.017e-09 0 5.02e-09 0.0014 5.023e-09 0 5.217e-09 0 5.22e-09 0.0014 5.223e-09 0 5.417e-09 0 5.42e-09 0.0014 5.423e-09 0 5.617e-09 0 5.62e-09 0.0014 5.623e-09 0 5.817e-09 0 5.82e-09 0.0014 5.823e-09 0 6.017e-09 0 6.02e-09 0.0014 6.023e-09 0 6.217e-09 0 6.22e-09 0.0014 6.223e-09 0 6.417e-09 0 6.42e-09 0.0014 6.423e-09 0 6.617e-09 0 6.62e-09 0.0014 6.623e-09 0 6.817e-09 0 6.82e-09 0.0014 6.823e-09 0 7.017e-09 0 7.02e-09 0.0014 7.023e-09 0 7.217e-09 0 7.22e-09 0.0014 7.223e-09 0 7.417e-09 0 7.42e-09 0.0014 7.423e-09 0 7.617e-09 0 7.62e-09 0.0014 7.623e-09 0 7.817e-09 0 7.82e-09 0.0014 7.823e-09 0 8.017e-09 0 8.02e-09 0.0014 8.023e-09 0 8.217e-09 0 8.22e-09 0.0014 8.223e-09 0 8.417e-09 0 8.42e-09 0.0014 8.423e-09 0 8.617e-09 0 8.62e-09 0.0014 8.623e-09 0 8.817e-09 0 8.82e-09 0.0014 8.823e-09 0 9.017e-09 0 9.02e-09 0.0014 9.023e-09 0 9.217e-09 0 9.22e-09 0.0014 9.223e-09 0 9.417e-09 0 9.42e-09 0.0014 9.423e-09 0 9.617e-09 0 9.62e-09 0.0014 9.623e-09 0 9.817e-09 0 9.82e-09 0.0014 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0014 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0014 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0014 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0014 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0014 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0014 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0014 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0014 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0014 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0014 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0014 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0014 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0014 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0014 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0014 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0014 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0014 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0014 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0014 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0014 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0014 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0014 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0014 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0014 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0014 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0014 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0014 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0014 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0014 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0014 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0014 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0014 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0014 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0014 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0014 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0014 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0014 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0014 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0014 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0014 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0014 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0014 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0014 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0014 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0014 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0014 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0014 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0014 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0014 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0014 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0014 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0014 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0014 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0014 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0014 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0014 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0014 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0014 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0014 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0014 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0014 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0014 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0014 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0014 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0014 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0014 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0014 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0014 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0014 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0014 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0014 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0014 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0014 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0014 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0014 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0014 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0014 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0014 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0014 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0014 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0014 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0014 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0014 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0014 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0014 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0014 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0014 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0014 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0014 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0014 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0014 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0014 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0014 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0014 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0014 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0014 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0014 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0014 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0014 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0014 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0014 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0014 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0014 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0014 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0014 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0014 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0014 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0014 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0014 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0014 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0014 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0014 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0014 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0014 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0014 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0014 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0014 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0014 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0014 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0014 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0014 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0014 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0014 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0014 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0014 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0014 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0014 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0014 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0014 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0014 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0014 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0014 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0014 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0014 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0014 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0014 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0014 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0014 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0014 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0014 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0014 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0014 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0014 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0014 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0014 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0014 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0014 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0014 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0014 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0014 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0014 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0014 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0014 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0014 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0014 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0014 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0014 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0014 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0014 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0014 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0014 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0014 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0014 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0014 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0014 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0014 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0014 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0014 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0014 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0014 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0014 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0014 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0014 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0014 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0014 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0014 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0014 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0014 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0014 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0014 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0014 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0014 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0014 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0014 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0014 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0014 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0014 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0014 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0014 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0014 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0014 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0014 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0014 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0014 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0014 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0014 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0014 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0014 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0014 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0014 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0014 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0014 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0014 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0014 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0014 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0014 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0014 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0014 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0014 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0014 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0014 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0014 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0014 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0014 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0014 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0014 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0014 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0014 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0014 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0014 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0014 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0014 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0014 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0014 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0014 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0014 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0014 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0014 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0014 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0014 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0014 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0014 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0014 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0014 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0014 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0014 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0014 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0014 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0014 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0014 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0014 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0014 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0014 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0014 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0014 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0014 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0014 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0014 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0014 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0014 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0014 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0014 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0014 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0014 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0014 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0014 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0014 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0014 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0014 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0014 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0014 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0014 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0014 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0014 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0014 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0014 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0014 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0014 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0014 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0014 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0014 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0014 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0014 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0014 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0014 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0014 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0014 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0014 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0014 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0014 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0014 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0014 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0014 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0014 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0014 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0014 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0014 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0014 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0014 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0014 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0014 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0014 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0014 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0014 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0014 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0014 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0014 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0014 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0014 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0014 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0014 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0014 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0014 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0014 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0014 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0014 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0014 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0014 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0014 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0014 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0014 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0014 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0014 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0014 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0014 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0014 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0014 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0014 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0014 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0014 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0014 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0014 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0014 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0014 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0014 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0014 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0014 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0014 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0014 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0014 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0014 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0014 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0014 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0014 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0014 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0014 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0014 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0014 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0014 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0014 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0014 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0014 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0014 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0014 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0014 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0014 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0014 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0014 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0014 7.9623e-08 0)
IT27|T 0 T27  PWL(0 0 1.7e-11 0 2e-11 0.0014 2.3e-11 0 2.17e-10 0 2.2e-10 0.0014 2.23e-10 0 4.17e-10 0 4.2e-10 0.0014 4.23e-10 0 6.17e-10 0 6.2e-10 0.0014 6.23e-10 0 8.17e-10 0 8.2e-10 0.0014 8.23e-10 0 1.017e-09 0 1.02e-09 0.0014 1.023e-09 0 1.217e-09 0 1.22e-09 0.0014 1.223e-09 0 1.417e-09 0 1.42e-09 0.0014 1.423e-09 0 1.617e-09 0 1.62e-09 0.0014 1.623e-09 0 1.817e-09 0 1.82e-09 0.0014 1.823e-09 0 2.017e-09 0 2.02e-09 0.0014 2.023e-09 0 2.217e-09 0 2.22e-09 0.0014 2.223e-09 0 2.417e-09 0 2.42e-09 0.0014 2.423e-09 0 2.617e-09 0 2.62e-09 0.0014 2.623e-09 0 2.817e-09 0 2.82e-09 0.0014 2.823e-09 0 3.017e-09 0 3.02e-09 0.0014 3.023e-09 0 3.217e-09 0 3.22e-09 0.0014 3.223e-09 0 3.417e-09 0 3.42e-09 0.0014 3.423e-09 0 3.617e-09 0 3.62e-09 0.0014 3.623e-09 0 3.817e-09 0 3.82e-09 0.0014 3.823e-09 0 4.017e-09 0 4.02e-09 0.0014 4.023e-09 0 4.217e-09 0 4.22e-09 0.0014 4.223e-09 0 4.417e-09 0 4.42e-09 0.0014 4.423e-09 0 4.617e-09 0 4.62e-09 0.0014 4.623e-09 0 4.817e-09 0 4.82e-09 0.0014 4.823e-09 0 5.017e-09 0 5.02e-09 0.0014 5.023e-09 0 5.217e-09 0 5.22e-09 0.0014 5.223e-09 0 5.417e-09 0 5.42e-09 0.0014 5.423e-09 0 5.617e-09 0 5.62e-09 0.0014 5.623e-09 0 5.817e-09 0 5.82e-09 0.0014 5.823e-09 0 6.017e-09 0 6.02e-09 0.0014 6.023e-09 0 6.217e-09 0 6.22e-09 0.0014 6.223e-09 0 6.417e-09 0 6.42e-09 0.0014 6.423e-09 0 6.617e-09 0 6.62e-09 0.0014 6.623e-09 0 6.817e-09 0 6.82e-09 0.0014 6.823e-09 0 7.017e-09 0 7.02e-09 0.0014 7.023e-09 0 7.217e-09 0 7.22e-09 0.0014 7.223e-09 0 7.417e-09 0 7.42e-09 0.0014 7.423e-09 0 7.617e-09 0 7.62e-09 0.0014 7.623e-09 0 7.817e-09 0 7.82e-09 0.0014 7.823e-09 0 8.017e-09 0 8.02e-09 0.0014 8.023e-09 0 8.217e-09 0 8.22e-09 0.0014 8.223e-09 0 8.417e-09 0 8.42e-09 0.0014 8.423e-09 0 8.617e-09 0 8.62e-09 0.0014 8.623e-09 0 8.817e-09 0 8.82e-09 0.0014 8.823e-09 0 9.017e-09 0 9.02e-09 0.0014 9.023e-09 0 9.217e-09 0 9.22e-09 0.0014 9.223e-09 0 9.417e-09 0 9.42e-09 0.0014 9.423e-09 0 9.617e-09 0 9.62e-09 0.0014 9.623e-09 0 9.817e-09 0 9.82e-09 0.0014 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0014 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0014 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0014 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0014 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0014 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0014 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0014 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0014 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0014 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0014 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0014 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0014 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0014 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0014 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0014 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0014 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0014 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0014 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0014 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0014 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0014 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0014 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0014 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0014 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0014 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0014 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0014 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0014 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0014 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0014 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0014 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0014 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0014 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0014 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0014 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0014 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0014 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0014 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0014 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0014 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0014 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0014 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0014 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0014 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0014 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0014 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0014 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0014 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0014 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0014 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0014 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0014 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0014 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0014 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0014 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0014 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0014 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0014 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0014 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0014 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0014 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0014 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0014 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0014 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0014 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0014 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0014 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0014 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0014 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0014 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0014 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0014 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0014 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0014 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0014 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0014 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0014 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0014 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0014 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0014 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0014 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0014 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0014 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0014 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0014 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0014 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0014 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0014 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0014 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0014 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0014 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0014 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0014 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0014 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0014 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0014 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0014 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0014 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0014 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0014 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0014 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0014 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0014 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0014 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0014 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0014 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0014 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0014 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0014 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0014 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0014 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0014 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0014 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0014 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0014 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0014 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0014 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0014 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0014 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0014 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0014 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0014 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0014 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0014 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0014 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0014 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0014 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0014 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0014 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0014 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0014 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0014 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0014 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0014 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0014 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0014 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0014 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0014 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0014 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0014 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0014 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0014 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0014 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0014 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0014 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0014 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0014 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0014 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0014 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0014 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0014 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0014 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0014 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0014 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0014 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0014 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0014 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0014 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0014 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0014 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0014 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0014 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0014 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0014 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0014 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0014 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0014 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0014 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0014 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0014 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0014 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0014 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0014 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0014 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0014 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0014 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0014 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0014 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0014 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0014 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0014 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0014 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0014 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0014 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0014 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0014 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0014 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0014 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0014 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0014 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0014 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0014 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0014 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0014 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0014 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0014 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0014 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0014 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0014 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0014 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0014 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0014 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0014 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0014 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0014 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0014 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0014 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0014 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0014 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0014 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0014 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0014 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0014 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0014 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0014 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0014 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0014 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0014 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0014 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0014 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0014 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0014 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0014 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0014 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0014 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0014 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0014 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0014 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0014 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0014 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0014 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0014 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0014 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0014 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0014 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0014 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0014 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0014 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0014 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0014 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0014 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0014 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0014 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0014 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0014 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0014 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0014 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0014 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0014 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0014 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0014 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0014 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0014 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0014 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0014 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0014 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0014 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0014 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0014 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0014 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0014 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0014 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0014 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0014 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0014 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0014 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0014 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0014 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0014 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0014 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0014 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0014 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0014 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0014 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0014 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0014 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0014 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0014 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0014 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0014 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0014 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0014 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0014 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0014 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0014 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0014 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0014 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0014 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0014 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0014 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0014 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0014 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0014 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0014 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0014 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0014 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0014 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0014 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0014 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0014 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0014 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0014 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0014 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0014 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0014 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0014 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0014 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0014 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0014 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0014 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0014 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0014 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0014 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0014 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0014 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0014 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0014 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0014 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0014 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0014 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0014 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0014 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0014 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0014 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0014 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0014 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0014 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0014 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0014 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0014 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0014 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0014 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0014 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0014 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0014 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0014 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0014 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0014 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0014 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0014 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0014 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0014 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0014 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0014 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0014 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0014 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0014 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0014 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0014 7.9623e-08 0)
IT28|T 0 T28  PWL(0 0 1.7e-11 0 2e-11 0.0028 2.3e-11 0 2.17e-10 0 2.2e-10 0.0028 2.23e-10 0 4.17e-10 0 4.2e-10 0.0028 4.23e-10 0 6.17e-10 0 6.2e-10 0.0028 6.23e-10 0 8.17e-10 0 8.2e-10 0.0028 8.23e-10 0 1.017e-09 0 1.02e-09 0.0028 1.023e-09 0 1.217e-09 0 1.22e-09 0.0028 1.223e-09 0 1.417e-09 0 1.42e-09 0.0028 1.423e-09 0 1.617e-09 0 1.62e-09 0.0028 1.623e-09 0 1.817e-09 0 1.82e-09 0.0028 1.823e-09 0 2.017e-09 0 2.02e-09 0.0028 2.023e-09 0 2.217e-09 0 2.22e-09 0.0028 2.223e-09 0 2.417e-09 0 2.42e-09 0.0028 2.423e-09 0 2.617e-09 0 2.62e-09 0.0028 2.623e-09 0 2.817e-09 0 2.82e-09 0.0028 2.823e-09 0 3.017e-09 0 3.02e-09 0.0028 3.023e-09 0 3.217e-09 0 3.22e-09 0.0028 3.223e-09 0 3.417e-09 0 3.42e-09 0.0028 3.423e-09 0 3.617e-09 0 3.62e-09 0.0028 3.623e-09 0 3.817e-09 0 3.82e-09 0.0028 3.823e-09 0 4.017e-09 0 4.02e-09 0.0028 4.023e-09 0 4.217e-09 0 4.22e-09 0.0028 4.223e-09 0 4.417e-09 0 4.42e-09 0.0028 4.423e-09 0 4.617e-09 0 4.62e-09 0.0028 4.623e-09 0 4.817e-09 0 4.82e-09 0.0028 4.823e-09 0 5.017e-09 0 5.02e-09 0.0028 5.023e-09 0 5.217e-09 0 5.22e-09 0.0028 5.223e-09 0 5.417e-09 0 5.42e-09 0.0028 5.423e-09 0 5.617e-09 0 5.62e-09 0.0028 5.623e-09 0 5.817e-09 0 5.82e-09 0.0028 5.823e-09 0 6.017e-09 0 6.02e-09 0.0028 6.023e-09 0 6.217e-09 0 6.22e-09 0.0028 6.223e-09 0 6.417e-09 0 6.42e-09 0.0028 6.423e-09 0 6.617e-09 0 6.62e-09 0.0028 6.623e-09 0 6.817e-09 0 6.82e-09 0.0028 6.823e-09 0 7.017e-09 0 7.02e-09 0.0028 7.023e-09 0 7.217e-09 0 7.22e-09 0.0028 7.223e-09 0 7.417e-09 0 7.42e-09 0.0028 7.423e-09 0 7.617e-09 0 7.62e-09 0.0028 7.623e-09 0 7.817e-09 0 7.82e-09 0.0028 7.823e-09 0 8.017e-09 0 8.02e-09 0.0028 8.023e-09 0 8.217e-09 0 8.22e-09 0.0028 8.223e-09 0 8.417e-09 0 8.42e-09 0.0028 8.423e-09 0 8.617e-09 0 8.62e-09 0.0028 8.623e-09 0 8.817e-09 0 8.82e-09 0.0028 8.823e-09 0 9.017e-09 0 9.02e-09 0.0028 9.023e-09 0 9.217e-09 0 9.22e-09 0.0028 9.223e-09 0 9.417e-09 0 9.42e-09 0.0028 9.423e-09 0 9.617e-09 0 9.62e-09 0.0028 9.623e-09 0 9.817e-09 0 9.82e-09 0.0028 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0028 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0028 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0028 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0028 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0028 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0028 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0028 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0028 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0028 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0028 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0028 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0028 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0028 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0028 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0028 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0028 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0028 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0028 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0028 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0028 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0028 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0028 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0028 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0028 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0028 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0028 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0028 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0028 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0028 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0028 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0028 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0028 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0028 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0028 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0028 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0028 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0028 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0028 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0028 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0028 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0028 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0028 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0028 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0028 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0028 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0028 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0028 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0028 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0028 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0028 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0028 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0028 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0028 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0028 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0028 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0028 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0028 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0028 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0028 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0028 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0028 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0028 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0028 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0028 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0028 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0028 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0028 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0028 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0028 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0028 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0028 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0028 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0028 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0028 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0028 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0028 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0028 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0028 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0028 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0028 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0028 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0028 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0028 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0028 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0028 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0028 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0028 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0028 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0028 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0028 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0028 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0028 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0028 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0028 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0028 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0028 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0028 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0028 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0028 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0028 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0028 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0028 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0028 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0028 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0028 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0028 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0028 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0028 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0028 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0028 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0028 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0028 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0028 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0028 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0028 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0028 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0028 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0028 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0028 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0028 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0028 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0028 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0028 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0028 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0028 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0028 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0028 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0028 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0028 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0028 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0028 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0028 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0028 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0028 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0028 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0028 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0028 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0028 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0028 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0028 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0028 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0028 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0028 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0028 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0028 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0028 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0028 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0028 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0028 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0028 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0028 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0028 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0028 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0028 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0028 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0028 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0028 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0028 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0028 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0028 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0028 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0028 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0028 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0028 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0028 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0028 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0028 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0028 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0028 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0028 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0028 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0028 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0028 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0028 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0028 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0028 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0028 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0028 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0028 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0028 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0028 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0028 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0028 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0028 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0028 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0028 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0028 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0028 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0028 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0028 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0028 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0028 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0028 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0028 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0028 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0028 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0028 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0028 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0028 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0028 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0028 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0028 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0028 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0028 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0028 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0028 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0028 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0028 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0028 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0028 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0028 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0028 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0028 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0028 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0028 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0028 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0028 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0028 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0028 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0028 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0028 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0028 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0028 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0028 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0028 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0028 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0028 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0028 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0028 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0028 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0028 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0028 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0028 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0028 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0028 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0028 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0028 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0028 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0028 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0028 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0028 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0028 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0028 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0028 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0028 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0028 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0028 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0028 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0028 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0028 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0028 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0028 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0028 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0028 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0028 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0028 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0028 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0028 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0028 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0028 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0028 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0028 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0028 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0028 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0028 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0028 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0028 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0028 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0028 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0028 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0028 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0028 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0028 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0028 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0028 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0028 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0028 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0028 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0028 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0028 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0028 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0028 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0028 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0028 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0028 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0028 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0028 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0028 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0028 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0028 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0028 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0028 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0028 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0028 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0028 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0028 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0028 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0028 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0028 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0028 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0028 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0028 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0028 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0028 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0028 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0028 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0028 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0028 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0028 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0028 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0028 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0028 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0028 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0028 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0028 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0028 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0028 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0028 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0028 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0028 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0028 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0028 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0028 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0028 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0028 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0028 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0028 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0028 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0028 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0028 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0028 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0028 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0028 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0028 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0028 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0028 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0028 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0028 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0028 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0028 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0028 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0028 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0028 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0028 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0028 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0028 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0028 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0028 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0028 7.9623e-08 0)
IT29|T 0 T29  PWL(0 0 1.7e-11 0 2e-11 0.0007 2.3e-11 0 2.17e-10 0 2.2e-10 0.0007 2.23e-10 0 4.17e-10 0 4.2e-10 0.0007 4.23e-10 0 6.17e-10 0 6.2e-10 0.0007 6.23e-10 0 8.17e-10 0 8.2e-10 0.0007 8.23e-10 0 1.017e-09 0 1.02e-09 0.0007 1.023e-09 0 1.217e-09 0 1.22e-09 0.0007 1.223e-09 0 1.417e-09 0 1.42e-09 0.0007 1.423e-09 0 1.617e-09 0 1.62e-09 0.0007 1.623e-09 0 1.817e-09 0 1.82e-09 0.0007 1.823e-09 0 2.017e-09 0 2.02e-09 0.0007 2.023e-09 0 2.217e-09 0 2.22e-09 0.0007 2.223e-09 0 2.417e-09 0 2.42e-09 0.0007 2.423e-09 0 2.617e-09 0 2.62e-09 0.0007 2.623e-09 0 2.817e-09 0 2.82e-09 0.0007 2.823e-09 0 3.017e-09 0 3.02e-09 0.0007 3.023e-09 0 3.217e-09 0 3.22e-09 0.0007 3.223e-09 0 3.417e-09 0 3.42e-09 0.0007 3.423e-09 0 3.617e-09 0 3.62e-09 0.0007 3.623e-09 0 3.817e-09 0 3.82e-09 0.0007 3.823e-09 0 4.017e-09 0 4.02e-09 0.0007 4.023e-09 0 4.217e-09 0 4.22e-09 0.0007 4.223e-09 0 4.417e-09 0 4.42e-09 0.0007 4.423e-09 0 4.617e-09 0 4.62e-09 0.0007 4.623e-09 0 4.817e-09 0 4.82e-09 0.0007 4.823e-09 0 5.017e-09 0 5.02e-09 0.0007 5.023e-09 0 5.217e-09 0 5.22e-09 0.0007 5.223e-09 0 5.417e-09 0 5.42e-09 0.0007 5.423e-09 0 5.617e-09 0 5.62e-09 0.0007 5.623e-09 0 5.817e-09 0 5.82e-09 0.0007 5.823e-09 0 6.017e-09 0 6.02e-09 0.0007 6.023e-09 0 6.217e-09 0 6.22e-09 0.0007 6.223e-09 0 6.417e-09 0 6.42e-09 0.0007 6.423e-09 0 6.617e-09 0 6.62e-09 0.0007 6.623e-09 0 6.817e-09 0 6.82e-09 0.0007 6.823e-09 0 7.017e-09 0 7.02e-09 0.0007 7.023e-09 0 7.217e-09 0 7.22e-09 0.0007 7.223e-09 0 7.417e-09 0 7.42e-09 0.0007 7.423e-09 0 7.617e-09 0 7.62e-09 0.0007 7.623e-09 0 7.817e-09 0 7.82e-09 0.0007 7.823e-09 0 8.017e-09 0 8.02e-09 0.0007 8.023e-09 0 8.217e-09 0 8.22e-09 0.0007 8.223e-09 0 8.417e-09 0 8.42e-09 0.0007 8.423e-09 0 8.617e-09 0 8.62e-09 0.0007 8.623e-09 0 8.817e-09 0 8.82e-09 0.0007 8.823e-09 0 9.017e-09 0 9.02e-09 0.0007 9.023e-09 0 9.217e-09 0 9.22e-09 0.0007 9.223e-09 0 9.417e-09 0 9.42e-09 0.0007 9.423e-09 0 9.617e-09 0 9.62e-09 0.0007 9.623e-09 0 9.817e-09 0 9.82e-09 0.0007 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0007 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0007 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0007 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0007 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0007 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0007 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0007 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0007 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0007 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0007 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0007 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0007 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0007 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0007 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0007 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0007 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0007 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0007 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0007 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0007 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0007 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0007 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0007 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0007 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0007 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0007 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0007 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0007 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0007 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0007 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0007 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0007 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0007 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0007 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0007 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0007 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0007 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0007 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0007 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0007 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0007 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0007 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0007 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0007 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0007 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0007 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0007 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0007 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0007 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0007 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0007 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0007 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0007 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0007 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0007 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0007 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0007 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0007 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0007 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0007 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0007 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0007 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0007 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0007 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0007 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0007 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0007 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0007 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0007 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0007 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0007 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0007 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0007 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0007 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0007 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0007 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0007 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0007 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0007 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0007 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0007 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0007 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0007 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0007 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0007 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0007 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0007 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0007 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0007 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0007 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0007 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0007 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0007 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0007 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0007 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0007 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0007 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0007 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0007 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0007 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0007 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0007 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0007 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0007 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0007 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0007 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0007 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0007 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0007 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0007 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0007 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0007 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0007 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0007 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0007 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0007 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0007 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0007 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0007 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0007 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0007 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0007 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0007 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0007 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0007 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0007 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0007 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0007 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0007 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0007 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0007 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0007 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0007 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0007 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0007 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0007 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0007 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0007 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0007 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0007 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0007 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0007 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0007 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0007 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0007 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0007 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0007 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0007 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0007 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0007 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0007 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0007 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0007 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0007 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0007 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0007 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0007 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0007 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0007 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0007 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0007 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0007 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0007 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0007 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0007 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0007 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0007 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0007 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0007 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0007 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0007 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0007 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0007 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0007 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0007 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0007 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0007 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0007 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0007 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0007 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0007 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0007 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0007 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0007 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0007 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0007 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0007 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0007 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0007 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0007 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0007 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0007 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0007 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0007 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0007 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0007 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0007 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0007 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0007 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0007 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0007 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0007 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0007 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0007 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0007 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0007 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0007 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0007 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0007 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0007 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0007 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0007 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0007 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0007 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0007 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0007 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0007 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0007 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0007 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0007 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0007 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0007 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0007 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0007 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0007 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0007 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0007 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0007 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0007 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0007 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0007 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0007 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0007 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0007 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0007 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0007 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0007 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0007 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0007 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0007 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0007 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0007 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0007 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0007 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0007 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0007 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0007 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0007 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0007 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0007 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0007 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0007 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0007 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0007 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0007 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0007 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0007 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0007 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0007 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0007 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0007 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0007 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0007 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0007 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0007 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0007 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0007 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0007 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0007 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0007 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0007 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0007 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0007 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0007 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0007 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0007 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0007 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0007 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0007 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0007 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0007 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0007 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0007 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0007 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0007 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0007 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0007 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0007 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0007 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0007 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0007 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0007 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0007 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0007 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0007 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0007 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0007 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0007 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0007 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0007 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0007 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0007 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0007 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0007 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0007 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0007 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0007 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0007 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0007 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0007 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0007 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0007 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0007 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0007 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0007 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0007 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0007 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0007 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0007 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0007 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0007 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0007 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0007 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0007 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0007 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0007 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0007 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0007 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0007 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0007 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0007 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0007 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0007 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0007 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0007 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0007 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0007 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0007 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0007 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0007 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0007 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0007 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0007 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0007 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0007 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0007 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0007 7.9623e-08 0)
L_IP3_12|1 IP3_1_OUT _IP3_12|A1  2.067833848e-12
L_IP3_12|2 _IP3_12|A1 _IP3_12|A2  4.135667696e-12
L_IP3_12|3 _IP3_12|A3 _IP3_12|A4  8.271335392e-12
L_IP3_12|T T29 _IP3_12|T1  2.067833848e-12
L_IP3_12|4 _IP3_12|T1 _IP3_12|T2  4.135667696e-12
L_IP3_12|5 _IP3_12|A4 _IP3_12|Q1  4.135667696e-12
L_IP3_12|6 _IP3_12|Q1 IP3_2_OUT_TX  2.067833848e-12
IT2A|T 0 T2A  PWL(0 0 1.7e-11 0 2e-11 0.0007 2.3e-11 0 2.17e-10 0 2.2e-10 0.0007 2.23e-10 0 4.17e-10 0 4.2e-10 0.0007 4.23e-10 0 6.17e-10 0 6.2e-10 0.0007 6.23e-10 0 8.17e-10 0 8.2e-10 0.0007 8.23e-10 0 1.017e-09 0 1.02e-09 0.0007 1.023e-09 0 1.217e-09 0 1.22e-09 0.0007 1.223e-09 0 1.417e-09 0 1.42e-09 0.0007 1.423e-09 0 1.617e-09 0 1.62e-09 0.0007 1.623e-09 0 1.817e-09 0 1.82e-09 0.0007 1.823e-09 0 2.017e-09 0 2.02e-09 0.0007 2.023e-09 0 2.217e-09 0 2.22e-09 0.0007 2.223e-09 0 2.417e-09 0 2.42e-09 0.0007 2.423e-09 0 2.617e-09 0 2.62e-09 0.0007 2.623e-09 0 2.817e-09 0 2.82e-09 0.0007 2.823e-09 0 3.017e-09 0 3.02e-09 0.0007 3.023e-09 0 3.217e-09 0 3.22e-09 0.0007 3.223e-09 0 3.417e-09 0 3.42e-09 0.0007 3.423e-09 0 3.617e-09 0 3.62e-09 0.0007 3.623e-09 0 3.817e-09 0 3.82e-09 0.0007 3.823e-09 0 4.017e-09 0 4.02e-09 0.0007 4.023e-09 0 4.217e-09 0 4.22e-09 0.0007 4.223e-09 0 4.417e-09 0 4.42e-09 0.0007 4.423e-09 0 4.617e-09 0 4.62e-09 0.0007 4.623e-09 0 4.817e-09 0 4.82e-09 0.0007 4.823e-09 0 5.017e-09 0 5.02e-09 0.0007 5.023e-09 0 5.217e-09 0 5.22e-09 0.0007 5.223e-09 0 5.417e-09 0 5.42e-09 0.0007 5.423e-09 0 5.617e-09 0 5.62e-09 0.0007 5.623e-09 0 5.817e-09 0 5.82e-09 0.0007 5.823e-09 0 6.017e-09 0 6.02e-09 0.0007 6.023e-09 0 6.217e-09 0 6.22e-09 0.0007 6.223e-09 0 6.417e-09 0 6.42e-09 0.0007 6.423e-09 0 6.617e-09 0 6.62e-09 0.0007 6.623e-09 0 6.817e-09 0 6.82e-09 0.0007 6.823e-09 0 7.017e-09 0 7.02e-09 0.0007 7.023e-09 0 7.217e-09 0 7.22e-09 0.0007 7.223e-09 0 7.417e-09 0 7.42e-09 0.0007 7.423e-09 0 7.617e-09 0 7.62e-09 0.0007 7.623e-09 0 7.817e-09 0 7.82e-09 0.0007 7.823e-09 0 8.017e-09 0 8.02e-09 0.0007 8.023e-09 0 8.217e-09 0 8.22e-09 0.0007 8.223e-09 0 8.417e-09 0 8.42e-09 0.0007 8.423e-09 0 8.617e-09 0 8.62e-09 0.0007 8.623e-09 0 8.817e-09 0 8.82e-09 0.0007 8.823e-09 0 9.017e-09 0 9.02e-09 0.0007 9.023e-09 0 9.217e-09 0 9.22e-09 0.0007 9.223e-09 0 9.417e-09 0 9.42e-09 0.0007 9.423e-09 0 9.617e-09 0 9.62e-09 0.0007 9.623e-09 0 9.817e-09 0 9.82e-09 0.0007 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0007 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0007 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0007 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0007 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0007 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0007 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0007 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0007 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0007 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0007 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0007 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0007 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0007 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0007 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0007 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0007 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0007 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0007 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0007 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0007 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0007 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0007 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0007 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0007 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0007 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0007 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0007 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0007 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0007 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0007 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0007 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0007 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0007 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0007 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0007 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0007 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0007 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0007 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0007 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0007 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0007 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0007 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0007 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0007 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0007 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0007 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0007 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0007 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0007 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0007 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0007 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0007 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0007 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0007 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0007 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0007 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0007 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0007 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0007 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0007 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0007 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0007 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0007 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0007 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0007 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0007 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0007 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0007 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0007 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0007 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0007 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0007 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0007 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0007 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0007 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0007 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0007 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0007 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0007 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0007 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0007 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0007 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0007 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0007 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0007 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0007 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0007 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0007 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0007 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0007 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0007 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0007 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0007 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0007 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0007 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0007 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0007 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0007 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0007 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0007 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0007 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0007 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0007 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0007 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0007 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0007 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0007 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0007 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0007 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0007 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0007 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0007 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0007 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0007 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0007 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0007 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0007 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0007 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0007 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0007 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0007 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0007 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0007 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0007 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0007 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0007 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0007 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0007 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0007 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0007 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0007 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0007 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0007 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0007 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0007 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0007 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0007 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0007 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0007 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0007 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0007 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0007 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0007 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0007 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0007 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0007 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0007 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0007 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0007 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0007 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0007 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0007 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0007 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0007 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0007 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0007 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0007 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0007 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0007 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0007 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0007 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0007 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0007 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0007 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0007 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0007 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0007 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0007 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0007 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0007 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0007 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0007 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0007 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0007 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0007 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0007 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0007 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0007 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0007 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0007 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0007 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0007 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0007 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0007 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0007 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0007 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0007 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0007 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0007 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0007 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0007 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0007 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0007 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0007 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0007 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0007 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0007 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0007 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0007 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0007 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0007 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0007 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0007 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0007 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0007 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0007 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0007 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0007 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0007 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0007 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0007 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0007 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0007 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0007 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0007 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0007 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0007 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0007 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0007 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0007 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0007 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0007 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0007 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0007 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0007 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0007 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0007 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0007 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0007 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0007 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0007 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0007 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0007 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0007 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0007 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0007 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0007 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0007 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0007 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0007 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0007 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0007 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0007 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0007 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0007 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0007 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0007 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0007 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0007 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0007 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0007 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0007 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0007 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0007 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0007 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0007 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0007 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0007 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0007 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0007 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0007 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0007 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0007 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0007 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0007 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0007 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0007 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0007 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0007 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0007 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0007 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0007 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0007 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0007 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0007 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0007 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0007 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0007 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0007 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0007 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0007 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0007 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0007 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0007 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0007 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0007 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0007 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0007 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0007 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0007 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0007 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0007 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0007 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0007 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0007 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0007 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0007 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0007 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0007 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0007 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0007 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0007 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0007 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0007 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0007 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0007 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0007 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0007 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0007 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0007 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0007 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0007 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0007 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0007 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0007 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0007 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0007 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0007 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0007 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0007 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0007 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0007 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0007 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0007 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0007 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0007 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0007 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0007 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0007 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0007 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0007 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0007 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0007 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0007 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0007 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0007 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0007 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0007 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0007 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0007 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0007 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0007 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0007 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0007 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0007 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0007 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0007 7.9623e-08 0)
L_IP5_12|1 IP5_1_OUT _IP5_12|A1  2.067833848e-12
L_IP5_12|2 _IP5_12|A1 _IP5_12|A2  4.135667696e-12
L_IP5_12|3 _IP5_12|A3 _IP5_12|A4  8.271335392e-12
L_IP5_12|T T2A _IP5_12|T1  2.067833848e-12
L_IP5_12|4 _IP5_12|T1 _IP5_12|T2  4.135667696e-12
L_IP5_12|5 _IP5_12|A4 _IP5_12|Q1  4.135667696e-12
L_IP5_12|6 _IP5_12|Q1 IP5_2_OUT_TX  2.067833848e-12
IT2B|T 0 T2B  PWL(0 0 1.7e-11 0 2e-11 0.0007 2.3e-11 0 2.17e-10 0 2.2e-10 0.0007 2.23e-10 0 4.17e-10 0 4.2e-10 0.0007 4.23e-10 0 6.17e-10 0 6.2e-10 0.0007 6.23e-10 0 8.17e-10 0 8.2e-10 0.0007 8.23e-10 0 1.017e-09 0 1.02e-09 0.0007 1.023e-09 0 1.217e-09 0 1.22e-09 0.0007 1.223e-09 0 1.417e-09 0 1.42e-09 0.0007 1.423e-09 0 1.617e-09 0 1.62e-09 0.0007 1.623e-09 0 1.817e-09 0 1.82e-09 0.0007 1.823e-09 0 2.017e-09 0 2.02e-09 0.0007 2.023e-09 0 2.217e-09 0 2.22e-09 0.0007 2.223e-09 0 2.417e-09 0 2.42e-09 0.0007 2.423e-09 0 2.617e-09 0 2.62e-09 0.0007 2.623e-09 0 2.817e-09 0 2.82e-09 0.0007 2.823e-09 0 3.017e-09 0 3.02e-09 0.0007 3.023e-09 0 3.217e-09 0 3.22e-09 0.0007 3.223e-09 0 3.417e-09 0 3.42e-09 0.0007 3.423e-09 0 3.617e-09 0 3.62e-09 0.0007 3.623e-09 0 3.817e-09 0 3.82e-09 0.0007 3.823e-09 0 4.017e-09 0 4.02e-09 0.0007 4.023e-09 0 4.217e-09 0 4.22e-09 0.0007 4.223e-09 0 4.417e-09 0 4.42e-09 0.0007 4.423e-09 0 4.617e-09 0 4.62e-09 0.0007 4.623e-09 0 4.817e-09 0 4.82e-09 0.0007 4.823e-09 0 5.017e-09 0 5.02e-09 0.0007 5.023e-09 0 5.217e-09 0 5.22e-09 0.0007 5.223e-09 0 5.417e-09 0 5.42e-09 0.0007 5.423e-09 0 5.617e-09 0 5.62e-09 0.0007 5.623e-09 0 5.817e-09 0 5.82e-09 0.0007 5.823e-09 0 6.017e-09 0 6.02e-09 0.0007 6.023e-09 0 6.217e-09 0 6.22e-09 0.0007 6.223e-09 0 6.417e-09 0 6.42e-09 0.0007 6.423e-09 0 6.617e-09 0 6.62e-09 0.0007 6.623e-09 0 6.817e-09 0 6.82e-09 0.0007 6.823e-09 0 7.017e-09 0 7.02e-09 0.0007 7.023e-09 0 7.217e-09 0 7.22e-09 0.0007 7.223e-09 0 7.417e-09 0 7.42e-09 0.0007 7.423e-09 0 7.617e-09 0 7.62e-09 0.0007 7.623e-09 0 7.817e-09 0 7.82e-09 0.0007 7.823e-09 0 8.017e-09 0 8.02e-09 0.0007 8.023e-09 0 8.217e-09 0 8.22e-09 0.0007 8.223e-09 0 8.417e-09 0 8.42e-09 0.0007 8.423e-09 0 8.617e-09 0 8.62e-09 0.0007 8.623e-09 0 8.817e-09 0 8.82e-09 0.0007 8.823e-09 0 9.017e-09 0 9.02e-09 0.0007 9.023e-09 0 9.217e-09 0 9.22e-09 0.0007 9.223e-09 0 9.417e-09 0 9.42e-09 0.0007 9.423e-09 0 9.617e-09 0 9.62e-09 0.0007 9.623e-09 0 9.817e-09 0 9.82e-09 0.0007 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0007 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0007 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0007 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0007 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0007 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0007 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0007 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0007 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0007 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0007 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0007 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0007 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0007 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0007 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0007 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0007 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0007 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0007 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0007 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0007 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0007 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0007 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0007 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0007 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0007 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0007 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0007 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0007 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0007 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0007 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0007 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0007 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0007 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0007 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0007 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0007 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0007 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0007 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0007 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0007 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0007 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0007 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0007 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0007 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0007 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0007 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0007 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0007 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0007 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0007 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0007 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0007 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0007 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0007 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0007 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0007 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0007 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0007 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0007 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0007 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0007 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0007 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0007 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0007 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0007 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0007 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0007 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0007 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0007 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0007 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0007 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0007 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0007 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0007 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0007 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0007 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0007 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0007 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0007 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0007 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0007 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0007 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0007 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0007 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0007 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0007 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0007 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0007 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0007 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0007 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0007 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0007 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0007 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0007 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0007 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0007 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0007 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0007 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0007 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0007 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0007 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0007 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0007 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0007 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0007 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0007 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0007 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0007 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0007 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0007 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0007 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0007 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0007 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0007 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0007 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0007 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0007 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0007 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0007 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0007 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0007 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0007 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0007 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0007 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0007 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0007 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0007 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0007 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0007 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0007 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0007 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0007 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0007 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0007 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0007 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0007 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0007 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0007 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0007 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0007 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0007 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0007 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0007 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0007 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0007 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0007 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0007 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0007 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0007 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0007 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0007 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0007 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0007 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0007 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0007 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0007 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0007 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0007 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0007 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0007 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0007 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0007 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0007 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0007 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0007 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0007 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0007 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0007 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0007 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0007 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0007 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0007 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0007 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0007 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0007 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0007 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0007 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0007 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0007 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0007 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0007 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0007 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0007 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0007 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0007 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0007 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0007 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0007 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0007 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0007 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0007 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0007 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0007 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0007 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0007 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0007 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0007 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0007 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0007 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0007 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0007 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0007 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0007 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0007 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0007 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0007 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0007 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0007 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0007 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0007 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0007 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0007 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0007 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0007 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0007 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0007 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0007 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0007 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0007 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0007 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0007 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0007 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0007 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0007 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0007 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0007 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0007 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0007 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0007 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0007 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0007 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0007 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0007 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0007 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0007 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0007 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0007 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0007 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0007 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0007 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0007 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0007 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0007 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0007 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0007 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0007 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0007 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0007 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0007 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0007 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0007 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0007 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0007 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0007 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0007 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0007 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0007 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0007 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0007 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0007 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0007 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0007 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0007 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0007 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0007 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0007 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0007 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0007 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0007 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0007 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0007 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0007 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0007 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0007 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0007 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0007 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0007 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0007 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0007 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0007 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0007 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0007 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0007 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0007 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0007 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0007 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0007 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0007 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0007 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0007 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0007 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0007 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0007 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0007 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0007 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0007 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0007 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0007 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0007 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0007 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0007 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0007 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0007 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0007 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0007 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0007 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0007 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0007 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0007 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0007 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0007 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0007 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0007 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0007 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0007 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0007 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0007 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0007 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0007 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0007 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0007 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0007 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0007 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0007 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0007 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0007 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0007 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0007 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0007 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0007 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0007 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0007 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0007 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0007 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0007 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0007 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0007 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0007 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0007 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0007 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0007 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0007 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0007 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0007 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0007 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0007 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0007 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0007 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0007 7.9623e-08 0)
L_IP7_12|1 IP7_1_OUT _IP7_12|A1  2.067833848e-12
L_IP7_12|2 _IP7_12|A1 _IP7_12|A2  4.135667696e-12
L_IP7_12|3 _IP7_12|A3 _IP7_12|A4  8.271335392e-12
L_IP7_12|T T2B _IP7_12|T1  2.067833848e-12
L_IP7_12|4 _IP7_12|T1 _IP7_12|T2  4.135667696e-12
L_IP7_12|5 _IP7_12|A4 _IP7_12|Q1  4.135667696e-12
L_IP7_12|6 _IP7_12|Q1 IP7_2_OUT_TX  2.067833848e-12
IT30|T 0 T30  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_S0_23|1 S0_2 _S0_23|A1  2.067833848e-12
L_S0_23|2 _S0_23|A1 _S0_23|A2  4.135667696e-12
L_S0_23|3 _S0_23|A3 _S0_23|A4  8.271335392e-12
L_S0_23|T T30 _S0_23|T1  2.067833848e-12
L_S0_23|4 _S0_23|T1 _S0_23|T2  4.135667696e-12
L_S0_23|5 _S0_23|A4 _S0_23|Q1  4.135667696e-12
L_S0_23|6 _S0_23|Q1 S0_3_TX  2.067833848e-12
IT31|T 0 T31  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_S1_23|1 S1_2 _S1_23|A1  2.067833848e-12
L_S1_23|2 _S1_23|A1 _S1_23|A2  4.135667696e-12
L_S1_23|3 _S1_23|A3 _S1_23|A4  8.271335392e-12
L_S1_23|T T31 _S1_23|T1  2.067833848e-12
L_S1_23|4 _S1_23|T1 _S1_23|T2  4.135667696e-12
L_S1_23|5 _S1_23|A4 _S1_23|Q1  4.135667696e-12
L_S1_23|6 _S1_23|Q1 S1_3_TX  2.067833848e-12
IT32|T 0 T32  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_S2_23|1 S2_2 _S2_23|A1  2.067833848e-12
L_S2_23|2 _S2_23|A1 _S2_23|A2  4.135667696e-12
L_S2_23|3 _S2_23|A3 _S2_23|A4  8.271335392e-12
L_S2_23|T T32 _S2_23|T1  2.067833848e-12
L_S2_23|4 _S2_23|T1 _S2_23|T2  4.135667696e-12
L_S2_23|5 _S2_23|A4 _S2_23|Q1  4.135667696e-12
L_S2_23|6 _S2_23|Q1 S2_3_TX  2.067833848e-12
IT33|T 0 T33  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_S3_23|A1 G2_2_OUT _S3_23|A1  2.067833848e-12
L_S3_23|A2 _S3_23|A1 _S3_23|A2  4.135667696e-12
L_S3_23|A3 _S3_23|A3 _S3_23|AB  8.271335392e-12
L_S3_23|B1 IP3_2_OUT _S3_23|B1  2.067833848e-12
L_S3_23|B2 _S3_23|B1 _S3_23|B2  4.135667696e-12
L_S3_23|B3 _S3_23|B3 _S3_23|AB  8.271335392e-12
L_S3_23|T1 T33 _S3_23|T1  2.067833848e-12
L_S3_23|T2 _S3_23|T1 _S3_23|T2  4.135667696e-12
L_S3_23|Q2 _S3_23|ABTQ _S3_23|Q1  4.135667696e-12
L_S3_23|Q1 _S3_23|Q1 S3_3_TX  2.067833848e-12
IT34|T 0 T34  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_S4_23|A1 G3_2_OUT _S4_23|A1  2.067833848e-12
L_S4_23|A2 _S4_23|A1 _S4_23|A2  4.135667696e-12
L_S4_23|A3 _S4_23|A3 _S4_23|AB  8.271335392e-12
L_S4_23|B1 P4_2_OUT _S4_23|B1  2.067833848e-12
L_S4_23|B2 _S4_23|B1 _S4_23|B2  4.135667696e-12
L_S4_23|B3 _S4_23|B3 _S4_23|AB  8.271335392e-12
L_S4_23|T1 T34 _S4_23|T1  2.067833848e-12
L_S4_23|T2 _S4_23|T1 _S4_23|T2  4.135667696e-12
L_S4_23|Q2 _S4_23|ABTQ _S4_23|Q1  4.135667696e-12
L_S4_23|Q1 _S4_23|Q1 S4_3_TX  2.067833848e-12
IT35|T 0 T35  PWL(0 0 7e-12 0 1e-11 0.0028 1.3e-11 0 2.07e-10 0 2.1e-10 0.0028 2.13e-10 0 4.07e-10 0 4.1e-10 0.0028 4.13e-10 0 6.07e-10 0 6.1e-10 0.0028 6.13e-10 0 8.07e-10 0 8.1e-10 0.0028 8.13e-10 0 1.007e-09 0 1.01e-09 0.0028 1.013e-09 0 1.207e-09 0 1.21e-09 0.0028 1.213e-09 0 1.407e-09 0 1.41e-09 0.0028 1.413e-09 0 1.607e-09 0 1.61e-09 0.0028 1.613e-09 0 1.807e-09 0 1.81e-09 0.0028 1.813e-09 0 2.007e-09 0 2.01e-09 0.0028 2.013e-09 0 2.207e-09 0 2.21e-09 0.0028 2.213e-09 0 2.407e-09 0 2.41e-09 0.0028 2.413e-09 0 2.607e-09 0 2.61e-09 0.0028 2.613e-09 0 2.807e-09 0 2.81e-09 0.0028 2.813e-09 0 3.007e-09 0 3.01e-09 0.0028 3.013e-09 0 3.207e-09 0 3.21e-09 0.0028 3.213e-09 0 3.407e-09 0 3.41e-09 0.0028 3.413e-09 0 3.607e-09 0 3.61e-09 0.0028 3.613e-09 0 3.807e-09 0 3.81e-09 0.0028 3.813e-09 0 4.007e-09 0 4.01e-09 0.0028 4.013e-09 0 4.207e-09 0 4.21e-09 0.0028 4.213e-09 0 4.407e-09 0 4.41e-09 0.0028 4.413e-09 0 4.607e-09 0 4.61e-09 0.0028 4.613e-09 0 4.807e-09 0 4.81e-09 0.0028 4.813e-09 0 5.007e-09 0 5.01e-09 0.0028 5.013e-09 0 5.207e-09 0 5.21e-09 0.0028 5.213e-09 0 5.407e-09 0 5.41e-09 0.0028 5.413e-09 0 5.607e-09 0 5.61e-09 0.0028 5.613e-09 0 5.807e-09 0 5.81e-09 0.0028 5.813e-09 0 6.007e-09 0 6.01e-09 0.0028 6.013e-09 0 6.207e-09 0 6.21e-09 0.0028 6.213e-09 0 6.407e-09 0 6.41e-09 0.0028 6.413e-09 0 6.607e-09 0 6.61e-09 0.0028 6.613e-09 0 6.807e-09 0 6.81e-09 0.0028 6.813e-09 0 7.007e-09 0 7.01e-09 0.0028 7.013e-09 0 7.207e-09 0 7.21e-09 0.0028 7.213e-09 0 7.407e-09 0 7.41e-09 0.0028 7.413e-09 0 7.607e-09 0 7.61e-09 0.0028 7.613e-09 0 7.807e-09 0 7.81e-09 0.0028 7.813e-09 0 8.007e-09 0 8.01e-09 0.0028 8.013e-09 0 8.207e-09 0 8.21e-09 0.0028 8.213e-09 0 8.407e-09 0 8.41e-09 0.0028 8.413e-09 0 8.607e-09 0 8.61e-09 0.0028 8.613e-09 0 8.807e-09 0 8.81e-09 0.0028 8.813e-09 0 9.007e-09 0 9.01e-09 0.0028 9.013e-09 0 9.207e-09 0 9.21e-09 0.0028 9.213e-09 0 9.407e-09 0 9.41e-09 0.0028 9.413e-09 0 9.607e-09 0 9.61e-09 0.0028 9.613e-09 0 9.807e-09 0 9.81e-09 0.0028 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0028 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0028 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0028 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0028 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0028 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0028 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0028 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0028 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0028 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0028 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0028 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0028 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0028 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0028 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0028 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0028 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0028 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0028 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0028 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0028 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0028 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0028 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0028 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0028 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0028 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0028 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0028 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0028 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0028 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0028 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0028 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0028 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0028 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0028 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0028 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0028 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0028 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0028 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0028 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0028 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0028 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0028 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0028 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0028 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0028 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0028 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0028 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0028 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0028 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0028 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0028 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0028 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0028 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0028 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0028 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0028 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0028 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0028 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0028 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0028 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0028 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0028 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0028 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0028 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0028 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0028 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0028 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0028 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0028 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0028 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0028 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0028 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0028 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0028 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0028 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0028 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0028 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0028 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0028 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0028 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0028 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0028 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0028 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0028 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0028 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0028 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0028 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0028 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0028 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0028 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0028 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0028 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0028 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0028 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0028 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0028 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0028 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0028 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0028 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0028 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0028 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0028 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0028 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0028 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0028 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0028 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0028 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0028 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0028 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0028 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0028 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0028 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0028 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0028 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0028 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0028 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0028 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0028 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0028 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0028 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0028 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0028 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0028 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0028 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0028 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0028 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0028 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0028 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0028 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0028 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0028 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0028 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0028 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0028 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0028 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0028 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0028 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0028 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0028 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0028 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0028 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0028 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0028 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0028 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0028 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0028 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0028 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0028 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0028 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0028 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0028 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0028 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0028 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0028 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0028 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0028 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0028 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0028 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0028 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0028 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0028 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0028 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0028 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0028 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0028 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0028 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0028 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0028 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0028 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0028 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0028 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0028 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0028 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0028 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0028 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0028 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0028 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0028 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0028 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0028 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0028 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0028 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0028 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0028 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0028 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0028 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0028 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0028 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0028 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0028 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0028 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0028 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0028 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0028 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0028 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0028 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0028 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0028 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0028 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0028 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0028 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0028 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0028 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0028 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0028 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0028 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0028 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0028 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0028 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0028 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0028 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0028 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0028 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0028 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0028 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0028 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0028 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0028 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0028 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0028 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0028 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0028 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0028 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0028 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0028 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0028 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0028 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0028 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0028 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0028 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0028 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0028 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0028 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0028 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0028 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0028 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0028 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0028 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0028 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0028 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0028 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0028 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0028 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0028 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0028 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0028 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0028 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0028 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0028 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0028 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0028 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0028 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0028 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0028 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0028 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0028 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0028 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0028 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0028 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0028 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0028 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0028 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0028 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0028 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0028 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0028 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0028 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0028 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0028 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0028 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0028 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0028 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0028 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0028 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0028 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0028 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0028 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0028 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0028 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0028 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0028 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0028 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0028 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0028 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0028 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0028 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0028 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0028 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0028 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0028 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0028 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0028 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0028 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0028 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0028 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0028 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0028 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0028 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0028 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0028 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0028 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0028 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0028 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0028 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0028 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0028 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0028 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0028 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0028 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0028 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0028 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0028 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0028 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0028 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0028 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0028 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0028 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0028 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0028 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0028 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0028 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0028 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0028 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0028 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0028 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0028 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0028 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0028 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0028 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0028 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0028 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0028 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0028 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0028 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0028 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0028 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0028 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0028 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0028 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0028 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0028 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0028 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0028 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0028 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0028 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0028 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0028 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0028 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0028 7.9613e-08 0)
IT36|T 0 T36  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_IP5_23|1 IP5_2_OUT _IP5_23|A1  2.067833848e-12
L_IP5_23|2 _IP5_23|A1 _IP5_23|A2  4.135667696e-12
L_IP5_23|3 _IP5_23|A3 _IP5_23|A4  8.271335392e-12
L_IP5_23|T T36 _IP5_23|T1  2.067833848e-12
L_IP5_23|4 _IP5_23|T1 _IP5_23|T2  4.135667696e-12
L_IP5_23|5 _IP5_23|A4 _IP5_23|Q1  4.135667696e-12
L_IP5_23|6 _IP5_23|Q1 IP5_3_OUT_TX  2.067833848e-12
IT37|T 0 T37  PWL(0 0 7e-12 0 1e-11 0.0028 1.3e-11 0 2.07e-10 0 2.1e-10 0.0028 2.13e-10 0 4.07e-10 0 4.1e-10 0.0028 4.13e-10 0 6.07e-10 0 6.1e-10 0.0028 6.13e-10 0 8.07e-10 0 8.1e-10 0.0028 8.13e-10 0 1.007e-09 0 1.01e-09 0.0028 1.013e-09 0 1.207e-09 0 1.21e-09 0.0028 1.213e-09 0 1.407e-09 0 1.41e-09 0.0028 1.413e-09 0 1.607e-09 0 1.61e-09 0.0028 1.613e-09 0 1.807e-09 0 1.81e-09 0.0028 1.813e-09 0 2.007e-09 0 2.01e-09 0.0028 2.013e-09 0 2.207e-09 0 2.21e-09 0.0028 2.213e-09 0 2.407e-09 0 2.41e-09 0.0028 2.413e-09 0 2.607e-09 0 2.61e-09 0.0028 2.613e-09 0 2.807e-09 0 2.81e-09 0.0028 2.813e-09 0 3.007e-09 0 3.01e-09 0.0028 3.013e-09 0 3.207e-09 0 3.21e-09 0.0028 3.213e-09 0 3.407e-09 0 3.41e-09 0.0028 3.413e-09 0 3.607e-09 0 3.61e-09 0.0028 3.613e-09 0 3.807e-09 0 3.81e-09 0.0028 3.813e-09 0 4.007e-09 0 4.01e-09 0.0028 4.013e-09 0 4.207e-09 0 4.21e-09 0.0028 4.213e-09 0 4.407e-09 0 4.41e-09 0.0028 4.413e-09 0 4.607e-09 0 4.61e-09 0.0028 4.613e-09 0 4.807e-09 0 4.81e-09 0.0028 4.813e-09 0 5.007e-09 0 5.01e-09 0.0028 5.013e-09 0 5.207e-09 0 5.21e-09 0.0028 5.213e-09 0 5.407e-09 0 5.41e-09 0.0028 5.413e-09 0 5.607e-09 0 5.61e-09 0.0028 5.613e-09 0 5.807e-09 0 5.81e-09 0.0028 5.813e-09 0 6.007e-09 0 6.01e-09 0.0028 6.013e-09 0 6.207e-09 0 6.21e-09 0.0028 6.213e-09 0 6.407e-09 0 6.41e-09 0.0028 6.413e-09 0 6.607e-09 0 6.61e-09 0.0028 6.613e-09 0 6.807e-09 0 6.81e-09 0.0028 6.813e-09 0 7.007e-09 0 7.01e-09 0.0028 7.013e-09 0 7.207e-09 0 7.21e-09 0.0028 7.213e-09 0 7.407e-09 0 7.41e-09 0.0028 7.413e-09 0 7.607e-09 0 7.61e-09 0.0028 7.613e-09 0 7.807e-09 0 7.81e-09 0.0028 7.813e-09 0 8.007e-09 0 8.01e-09 0.0028 8.013e-09 0 8.207e-09 0 8.21e-09 0.0028 8.213e-09 0 8.407e-09 0 8.41e-09 0.0028 8.413e-09 0 8.607e-09 0 8.61e-09 0.0028 8.613e-09 0 8.807e-09 0 8.81e-09 0.0028 8.813e-09 0 9.007e-09 0 9.01e-09 0.0028 9.013e-09 0 9.207e-09 0 9.21e-09 0.0028 9.213e-09 0 9.407e-09 0 9.41e-09 0.0028 9.413e-09 0 9.607e-09 0 9.61e-09 0.0028 9.613e-09 0 9.807e-09 0 9.81e-09 0.0028 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0028 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0028 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0028 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0028 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0028 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0028 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0028 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0028 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0028 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0028 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0028 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0028 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0028 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0028 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0028 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0028 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0028 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0028 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0028 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0028 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0028 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0028 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0028 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0028 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0028 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0028 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0028 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0028 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0028 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0028 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0028 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0028 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0028 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0028 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0028 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0028 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0028 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0028 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0028 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0028 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0028 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0028 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0028 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0028 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0028 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0028 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0028 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0028 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0028 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0028 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0028 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0028 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0028 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0028 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0028 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0028 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0028 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0028 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0028 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0028 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0028 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0028 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0028 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0028 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0028 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0028 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0028 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0028 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0028 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0028 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0028 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0028 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0028 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0028 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0028 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0028 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0028 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0028 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0028 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0028 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0028 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0028 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0028 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0028 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0028 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0028 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0028 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0028 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0028 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0028 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0028 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0028 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0028 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0028 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0028 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0028 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0028 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0028 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0028 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0028 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0028 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0028 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0028 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0028 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0028 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0028 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0028 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0028 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0028 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0028 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0028 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0028 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0028 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0028 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0028 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0028 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0028 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0028 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0028 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0028 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0028 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0028 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0028 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0028 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0028 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0028 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0028 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0028 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0028 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0028 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0028 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0028 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0028 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0028 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0028 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0028 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0028 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0028 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0028 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0028 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0028 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0028 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0028 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0028 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0028 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0028 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0028 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0028 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0028 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0028 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0028 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0028 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0028 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0028 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0028 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0028 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0028 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0028 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0028 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0028 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0028 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0028 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0028 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0028 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0028 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0028 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0028 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0028 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0028 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0028 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0028 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0028 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0028 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0028 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0028 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0028 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0028 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0028 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0028 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0028 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0028 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0028 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0028 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0028 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0028 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0028 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0028 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0028 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0028 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0028 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0028 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0028 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0028 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0028 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0028 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0028 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0028 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0028 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0028 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0028 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0028 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0028 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0028 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0028 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0028 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0028 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0028 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0028 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0028 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0028 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0028 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0028 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0028 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0028 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0028 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0028 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0028 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0028 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0028 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0028 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0028 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0028 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0028 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0028 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0028 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0028 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0028 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0028 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0028 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0028 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0028 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0028 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0028 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0028 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0028 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0028 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0028 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0028 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0028 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0028 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0028 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0028 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0028 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0028 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0028 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0028 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0028 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0028 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0028 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0028 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0028 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0028 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0028 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0028 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0028 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0028 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0028 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0028 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0028 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0028 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0028 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0028 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0028 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0028 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0028 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0028 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0028 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0028 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0028 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0028 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0028 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0028 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0028 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0028 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0028 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0028 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0028 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0028 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0028 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0028 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0028 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0028 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0028 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0028 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0028 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0028 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0028 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0028 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0028 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0028 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0028 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0028 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0028 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0028 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0028 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0028 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0028 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0028 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0028 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0028 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0028 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0028 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0028 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0028 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0028 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0028 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0028 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0028 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0028 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0028 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0028 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0028 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0028 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0028 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0028 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0028 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0028 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0028 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0028 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0028 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0028 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0028 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0028 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0028 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0028 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0028 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0028 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0028 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0028 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0028 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0028 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0028 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0028 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0028 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0028 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0028 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0028 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0028 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0028 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0028 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0028 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0028 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0028 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0028 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0028 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0028 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0028 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0028 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0028 7.9613e-08 0)
IT38|T 0 T38  PWL(0 0 7e-12 0 1e-11 0.0014 1.3e-11 0 2.07e-10 0 2.1e-10 0.0014 2.13e-10 0 4.07e-10 0 4.1e-10 0.0014 4.13e-10 0 6.07e-10 0 6.1e-10 0.0014 6.13e-10 0 8.07e-10 0 8.1e-10 0.0014 8.13e-10 0 1.007e-09 0 1.01e-09 0.0014 1.013e-09 0 1.207e-09 0 1.21e-09 0.0014 1.213e-09 0 1.407e-09 0 1.41e-09 0.0014 1.413e-09 0 1.607e-09 0 1.61e-09 0.0014 1.613e-09 0 1.807e-09 0 1.81e-09 0.0014 1.813e-09 0 2.007e-09 0 2.01e-09 0.0014 2.013e-09 0 2.207e-09 0 2.21e-09 0.0014 2.213e-09 0 2.407e-09 0 2.41e-09 0.0014 2.413e-09 0 2.607e-09 0 2.61e-09 0.0014 2.613e-09 0 2.807e-09 0 2.81e-09 0.0014 2.813e-09 0 3.007e-09 0 3.01e-09 0.0014 3.013e-09 0 3.207e-09 0 3.21e-09 0.0014 3.213e-09 0 3.407e-09 0 3.41e-09 0.0014 3.413e-09 0 3.607e-09 0 3.61e-09 0.0014 3.613e-09 0 3.807e-09 0 3.81e-09 0.0014 3.813e-09 0 4.007e-09 0 4.01e-09 0.0014 4.013e-09 0 4.207e-09 0 4.21e-09 0.0014 4.213e-09 0 4.407e-09 0 4.41e-09 0.0014 4.413e-09 0 4.607e-09 0 4.61e-09 0.0014 4.613e-09 0 4.807e-09 0 4.81e-09 0.0014 4.813e-09 0 5.007e-09 0 5.01e-09 0.0014 5.013e-09 0 5.207e-09 0 5.21e-09 0.0014 5.213e-09 0 5.407e-09 0 5.41e-09 0.0014 5.413e-09 0 5.607e-09 0 5.61e-09 0.0014 5.613e-09 0 5.807e-09 0 5.81e-09 0.0014 5.813e-09 0 6.007e-09 0 6.01e-09 0.0014 6.013e-09 0 6.207e-09 0 6.21e-09 0.0014 6.213e-09 0 6.407e-09 0 6.41e-09 0.0014 6.413e-09 0 6.607e-09 0 6.61e-09 0.0014 6.613e-09 0 6.807e-09 0 6.81e-09 0.0014 6.813e-09 0 7.007e-09 0 7.01e-09 0.0014 7.013e-09 0 7.207e-09 0 7.21e-09 0.0014 7.213e-09 0 7.407e-09 0 7.41e-09 0.0014 7.413e-09 0 7.607e-09 0 7.61e-09 0.0014 7.613e-09 0 7.807e-09 0 7.81e-09 0.0014 7.813e-09 0 8.007e-09 0 8.01e-09 0.0014 8.013e-09 0 8.207e-09 0 8.21e-09 0.0014 8.213e-09 0 8.407e-09 0 8.41e-09 0.0014 8.413e-09 0 8.607e-09 0 8.61e-09 0.0014 8.613e-09 0 8.807e-09 0 8.81e-09 0.0014 8.813e-09 0 9.007e-09 0 9.01e-09 0.0014 9.013e-09 0 9.207e-09 0 9.21e-09 0.0014 9.213e-09 0 9.407e-09 0 9.41e-09 0.0014 9.413e-09 0 9.607e-09 0 9.61e-09 0.0014 9.613e-09 0 9.807e-09 0 9.81e-09 0.0014 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0014 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0014 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0014 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0014 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0014 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0014 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0014 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0014 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0014 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0014 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0014 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0014 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0014 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0014 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0014 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0014 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0014 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0014 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0014 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0014 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0014 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0014 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0014 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0014 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0014 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0014 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0014 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0014 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0014 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0014 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0014 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0014 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0014 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0014 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0014 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0014 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0014 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0014 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0014 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0014 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0014 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0014 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0014 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0014 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0014 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0014 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0014 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0014 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0014 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0014 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0014 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0014 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0014 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0014 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0014 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0014 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0014 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0014 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0014 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0014 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0014 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0014 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0014 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0014 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0014 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0014 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0014 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0014 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0014 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0014 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0014 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0014 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0014 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0014 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0014 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0014 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0014 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0014 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0014 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0014 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0014 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0014 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0014 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0014 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0014 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0014 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0014 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0014 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0014 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0014 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0014 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0014 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0014 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0014 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0014 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0014 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0014 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0014 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0014 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0014 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0014 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0014 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0014 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0014 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0014 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0014 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0014 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0014 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0014 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0014 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0014 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0014 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0014 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0014 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0014 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0014 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0014 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0014 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0014 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0014 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0014 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0014 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0014 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0014 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0014 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0014 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0014 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0014 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0014 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0014 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0014 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0014 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0014 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0014 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0014 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0014 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0014 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0014 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0014 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0014 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0014 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0014 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0014 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0014 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0014 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0014 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0014 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0014 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0014 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0014 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0014 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0014 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0014 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0014 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0014 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0014 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0014 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0014 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0014 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0014 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0014 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0014 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0014 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0014 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0014 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0014 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0014 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0014 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0014 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0014 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0014 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0014 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0014 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0014 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0014 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0014 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0014 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0014 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0014 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0014 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0014 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0014 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0014 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0014 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0014 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0014 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0014 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0014 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0014 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0014 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0014 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0014 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0014 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0014 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0014 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0014 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0014 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0014 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0014 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0014 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0014 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0014 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0014 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0014 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0014 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0014 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0014 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0014 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0014 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0014 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0014 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0014 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0014 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0014 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0014 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0014 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0014 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0014 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0014 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0014 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0014 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0014 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0014 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0014 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0014 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0014 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0014 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0014 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0014 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0014 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0014 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0014 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0014 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0014 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0014 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0014 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0014 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0014 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0014 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0014 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0014 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0014 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0014 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0014 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0014 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0014 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0014 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0014 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0014 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0014 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0014 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0014 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0014 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0014 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0014 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0014 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0014 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0014 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0014 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0014 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0014 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0014 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0014 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0014 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0014 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0014 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0014 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0014 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0014 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0014 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0014 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0014 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0014 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0014 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0014 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0014 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0014 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0014 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0014 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0014 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0014 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0014 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0014 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0014 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0014 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0014 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0014 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0014 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0014 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0014 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0014 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0014 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0014 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0014 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0014 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0014 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0014 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0014 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0014 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0014 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0014 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0014 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0014 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0014 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0014 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0014 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0014 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0014 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0014 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0014 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0014 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0014 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0014 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0014 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0014 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0014 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0014 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0014 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0014 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0014 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0014 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0014 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0014 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0014 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0014 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0014 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0014 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0014 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0014 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0014 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0014 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0014 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0014 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0014 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0014 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0014 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0014 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0014 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0014 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0014 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0014 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0014 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0014 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0014 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0014 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0014 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0014 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0014 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0014 7.9613e-08 0)
IT39|T 0 T39  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_IP7_23|1 IP7_2_OUT _IP7_23|A1  2.067833848e-12
L_IP7_23|2 _IP7_23|A1 _IP7_23|A2  4.135667696e-12
L_IP7_23|3 _IP7_23|A3 _IP7_23|A4  8.271335392e-12
L_IP7_23|T T39 _IP7_23|T1  2.067833848e-12
L_IP7_23|4 _IP7_23|T1 _IP7_23|T2  4.135667696e-12
L_IP7_23|5 _IP7_23|A4 _IP7_23|Q1  4.135667696e-12
L_IP7_23|6 _IP7_23|Q1 IP7_3_OUT_TX  2.067833848e-12
IT3A|T 0 T3A  PWL(0 0 7e-12 0 1e-11 0.0028 1.3e-11 0 2.07e-10 0 2.1e-10 0.0028 2.13e-10 0 4.07e-10 0 4.1e-10 0.0028 4.13e-10 0 6.07e-10 0 6.1e-10 0.0028 6.13e-10 0 8.07e-10 0 8.1e-10 0.0028 8.13e-10 0 1.007e-09 0 1.01e-09 0.0028 1.013e-09 0 1.207e-09 0 1.21e-09 0.0028 1.213e-09 0 1.407e-09 0 1.41e-09 0.0028 1.413e-09 0 1.607e-09 0 1.61e-09 0.0028 1.613e-09 0 1.807e-09 0 1.81e-09 0.0028 1.813e-09 0 2.007e-09 0 2.01e-09 0.0028 2.013e-09 0 2.207e-09 0 2.21e-09 0.0028 2.213e-09 0 2.407e-09 0 2.41e-09 0.0028 2.413e-09 0 2.607e-09 0 2.61e-09 0.0028 2.613e-09 0 2.807e-09 0 2.81e-09 0.0028 2.813e-09 0 3.007e-09 0 3.01e-09 0.0028 3.013e-09 0 3.207e-09 0 3.21e-09 0.0028 3.213e-09 0 3.407e-09 0 3.41e-09 0.0028 3.413e-09 0 3.607e-09 0 3.61e-09 0.0028 3.613e-09 0 3.807e-09 0 3.81e-09 0.0028 3.813e-09 0 4.007e-09 0 4.01e-09 0.0028 4.013e-09 0 4.207e-09 0 4.21e-09 0.0028 4.213e-09 0 4.407e-09 0 4.41e-09 0.0028 4.413e-09 0 4.607e-09 0 4.61e-09 0.0028 4.613e-09 0 4.807e-09 0 4.81e-09 0.0028 4.813e-09 0 5.007e-09 0 5.01e-09 0.0028 5.013e-09 0 5.207e-09 0 5.21e-09 0.0028 5.213e-09 0 5.407e-09 0 5.41e-09 0.0028 5.413e-09 0 5.607e-09 0 5.61e-09 0.0028 5.613e-09 0 5.807e-09 0 5.81e-09 0.0028 5.813e-09 0 6.007e-09 0 6.01e-09 0.0028 6.013e-09 0 6.207e-09 0 6.21e-09 0.0028 6.213e-09 0 6.407e-09 0 6.41e-09 0.0028 6.413e-09 0 6.607e-09 0 6.61e-09 0.0028 6.613e-09 0 6.807e-09 0 6.81e-09 0.0028 6.813e-09 0 7.007e-09 0 7.01e-09 0.0028 7.013e-09 0 7.207e-09 0 7.21e-09 0.0028 7.213e-09 0 7.407e-09 0 7.41e-09 0.0028 7.413e-09 0 7.607e-09 0 7.61e-09 0.0028 7.613e-09 0 7.807e-09 0 7.81e-09 0.0028 7.813e-09 0 8.007e-09 0 8.01e-09 0.0028 8.013e-09 0 8.207e-09 0 8.21e-09 0.0028 8.213e-09 0 8.407e-09 0 8.41e-09 0.0028 8.413e-09 0 8.607e-09 0 8.61e-09 0.0028 8.613e-09 0 8.807e-09 0 8.81e-09 0.0028 8.813e-09 0 9.007e-09 0 9.01e-09 0.0028 9.013e-09 0 9.207e-09 0 9.21e-09 0.0028 9.213e-09 0 9.407e-09 0 9.41e-09 0.0028 9.413e-09 0 9.607e-09 0 9.61e-09 0.0028 9.613e-09 0 9.807e-09 0 9.81e-09 0.0028 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0028 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0028 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0028 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0028 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0028 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0028 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0028 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0028 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0028 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0028 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0028 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0028 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0028 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0028 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0028 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0028 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0028 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0028 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0028 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0028 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0028 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0028 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0028 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0028 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0028 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0028 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0028 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0028 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0028 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0028 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0028 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0028 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0028 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0028 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0028 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0028 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0028 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0028 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0028 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0028 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0028 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0028 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0028 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0028 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0028 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0028 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0028 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0028 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0028 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0028 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0028 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0028 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0028 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0028 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0028 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0028 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0028 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0028 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0028 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0028 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0028 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0028 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0028 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0028 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0028 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0028 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0028 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0028 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0028 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0028 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0028 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0028 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0028 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0028 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0028 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0028 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0028 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0028 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0028 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0028 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0028 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0028 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0028 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0028 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0028 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0028 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0028 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0028 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0028 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0028 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0028 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0028 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0028 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0028 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0028 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0028 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0028 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0028 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0028 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0028 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0028 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0028 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0028 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0028 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0028 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0028 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0028 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0028 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0028 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0028 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0028 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0028 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0028 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0028 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0028 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0028 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0028 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0028 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0028 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0028 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0028 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0028 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0028 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0028 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0028 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0028 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0028 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0028 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0028 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0028 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0028 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0028 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0028 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0028 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0028 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0028 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0028 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0028 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0028 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0028 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0028 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0028 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0028 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0028 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0028 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0028 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0028 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0028 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0028 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0028 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0028 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0028 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0028 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0028 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0028 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0028 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0028 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0028 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0028 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0028 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0028 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0028 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0028 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0028 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0028 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0028 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0028 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0028 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0028 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0028 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0028 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0028 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0028 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0028 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0028 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0028 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0028 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0028 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0028 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0028 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0028 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0028 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0028 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0028 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0028 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0028 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0028 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0028 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0028 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0028 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0028 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0028 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0028 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0028 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0028 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0028 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0028 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0028 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0028 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0028 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0028 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0028 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0028 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0028 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0028 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0028 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0028 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0028 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0028 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0028 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0028 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0028 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0028 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0028 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0028 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0028 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0028 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0028 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0028 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0028 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0028 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0028 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0028 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0028 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0028 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0028 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0028 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0028 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0028 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0028 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0028 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0028 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0028 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0028 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0028 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0028 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0028 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0028 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0028 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0028 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0028 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0028 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0028 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0028 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0028 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0028 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0028 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0028 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0028 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0028 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0028 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0028 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0028 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0028 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0028 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0028 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0028 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0028 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0028 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0028 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0028 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0028 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0028 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0028 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0028 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0028 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0028 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0028 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0028 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0028 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0028 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0028 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0028 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0028 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0028 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0028 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0028 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0028 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0028 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0028 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0028 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0028 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0028 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0028 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0028 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0028 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0028 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0028 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0028 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0028 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0028 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0028 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0028 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0028 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0028 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0028 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0028 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0028 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0028 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0028 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0028 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0028 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0028 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0028 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0028 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0028 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0028 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0028 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0028 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0028 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0028 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0028 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0028 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0028 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0028 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0028 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0028 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0028 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0028 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0028 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0028 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0028 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0028 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0028 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0028 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0028 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0028 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0028 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0028 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0028 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0028 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0028 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0028 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0028 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0028 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0028 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0028 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0028 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0028 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0028 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0028 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0028 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0028 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0028 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0028 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0028 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0028 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0028 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0028 7.9613e-08 0)
IT40|T 0 T40  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S0_34|1 S0_3 _S0_34|A1  2.067833848e-12
L_S0_34|2 _S0_34|A1 _S0_34|A2  4.135667696e-12
L_S0_34|3 _S0_34|A3 _S0_34|A4  8.271335392e-12
L_S0_34|T T40 _S0_34|T1  2.067833848e-12
L_S0_34|4 _S0_34|T1 _S0_34|T2  4.135667696e-12
L_S0_34|5 _S0_34|A4 _S0_34|Q1  4.135667696e-12
L_S0_34|6 _S0_34|Q1 S0_4_TX  2.067833848e-12
IT41|T 0 T41  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S1_34|1 S1_3 _S1_34|A1  2.067833848e-12
L_S1_34|2 _S1_34|A1 _S1_34|A2  4.135667696e-12
L_S1_34|3 _S1_34|A3 _S1_34|A4  8.271335392e-12
L_S1_34|T T41 _S1_34|T1  2.067833848e-12
L_S1_34|4 _S1_34|T1 _S1_34|T2  4.135667696e-12
L_S1_34|5 _S1_34|A4 _S1_34|Q1  4.135667696e-12
L_S1_34|6 _S1_34|Q1 S1_4_TX  2.067833848e-12
IT42|T 0 T42  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S2_34|1 S2_3 _S2_34|A1  2.067833848e-12
L_S2_34|2 _S2_34|A1 _S2_34|A2  4.135667696e-12
L_S2_34|3 _S2_34|A3 _S2_34|A4  8.271335392e-12
L_S2_34|T T42 _S2_34|T1  2.067833848e-12
L_S2_34|4 _S2_34|T1 _S2_34|T2  4.135667696e-12
L_S2_34|5 _S2_34|A4 _S2_34|Q1  4.135667696e-12
L_S2_34|6 _S2_34|Q1 S2_4_TX  2.067833848e-12
IT43|T 0 T43  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S3_34|1 S3_3 _S3_34|A1  2.067833848e-12
L_S3_34|2 _S3_34|A1 _S3_34|A2  4.135667696e-12
L_S3_34|3 _S3_34|A3 _S3_34|A4  8.271335392e-12
L_S3_34|T T43 _S3_34|T1  2.067833848e-12
L_S3_34|4 _S3_34|T1 _S3_34|T2  4.135667696e-12
L_S3_34|5 _S3_34|A4 _S3_34|Q1  4.135667696e-12
L_S3_34|6 _S3_34|Q1 S3_4_TX  2.067833848e-12
IT44|T 0 T44  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S4_34|1 S4_3 _S4_34|A1  2.067833848e-12
L_S4_34|2 _S4_34|A1 _S4_34|A2  4.135667696e-12
L_S4_34|3 _S4_34|A3 _S4_34|A4  8.271335392e-12
L_S4_34|T T44 _S4_34|T1  2.067833848e-12
L_S4_34|4 _S4_34|T1 _S4_34|T2  4.135667696e-12
L_S4_34|5 _S4_34|A4 _S4_34|Q1  4.135667696e-12
L_S4_34|6 _S4_34|Q1 S4_4_TX  2.067833848e-12
IT45|T 0 T45  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S5_34|A1 G4_3_OUT _S5_34|A1  2.067833848e-12
L_S5_34|A2 _S5_34|A1 _S5_34|A2  4.135667696e-12
L_S5_34|A3 _S5_34|A3 _S5_34|AB  8.271335392e-12
L_S5_34|B1 IP5_3_OUT _S5_34|B1  2.067833848e-12
L_S5_34|B2 _S5_34|B1 _S5_34|B2  4.135667696e-12
L_S5_34|B3 _S5_34|B3 _S5_34|AB  8.271335392e-12
L_S5_34|T1 T45 _S5_34|T1  2.067833848e-12
L_S5_34|T2 _S5_34|T1 _S5_34|T2  4.135667696e-12
L_S5_34|Q2 _S5_34|ABTQ _S5_34|Q1  4.135667696e-12
L_S5_34|Q1 _S5_34|Q1 S5_4_TX  2.067833848e-12
IT46|T 0 T46  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S6_34|A1 G5_3_OUT _S6_34|A1  2.067833848e-12
L_S6_34|A2 _S6_34|A1 _S6_34|A2  4.135667696e-12
L_S6_34|A3 _S6_34|A3 _S6_34|AB  8.271335392e-12
L_S6_34|B1 P6_3_OUT _S6_34|B1  2.067833848e-12
L_S6_34|B2 _S6_34|B1 _S6_34|B2  4.135667696e-12
L_S6_34|B3 _S6_34|B3 _S6_34|AB  8.271335392e-12
L_S6_34|T1 T46 _S6_34|T1  2.067833848e-12
L_S6_34|T2 _S6_34|T1 _S6_34|T2  4.135667696e-12
L_S6_34|Q2 _S6_34|ABTQ _S6_34|Q1  4.135667696e-12
L_S6_34|Q1 _S6_34|Q1 S6_4_TX  2.067833848e-12
IT47|T 0 T47  PWL(0 0 -3e-12 0 0 0.0028 3e-12 0 1.97e-10 0 2e-10 0.0028 2.03e-10 0 3.97e-10 0 4e-10 0.0028 4.03e-10 0 5.97e-10 0 6e-10 0.0028 6.03e-10 0 7.97e-10 0 8e-10 0.0028 8.03e-10 0 9.97e-10 0 1e-09 0.0028 1.003e-09 0 1.197e-09 0 1.2e-09 0.0028 1.203e-09 0 1.397e-09 0 1.4e-09 0.0028 1.403e-09 0 1.597e-09 0 1.6e-09 0.0028 1.603e-09 0 1.797e-09 0 1.8e-09 0.0028 1.803e-09 0 1.997e-09 0 2e-09 0.0028 2.003e-09 0 2.197e-09 0 2.2e-09 0.0028 2.203e-09 0 2.397e-09 0 2.4e-09 0.0028 2.403e-09 0 2.597e-09 0 2.6e-09 0.0028 2.603e-09 0 2.797e-09 0 2.8e-09 0.0028 2.803e-09 0 2.997e-09 0 3e-09 0.0028 3.003e-09 0 3.197e-09 0 3.2e-09 0.0028 3.203e-09 0 3.397e-09 0 3.4e-09 0.0028 3.403e-09 0 3.597e-09 0 3.6e-09 0.0028 3.603e-09 0 3.797e-09 0 3.8e-09 0.0028 3.803e-09 0 3.997e-09 0 4e-09 0.0028 4.003e-09 0 4.197e-09 0 4.2e-09 0.0028 4.203e-09 0 4.397e-09 0 4.4e-09 0.0028 4.403e-09 0 4.597e-09 0 4.6e-09 0.0028 4.603e-09 0 4.797e-09 0 4.8e-09 0.0028 4.803e-09 0 4.997e-09 0 5e-09 0.0028 5.003e-09 0 5.197e-09 0 5.2e-09 0.0028 5.203e-09 0 5.397e-09 0 5.4e-09 0.0028 5.403e-09 0 5.597e-09 0 5.6e-09 0.0028 5.603e-09 0 5.797e-09 0 5.8e-09 0.0028 5.803e-09 0 5.997e-09 0 6e-09 0.0028 6.003e-09 0 6.197e-09 0 6.2e-09 0.0028 6.203e-09 0 6.397e-09 0 6.4e-09 0.0028 6.403e-09 0 6.597e-09 0 6.6e-09 0.0028 6.603e-09 0 6.797e-09 0 6.8e-09 0.0028 6.803e-09 0 6.997e-09 0 7e-09 0.0028 7.003e-09 0 7.197e-09 0 7.2e-09 0.0028 7.203e-09 0 7.397e-09 0 7.4e-09 0.0028 7.403e-09 0 7.597e-09 0 7.6e-09 0.0028 7.603e-09 0 7.797e-09 0 7.8e-09 0.0028 7.803e-09 0 7.997e-09 0 8e-09 0.0028 8.003e-09 0 8.197e-09 0 8.2e-09 0.0028 8.203e-09 0 8.397e-09 0 8.4e-09 0.0028 8.403e-09 0 8.597e-09 0 8.6e-09 0.0028 8.603e-09 0 8.797e-09 0 8.8e-09 0.0028 8.803e-09 0 8.997e-09 0 9e-09 0.0028 9.003e-09 0 9.197e-09 0 9.2e-09 0.0028 9.203e-09 0 9.397e-09 0 9.4e-09 0.0028 9.403e-09 0 9.597e-09 0 9.6e-09 0.0028 9.603e-09 0 9.797e-09 0 9.8e-09 0.0028 9.803e-09 0 9.997e-09 0 1e-08 0.0028 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0028 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0028 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0028 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0028 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0028 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0028 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0028 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0028 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0028 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0028 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0028 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0028 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0028 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0028 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0028 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0028 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0028 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0028 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0028 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0028 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0028 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0028 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0028 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0028 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0028 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0028 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0028 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0028 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0028 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0028 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0028 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0028 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0028 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0028 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0028 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0028 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0028 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0028 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0028 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0028 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0028 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0028 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0028 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0028 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0028 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0028 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0028 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0028 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0028 1.9803e-08 0 1.9997e-08 0 2e-08 0.0028 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0028 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0028 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0028 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0028 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0028 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0028 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0028 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0028 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0028 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0028 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0028 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0028 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0028 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0028 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0028 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0028 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0028 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0028 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0028 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0028 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0028 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0028 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0028 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0028 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0028 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0028 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0028 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0028 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0028 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0028 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0028 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0028 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0028 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0028 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0028 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0028 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0028 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0028 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0028 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0028 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0028 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0028 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0028 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0028 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0028 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0028 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0028 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0028 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0028 2.9803e-08 0 2.9997e-08 0 3e-08 0.0028 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0028 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0028 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0028 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0028 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0028 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0028 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0028 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0028 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0028 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0028 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0028 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0028 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0028 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0028 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0028 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0028 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0028 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0028 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0028 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0028 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0028 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0028 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0028 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0028 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0028 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0028 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0028 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0028 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0028 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0028 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0028 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0028 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0028 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0028 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0028 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0028 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0028 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0028 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0028 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0028 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0028 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0028 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0028 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0028 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0028 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0028 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0028 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0028 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0028 3.9803e-08 0 3.9997e-08 0 4e-08 0.0028 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0028 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0028 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0028 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0028 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0028 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0028 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0028 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0028 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0028 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0028 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0028 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0028 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0028 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0028 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0028 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0028 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0028 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0028 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0028 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0028 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0028 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0028 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0028 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0028 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0028 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0028 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0028 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0028 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0028 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0028 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0028 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0028 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0028 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0028 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0028 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0028 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0028 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0028 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0028 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0028 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0028 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0028 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0028 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0028 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0028 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0028 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0028 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0028 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0028 4.9803e-08 0 4.9997e-08 0 5e-08 0.0028 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0028 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0028 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0028 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0028 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0028 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0028 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0028 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0028 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0028 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0028 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0028 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0028 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0028 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0028 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0028 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0028 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0028 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0028 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0028 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0028 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0028 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0028 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0028 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0028 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0028 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0028 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0028 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0028 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0028 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0028 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0028 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0028 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0028 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0028 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0028 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0028 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0028 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0028 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0028 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0028 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0028 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0028 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0028 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0028 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0028 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0028 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0028 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0028 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0028 5.9803e-08 0 5.9997e-08 0 6e-08 0.0028 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0028 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0028 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0028 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0028 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0028 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0028 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0028 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0028 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0028 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0028 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0028 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0028 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0028 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0028 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0028 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0028 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0028 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0028 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0028 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0028 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0028 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0028 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0028 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0028 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0028 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0028 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0028 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0028 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0028 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0028 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0028 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0028 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0028 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0028 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0028 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0028 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0028 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0028 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0028 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0028 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0028 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0028 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0028 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0028 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0028 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0028 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0028 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0028 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0028 6.9803e-08 0 6.9997e-08 0 7e-08 0.0028 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0028 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0028 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0028 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0028 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0028 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0028 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0028 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0028 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0028 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0028 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0028 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0028 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0028 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0028 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0028 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0028 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0028 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0028 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0028 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0028 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0028 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0028 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0028 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0028 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0028 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0028 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0028 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0028 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0028 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0028 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0028 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0028 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0028 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0028 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0028 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0028 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0028 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0028 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0028 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0028 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0028 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0028 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0028 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0028 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0028 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0028 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0028 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0028 7.9603e-08 0)
IT48|T 0 T48  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_IP7_34|1 IP7_3_OUT _IP7_34|A1  2.067833848e-12
L_IP7_34|2 _IP7_34|A1 _IP7_34|A2  4.135667696e-12
L_IP7_34|3 _IP7_34|A3 _IP7_34|A4  8.271335392e-12
L_IP7_34|T T48 _IP7_34|T1  2.067833848e-12
L_IP7_34|4 _IP7_34|T1 _IP7_34|T2  4.135667696e-12
L_IP7_34|5 _IP7_34|A4 _IP7_34|Q1  4.135667696e-12
L_IP7_34|6 _IP7_34|Q1 IP7_4_OUT_TX  2.067833848e-12
IT49|T 0 T49  PWL(0 0 -3e-12 0 0 0.0007 3e-12 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9997e-08 0 4e-08 0.0007 4.0003e-08 0 4.0197e-08 0 4.02e-08 0.0007 4.0203e-08 0 4.0397e-08 0 4.04e-08 0.0007 4.0403e-08 0 4.0597e-08 0 4.06e-08 0.0007 4.0603e-08 0 4.0797e-08 0 4.08e-08 0.0007 4.0803e-08 0 4.0997e-08 0 4.1e-08 0.0007 4.1003e-08 0 4.1197e-08 0 4.12e-08 0.0007 4.1203e-08 0 4.1397e-08 0 4.14e-08 0.0007 4.1403e-08 0 4.1597e-08 0 4.16e-08 0.0007 4.1603e-08 0 4.1797e-08 0 4.18e-08 0.0007 4.1803e-08 0 4.1997e-08 0 4.2e-08 0.0007 4.2003e-08 0 4.2197e-08 0 4.22e-08 0.0007 4.2203e-08 0 4.2397e-08 0 4.24e-08 0.0007 4.2403e-08 0 4.2597e-08 0 4.26e-08 0.0007 4.2603e-08 0 4.2797e-08 0 4.28e-08 0.0007 4.2803e-08 0 4.2997e-08 0 4.3e-08 0.0007 4.3003e-08 0 4.3197e-08 0 4.32e-08 0.0007 4.3203e-08 0 4.3397e-08 0 4.34e-08 0.0007 4.3403e-08 0 4.3597e-08 0 4.36e-08 0.0007 4.3603e-08 0 4.3797e-08 0 4.38e-08 0.0007 4.3803e-08 0 4.3997e-08 0 4.4e-08 0.0007 4.4003e-08 0 4.4197e-08 0 4.42e-08 0.0007 4.4203e-08 0 4.4397e-08 0 4.44e-08 0.0007 4.4403e-08 0 4.4597e-08 0 4.46e-08 0.0007 4.4603e-08 0 4.4797e-08 0 4.48e-08 0.0007 4.4803e-08 0 4.4997e-08 0 4.5e-08 0.0007 4.5003e-08 0 4.5197e-08 0 4.52e-08 0.0007 4.5203e-08 0 4.5397e-08 0 4.54e-08 0.0007 4.5403e-08 0 4.5597e-08 0 4.56e-08 0.0007 4.5603e-08 0 4.5797e-08 0 4.58e-08 0.0007 4.5803e-08 0 4.5997e-08 0 4.6e-08 0.0007 4.6003e-08 0 4.6197e-08 0 4.62e-08 0.0007 4.6203e-08 0 4.6397e-08 0 4.64e-08 0.0007 4.6403e-08 0 4.6597e-08 0 4.66e-08 0.0007 4.6603e-08 0 4.6797e-08 0 4.68e-08 0.0007 4.6803e-08 0 4.6997e-08 0 4.7e-08 0.0007 4.7003e-08 0 4.7197e-08 0 4.72e-08 0.0007 4.7203e-08 0 4.7397e-08 0 4.74e-08 0.0007 4.7403e-08 0 4.7597e-08 0 4.76e-08 0.0007 4.7603e-08 0 4.7797e-08 0 4.78e-08 0.0007 4.7803e-08 0 4.7997e-08 0 4.8e-08 0.0007 4.8003e-08 0 4.8197e-08 0 4.82e-08 0.0007 4.8203e-08 0 4.8397e-08 0 4.84e-08 0.0007 4.8403e-08 0 4.8597e-08 0 4.86e-08 0.0007 4.8603e-08 0 4.8797e-08 0 4.88e-08 0.0007 4.8803e-08 0 4.8997e-08 0 4.9e-08 0.0007 4.9003e-08 0 4.9197e-08 0 4.92e-08 0.0007 4.9203e-08 0 4.9397e-08 0 4.94e-08 0.0007 4.9403e-08 0 4.9597e-08 0 4.96e-08 0.0007 4.9603e-08 0 4.9797e-08 0 4.98e-08 0.0007 4.9803e-08 0 4.9997e-08 0 5e-08 0.0007 5.0003e-08 0 5.0197e-08 0 5.02e-08 0.0007 5.0203e-08 0 5.0397e-08 0 5.04e-08 0.0007 5.0403e-08 0 5.0597e-08 0 5.06e-08 0.0007 5.0603e-08 0 5.0797e-08 0 5.08e-08 0.0007 5.0803e-08 0 5.0997e-08 0 5.1e-08 0.0007 5.1003e-08 0 5.1197e-08 0 5.12e-08 0.0007 5.1203e-08 0 5.1397e-08 0 5.14e-08 0.0007 5.1403e-08 0 5.1597e-08 0 5.16e-08 0.0007 5.1603e-08 0 5.1797e-08 0 5.18e-08 0.0007 5.1803e-08 0 5.1997e-08 0 5.2e-08 0.0007 5.2003e-08 0 5.2197e-08 0 5.22e-08 0.0007 5.2203e-08 0 5.2397e-08 0 5.24e-08 0.0007 5.2403e-08 0 5.2597e-08 0 5.26e-08 0.0007 5.2603e-08 0 5.2797e-08 0 5.28e-08 0.0007 5.2803e-08 0 5.2997e-08 0 5.3e-08 0.0007 5.3003e-08 0 5.3197e-08 0 5.32e-08 0.0007 5.3203e-08 0 5.3397e-08 0 5.34e-08 0.0007 5.3403e-08 0 5.3597e-08 0 5.36e-08 0.0007 5.3603e-08 0 5.3797e-08 0 5.38e-08 0.0007 5.3803e-08 0 5.3997e-08 0 5.4e-08 0.0007 5.4003e-08 0 5.4197e-08 0 5.42e-08 0.0007 5.4203e-08 0 5.4397e-08 0 5.44e-08 0.0007 5.4403e-08 0 5.4597e-08 0 5.46e-08 0.0007 5.4603e-08 0 5.4797e-08 0 5.48e-08 0.0007 5.4803e-08 0 5.4997e-08 0 5.5e-08 0.0007 5.5003e-08 0 5.5197e-08 0 5.52e-08 0.0007 5.5203e-08 0 5.5397e-08 0 5.54e-08 0.0007 5.5403e-08 0 5.5597e-08 0 5.56e-08 0.0007 5.5603e-08 0 5.5797e-08 0 5.58e-08 0.0007 5.5803e-08 0 5.5997e-08 0 5.6e-08 0.0007 5.6003e-08 0 5.6197e-08 0 5.62e-08 0.0007 5.6203e-08 0 5.6397e-08 0 5.64e-08 0.0007 5.6403e-08 0 5.6597e-08 0 5.66e-08 0.0007 5.6603e-08 0 5.6797e-08 0 5.68e-08 0.0007 5.6803e-08 0 5.6997e-08 0 5.7e-08 0.0007 5.7003e-08 0 5.7197e-08 0 5.72e-08 0.0007 5.7203e-08 0 5.7397e-08 0 5.74e-08 0.0007 5.7403e-08 0 5.7597e-08 0 5.76e-08 0.0007 5.7603e-08 0 5.7797e-08 0 5.78e-08 0.0007 5.7803e-08 0 5.7997e-08 0 5.8e-08 0.0007 5.8003e-08 0 5.8197e-08 0 5.82e-08 0.0007 5.8203e-08 0 5.8397e-08 0 5.84e-08 0.0007 5.8403e-08 0 5.8597e-08 0 5.86e-08 0.0007 5.8603e-08 0 5.8797e-08 0 5.88e-08 0.0007 5.8803e-08 0 5.8997e-08 0 5.9e-08 0.0007 5.9003e-08 0 5.9197e-08 0 5.92e-08 0.0007 5.9203e-08 0 5.9397e-08 0 5.94e-08 0.0007 5.9403e-08 0 5.9597e-08 0 5.96e-08 0.0007 5.9603e-08 0 5.9797e-08 0 5.98e-08 0.0007 5.9803e-08 0 5.9997e-08 0 6e-08 0.0007 6.0003e-08 0 6.0197e-08 0 6.02e-08 0.0007 6.0203e-08 0 6.0397e-08 0 6.04e-08 0.0007 6.0403e-08 0 6.0597e-08 0 6.06e-08 0.0007 6.0603e-08 0 6.0797e-08 0 6.08e-08 0.0007 6.0803e-08 0 6.0997e-08 0 6.1e-08 0.0007 6.1003e-08 0 6.1197e-08 0 6.12e-08 0.0007 6.1203e-08 0 6.1397e-08 0 6.14e-08 0.0007 6.1403e-08 0 6.1597e-08 0 6.16e-08 0.0007 6.1603e-08 0 6.1797e-08 0 6.18e-08 0.0007 6.1803e-08 0 6.1997e-08 0 6.2e-08 0.0007 6.2003e-08 0 6.2197e-08 0 6.22e-08 0.0007 6.2203e-08 0 6.2397e-08 0 6.24e-08 0.0007 6.2403e-08 0 6.2597e-08 0 6.26e-08 0.0007 6.2603e-08 0 6.2797e-08 0 6.28e-08 0.0007 6.2803e-08 0 6.2997e-08 0 6.3e-08 0.0007 6.3003e-08 0 6.3197e-08 0 6.32e-08 0.0007 6.3203e-08 0 6.3397e-08 0 6.34e-08 0.0007 6.3403e-08 0 6.3597e-08 0 6.36e-08 0.0007 6.3603e-08 0 6.3797e-08 0 6.38e-08 0.0007 6.3803e-08 0 6.3997e-08 0 6.4e-08 0.0007 6.4003e-08 0 6.4197e-08 0 6.42e-08 0.0007 6.4203e-08 0 6.4397e-08 0 6.44e-08 0.0007 6.4403e-08 0 6.4597e-08 0 6.46e-08 0.0007 6.4603e-08 0 6.4797e-08 0 6.48e-08 0.0007 6.4803e-08 0 6.4997e-08 0 6.5e-08 0.0007 6.5003e-08 0 6.5197e-08 0 6.52e-08 0.0007 6.5203e-08 0 6.5397e-08 0 6.54e-08 0.0007 6.5403e-08 0 6.5597e-08 0 6.56e-08 0.0007 6.5603e-08 0 6.5797e-08 0 6.58e-08 0.0007 6.5803e-08 0 6.5997e-08 0 6.6e-08 0.0007 6.6003e-08 0 6.6197e-08 0 6.62e-08 0.0007 6.6203e-08 0 6.6397e-08 0 6.64e-08 0.0007 6.6403e-08 0 6.6597e-08 0 6.66e-08 0.0007 6.6603e-08 0 6.6797e-08 0 6.68e-08 0.0007 6.6803e-08 0 6.6997e-08 0 6.7e-08 0.0007 6.7003e-08 0 6.7197e-08 0 6.72e-08 0.0007 6.7203e-08 0 6.7397e-08 0 6.74e-08 0.0007 6.7403e-08 0 6.7597e-08 0 6.76e-08 0.0007 6.7603e-08 0 6.7797e-08 0 6.78e-08 0.0007 6.7803e-08 0 6.7997e-08 0 6.8e-08 0.0007 6.8003e-08 0 6.8197e-08 0 6.82e-08 0.0007 6.8203e-08 0 6.8397e-08 0 6.84e-08 0.0007 6.8403e-08 0 6.8597e-08 0 6.86e-08 0.0007 6.8603e-08 0 6.8797e-08 0 6.88e-08 0.0007 6.8803e-08 0 6.8997e-08 0 6.9e-08 0.0007 6.9003e-08 0 6.9197e-08 0 6.92e-08 0.0007 6.9203e-08 0 6.9397e-08 0 6.94e-08 0.0007 6.9403e-08 0 6.9597e-08 0 6.96e-08 0.0007 6.9603e-08 0 6.9797e-08 0 6.98e-08 0.0007 6.9803e-08 0 6.9997e-08 0 7e-08 0.0007 7.0003e-08 0 7.0197e-08 0 7.02e-08 0.0007 7.0203e-08 0 7.0397e-08 0 7.04e-08 0.0007 7.0403e-08 0 7.0597e-08 0 7.06e-08 0.0007 7.0603e-08 0 7.0797e-08 0 7.08e-08 0.0007 7.0803e-08 0 7.0997e-08 0 7.1e-08 0.0007 7.1003e-08 0 7.1197e-08 0 7.12e-08 0.0007 7.1203e-08 0 7.1397e-08 0 7.14e-08 0.0007 7.1403e-08 0 7.1597e-08 0 7.16e-08 0.0007 7.1603e-08 0 7.1797e-08 0 7.18e-08 0.0007 7.1803e-08 0 7.1997e-08 0 7.2e-08 0.0007 7.2003e-08 0 7.2197e-08 0 7.22e-08 0.0007 7.2203e-08 0 7.2397e-08 0 7.24e-08 0.0007 7.2403e-08 0 7.2597e-08 0 7.26e-08 0.0007 7.2603e-08 0 7.2797e-08 0 7.28e-08 0.0007 7.2803e-08 0 7.2997e-08 0 7.3e-08 0.0007 7.3003e-08 0 7.3197e-08 0 7.32e-08 0.0007 7.3203e-08 0 7.3397e-08 0 7.34e-08 0.0007 7.3403e-08 0 7.3597e-08 0 7.36e-08 0.0007 7.3603e-08 0 7.3797e-08 0 7.38e-08 0.0007 7.3803e-08 0 7.3997e-08 0 7.4e-08 0.0007 7.4003e-08 0 7.4197e-08 0 7.42e-08 0.0007 7.4203e-08 0 7.4397e-08 0 7.44e-08 0.0007 7.4403e-08 0 7.4597e-08 0 7.46e-08 0.0007 7.4603e-08 0 7.4797e-08 0 7.48e-08 0.0007 7.4803e-08 0 7.4997e-08 0 7.5e-08 0.0007 7.5003e-08 0 7.5197e-08 0 7.52e-08 0.0007 7.5203e-08 0 7.5397e-08 0 7.54e-08 0.0007 7.5403e-08 0 7.5597e-08 0 7.56e-08 0.0007 7.5603e-08 0 7.5797e-08 0 7.58e-08 0.0007 7.5803e-08 0 7.5997e-08 0 7.6e-08 0.0007 7.6003e-08 0 7.6197e-08 0 7.62e-08 0.0007 7.6203e-08 0 7.6397e-08 0 7.64e-08 0.0007 7.6403e-08 0 7.6597e-08 0 7.66e-08 0.0007 7.6603e-08 0 7.6797e-08 0 7.68e-08 0.0007 7.6803e-08 0 7.6997e-08 0 7.7e-08 0.0007 7.7003e-08 0 7.7197e-08 0 7.72e-08 0.0007 7.7203e-08 0 7.7397e-08 0 7.74e-08 0.0007 7.7403e-08 0 7.7597e-08 0 7.76e-08 0.0007 7.7603e-08 0 7.7797e-08 0 7.78e-08 0.0007 7.7803e-08 0 7.7997e-08 0 7.8e-08 0.0007 7.8003e-08 0 7.8197e-08 0 7.82e-08 0.0007 7.8203e-08 0 7.8397e-08 0 7.84e-08 0.0007 7.8403e-08 0 7.8597e-08 0 7.86e-08 0.0007 7.8603e-08 0 7.8797e-08 0 7.88e-08 0.0007 7.8803e-08 0 7.8997e-08 0 7.9e-08 0.0007 7.9003e-08 0 7.9197e-08 0 7.92e-08 0.0007 7.9203e-08 0 7.9397e-08 0 7.94e-08 0.0007 7.9403e-08 0 7.9597e-08 0 7.96e-08 0.0007 7.9603e-08 0)
L_S8_34|1 S8_3 _S8_34|A1  2.067833848e-12
L_S8_34|2 _S8_34|A1 _S8_34|A2  4.135667696e-12
L_S8_34|3 _S8_34|A3 _S8_34|A4  8.271335392e-12
L_S8_34|T T49 _S8_34|T1  2.067833848e-12
L_S8_34|4 _S8_34|T1 _S8_34|T2  4.135667696e-12
L_S8_34|5 _S8_34|A4 _S8_34|Q1  4.135667696e-12
L_S8_34|6 _S8_34|Q1 S8_4_TX  2.067833848e-12
IT50|T 0 T50  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S0_45|1 S0_4 _S0_45|A1  2.067833848e-12
L_S0_45|2 _S0_45|A1 _S0_45|A2  4.135667696e-12
L_S0_45|3 _S0_45|A3 _S0_45|A4  8.271335392e-12
L_S0_45|T T50 _S0_45|T1  2.067833848e-12
L_S0_45|4 _S0_45|T1 _S0_45|T2  4.135667696e-12
L_S0_45|5 _S0_45|A4 _S0_45|Q1  4.135667696e-12
L_S0_45|6 _S0_45|Q1 S0_5_TX  2.067833848e-12
IT51|T 0 T51  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S1_45|1 S1_4 _S1_45|A1  2.067833848e-12
L_S1_45|2 _S1_45|A1 _S1_45|A2  4.135667696e-12
L_S1_45|3 _S1_45|A3 _S1_45|A4  8.271335392e-12
L_S1_45|T T51 _S1_45|T1  2.067833848e-12
L_S1_45|4 _S1_45|T1 _S1_45|T2  4.135667696e-12
L_S1_45|5 _S1_45|A4 _S1_45|Q1  4.135667696e-12
L_S1_45|6 _S1_45|Q1 S1_5_TX  2.067833848e-12
IT52|T 0 T52  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S2_45|1 S2_4 _S2_45|A1  2.067833848e-12
L_S2_45|2 _S2_45|A1 _S2_45|A2  4.135667696e-12
L_S2_45|3 _S2_45|A3 _S2_45|A4  8.271335392e-12
L_S2_45|T T52 _S2_45|T1  2.067833848e-12
L_S2_45|4 _S2_45|T1 _S2_45|T2  4.135667696e-12
L_S2_45|5 _S2_45|A4 _S2_45|Q1  4.135667696e-12
L_S2_45|6 _S2_45|Q1 S2_5_TX  2.067833848e-12
IT53|T 0 T53  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S3_45|1 S3_4 _S3_45|A1  2.067833848e-12
L_S3_45|2 _S3_45|A1 _S3_45|A2  4.135667696e-12
L_S3_45|3 _S3_45|A3 _S3_45|A4  8.271335392e-12
L_S3_45|T T53 _S3_45|T1  2.067833848e-12
L_S3_45|4 _S3_45|T1 _S3_45|T2  4.135667696e-12
L_S3_45|5 _S3_45|A4 _S3_45|Q1  4.135667696e-12
L_S3_45|6 _S3_45|Q1 S3_5_TX  2.067833848e-12
IT54|T 0 T54  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S4_45|1 S4_4 _S4_45|A1  2.067833848e-12
L_S4_45|2 _S4_45|A1 _S4_45|A2  4.135667696e-12
L_S4_45|3 _S4_45|A3 _S4_45|A4  8.271335392e-12
L_S4_45|T T54 _S4_45|T1  2.067833848e-12
L_S4_45|4 _S4_45|T1 _S4_45|T2  4.135667696e-12
L_S4_45|5 _S4_45|A4 _S4_45|Q1  4.135667696e-12
L_S4_45|6 _S4_45|Q1 S4_5_TX  2.067833848e-12
IT55|T 0 T55  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S5_45|1 S5_4 _S5_45|A1  2.067833848e-12
L_S5_45|2 _S5_45|A1 _S5_45|A2  4.135667696e-12
L_S5_45|3 _S5_45|A3 _S5_45|A4  8.271335392e-12
L_S5_45|T T55 _S5_45|T1  2.067833848e-12
L_S5_45|4 _S5_45|T1 _S5_45|T2  4.135667696e-12
L_S5_45|5 _S5_45|A4 _S5_45|Q1  4.135667696e-12
L_S5_45|6 _S5_45|Q1 S5_5_TX  2.067833848e-12
IT56|T 0 T56  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S6_45|1 S6_4 _S6_45|A1  2.067833848e-12
L_S6_45|2 _S6_45|A1 _S6_45|A2  4.135667696e-12
L_S6_45|3 _S6_45|A3 _S6_45|A4  8.271335392e-12
L_S6_45|T T56 _S6_45|T1  2.067833848e-12
L_S6_45|4 _S6_45|T1 _S6_45|T2  4.135667696e-12
L_S6_45|5 _S6_45|A4 _S6_45|Q1  4.135667696e-12
L_S6_45|6 _S6_45|Q1 S6_5_TX  2.067833848e-12
IT57|T 0 T57  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S7_45|A1 G6_4_OUT _S7_45|A1  2.067833848e-12
L_S7_45|A2 _S7_45|A1 _S7_45|A2  4.135667696e-12
L_S7_45|A3 _S7_45|A3 _S7_45|AB  8.271335392e-12
L_S7_45|B1 IP7_4_OUT _S7_45|B1  2.067833848e-12
L_S7_45|B2 _S7_45|B1 _S7_45|B2  4.135667696e-12
L_S7_45|B3 _S7_45|B3 _S7_45|AB  8.271335392e-12
L_S7_45|T1 T57 _S7_45|T1  2.067833848e-12
L_S7_45|T2 _S7_45|T1 _S7_45|T2  4.135667696e-12
L_S7_45|Q2 _S7_45|ABTQ _S7_45|Q1  4.135667696e-12
L_S7_45|Q1 _S7_45|Q1 S7_4_TX  2.067833848e-12
IT58|T 0 T58  PWL(0 0 -1.3e-11 0 -1e-11 0.0007 -7e-12 0 1.87e-10 0 1.9e-10 0.0007 1.93e-10 0 3.87e-10 0 3.9e-10 0.0007 3.93e-10 0 5.87e-10 0 5.9e-10 0.0007 5.93e-10 0 7.87e-10 0 7.9e-10 0.0007 7.93e-10 0 9.87e-10 0 9.9e-10 0.0007 9.93e-10 0 1.187e-09 0 1.19e-09 0.0007 1.193e-09 0 1.387e-09 0 1.39e-09 0.0007 1.393e-09 0 1.587e-09 0 1.59e-09 0.0007 1.593e-09 0 1.787e-09 0 1.79e-09 0.0007 1.793e-09 0 1.987e-09 0 1.99e-09 0.0007 1.993e-09 0 2.187e-09 0 2.19e-09 0.0007 2.193e-09 0 2.387e-09 0 2.39e-09 0.0007 2.393e-09 0 2.587e-09 0 2.59e-09 0.0007 2.593e-09 0 2.787e-09 0 2.79e-09 0.0007 2.793e-09 0 2.987e-09 0 2.99e-09 0.0007 2.993e-09 0 3.187e-09 0 3.19e-09 0.0007 3.193e-09 0 3.387e-09 0 3.39e-09 0.0007 3.393e-09 0 3.587e-09 0 3.59e-09 0.0007 3.593e-09 0 3.787e-09 0 3.79e-09 0.0007 3.793e-09 0 3.987e-09 0 3.99e-09 0.0007 3.993e-09 0 4.187e-09 0 4.19e-09 0.0007 4.193e-09 0 4.387e-09 0 4.39e-09 0.0007 4.393e-09 0 4.587e-09 0 4.59e-09 0.0007 4.593e-09 0 4.787e-09 0 4.79e-09 0.0007 4.793e-09 0 4.987e-09 0 4.99e-09 0.0007 4.993e-09 0 5.187e-09 0 5.19e-09 0.0007 5.193e-09 0 5.387e-09 0 5.39e-09 0.0007 5.393e-09 0 5.587e-09 0 5.59e-09 0.0007 5.593e-09 0 5.787e-09 0 5.79e-09 0.0007 5.793e-09 0 5.987e-09 0 5.99e-09 0.0007 5.993e-09 0 6.187e-09 0 6.19e-09 0.0007 6.193e-09 0 6.387e-09 0 6.39e-09 0.0007 6.393e-09 0 6.587e-09 0 6.59e-09 0.0007 6.593e-09 0 6.787e-09 0 6.79e-09 0.0007 6.793e-09 0 6.987e-09 0 6.99e-09 0.0007 6.993e-09 0 7.187e-09 0 7.19e-09 0.0007 7.193e-09 0 7.387e-09 0 7.39e-09 0.0007 7.393e-09 0 7.587e-09 0 7.59e-09 0.0007 7.593e-09 0 7.787e-09 0 7.79e-09 0.0007 7.793e-09 0 7.987e-09 0 7.99e-09 0.0007 7.993e-09 0 8.187e-09 0 8.19e-09 0.0007 8.193e-09 0 8.387e-09 0 8.39e-09 0.0007 8.393e-09 0 8.587e-09 0 8.59e-09 0.0007 8.593e-09 0 8.787e-09 0 8.79e-09 0.0007 8.793e-09 0 8.987e-09 0 8.99e-09 0.0007 8.993e-09 0 9.187e-09 0 9.19e-09 0.0007 9.193e-09 0 9.387e-09 0 9.39e-09 0.0007 9.393e-09 0 9.587e-09 0 9.59e-09 0.0007 9.593e-09 0 9.787e-09 0 9.79e-09 0.0007 9.793e-09 0 9.987e-09 0 9.99e-09 0.0007 9.993e-09 0 1.0187e-08 0 1.019e-08 0.0007 1.0193e-08 0 1.0387e-08 0 1.039e-08 0.0007 1.0393e-08 0 1.0587e-08 0 1.059e-08 0.0007 1.0593e-08 0 1.0787e-08 0 1.079e-08 0.0007 1.0793e-08 0 1.0987e-08 0 1.099e-08 0.0007 1.0993e-08 0 1.1187e-08 0 1.119e-08 0.0007 1.1193e-08 0 1.1387e-08 0 1.139e-08 0.0007 1.1393e-08 0 1.1587e-08 0 1.159e-08 0.0007 1.1593e-08 0 1.1787e-08 0 1.179e-08 0.0007 1.1793e-08 0 1.1987e-08 0 1.199e-08 0.0007 1.1993e-08 0 1.2187e-08 0 1.219e-08 0.0007 1.2193e-08 0 1.2387e-08 0 1.239e-08 0.0007 1.2393e-08 0 1.2587e-08 0 1.259e-08 0.0007 1.2593e-08 0 1.2787e-08 0 1.279e-08 0.0007 1.2793e-08 0 1.2987e-08 0 1.299e-08 0.0007 1.2993e-08 0 1.3187e-08 0 1.319e-08 0.0007 1.3193e-08 0 1.3387e-08 0 1.339e-08 0.0007 1.3393e-08 0 1.3587e-08 0 1.359e-08 0.0007 1.3593e-08 0 1.3787e-08 0 1.379e-08 0.0007 1.3793e-08 0 1.3987e-08 0 1.399e-08 0.0007 1.3993e-08 0 1.4187e-08 0 1.419e-08 0.0007 1.4193e-08 0 1.4387e-08 0 1.439e-08 0.0007 1.4393e-08 0 1.4587e-08 0 1.459e-08 0.0007 1.4593e-08 0 1.4787e-08 0 1.479e-08 0.0007 1.4793e-08 0 1.4987e-08 0 1.499e-08 0.0007 1.4993e-08 0 1.5187e-08 0 1.519e-08 0.0007 1.5193e-08 0 1.5387e-08 0 1.539e-08 0.0007 1.5393e-08 0 1.5587e-08 0 1.559e-08 0.0007 1.5593e-08 0 1.5787e-08 0 1.579e-08 0.0007 1.5793e-08 0 1.5987e-08 0 1.599e-08 0.0007 1.5993e-08 0 1.6187e-08 0 1.619e-08 0.0007 1.6193e-08 0 1.6387e-08 0 1.639e-08 0.0007 1.6393e-08 0 1.6587e-08 0 1.659e-08 0.0007 1.6593e-08 0 1.6787e-08 0 1.679e-08 0.0007 1.6793e-08 0 1.6987e-08 0 1.699e-08 0.0007 1.6993e-08 0 1.7187e-08 0 1.719e-08 0.0007 1.7193e-08 0 1.7387e-08 0 1.739e-08 0.0007 1.7393e-08 0 1.7587e-08 0 1.759e-08 0.0007 1.7593e-08 0 1.7787e-08 0 1.779e-08 0.0007 1.7793e-08 0 1.7987e-08 0 1.799e-08 0.0007 1.7993e-08 0 1.8187e-08 0 1.819e-08 0.0007 1.8193e-08 0 1.8387e-08 0 1.839e-08 0.0007 1.8393e-08 0 1.8587e-08 0 1.859e-08 0.0007 1.8593e-08 0 1.8787e-08 0 1.879e-08 0.0007 1.8793e-08 0 1.8987e-08 0 1.899e-08 0.0007 1.8993e-08 0 1.9187e-08 0 1.919e-08 0.0007 1.9193e-08 0 1.9387e-08 0 1.939e-08 0.0007 1.9393e-08 0 1.9587e-08 0 1.959e-08 0.0007 1.9593e-08 0 1.9787e-08 0 1.979e-08 0.0007 1.9793e-08 0 1.9987e-08 0 1.999e-08 0.0007 1.9993e-08 0 2.0187e-08 0 2.019e-08 0.0007 2.0193e-08 0 2.0387e-08 0 2.039e-08 0.0007 2.0393e-08 0 2.0587e-08 0 2.059e-08 0.0007 2.0593e-08 0 2.0787e-08 0 2.079e-08 0.0007 2.0793e-08 0 2.0987e-08 0 2.099e-08 0.0007 2.0993e-08 0 2.1187e-08 0 2.119e-08 0.0007 2.1193e-08 0 2.1387e-08 0 2.139e-08 0.0007 2.1393e-08 0 2.1587e-08 0 2.159e-08 0.0007 2.1593e-08 0 2.1787e-08 0 2.179e-08 0.0007 2.1793e-08 0 2.1987e-08 0 2.199e-08 0.0007 2.1993e-08 0 2.2187e-08 0 2.219e-08 0.0007 2.2193e-08 0 2.2387e-08 0 2.239e-08 0.0007 2.2393e-08 0 2.2587e-08 0 2.259e-08 0.0007 2.2593e-08 0 2.2787e-08 0 2.279e-08 0.0007 2.2793e-08 0 2.2987e-08 0 2.299e-08 0.0007 2.2993e-08 0 2.3187e-08 0 2.319e-08 0.0007 2.3193e-08 0 2.3387e-08 0 2.339e-08 0.0007 2.3393e-08 0 2.3587e-08 0 2.359e-08 0.0007 2.3593e-08 0 2.3787e-08 0 2.379e-08 0.0007 2.3793e-08 0 2.3987e-08 0 2.399e-08 0.0007 2.3993e-08 0 2.4187e-08 0 2.419e-08 0.0007 2.4193e-08 0 2.4387e-08 0 2.439e-08 0.0007 2.4393e-08 0 2.4587e-08 0 2.459e-08 0.0007 2.4593e-08 0 2.4787e-08 0 2.479e-08 0.0007 2.4793e-08 0 2.4987e-08 0 2.499e-08 0.0007 2.4993e-08 0 2.5187e-08 0 2.519e-08 0.0007 2.5193e-08 0 2.5387e-08 0 2.539e-08 0.0007 2.5393e-08 0 2.5587e-08 0 2.559e-08 0.0007 2.5593e-08 0 2.5787e-08 0 2.579e-08 0.0007 2.5793e-08 0 2.5987e-08 0 2.599e-08 0.0007 2.5993e-08 0 2.6187e-08 0 2.619e-08 0.0007 2.6193e-08 0 2.6387e-08 0 2.639e-08 0.0007 2.6393e-08 0 2.6587e-08 0 2.659e-08 0.0007 2.6593e-08 0 2.6787e-08 0 2.679e-08 0.0007 2.6793e-08 0 2.6987e-08 0 2.699e-08 0.0007 2.6993e-08 0 2.7187e-08 0 2.719e-08 0.0007 2.7193e-08 0 2.7387e-08 0 2.739e-08 0.0007 2.7393e-08 0 2.7587e-08 0 2.759e-08 0.0007 2.7593e-08 0 2.7787e-08 0 2.779e-08 0.0007 2.7793e-08 0 2.7987e-08 0 2.799e-08 0.0007 2.7993e-08 0 2.8187e-08 0 2.819e-08 0.0007 2.8193e-08 0 2.8387e-08 0 2.839e-08 0.0007 2.8393e-08 0 2.8587e-08 0 2.859e-08 0.0007 2.8593e-08 0 2.8787e-08 0 2.879e-08 0.0007 2.8793e-08 0 2.8987e-08 0 2.899e-08 0.0007 2.8993e-08 0 2.9187e-08 0 2.919e-08 0.0007 2.9193e-08 0 2.9387e-08 0 2.939e-08 0.0007 2.9393e-08 0 2.9587e-08 0 2.959e-08 0.0007 2.9593e-08 0 2.9787e-08 0 2.979e-08 0.0007 2.9793e-08 0 2.9987e-08 0 2.999e-08 0.0007 2.9993e-08 0 3.0187e-08 0 3.019e-08 0.0007 3.0193e-08 0 3.0387e-08 0 3.039e-08 0.0007 3.0393e-08 0 3.0587e-08 0 3.059e-08 0.0007 3.0593e-08 0 3.0787e-08 0 3.079e-08 0.0007 3.0793e-08 0 3.0987e-08 0 3.099e-08 0.0007 3.0993e-08 0 3.1187e-08 0 3.119e-08 0.0007 3.1193e-08 0 3.1387e-08 0 3.139e-08 0.0007 3.1393e-08 0 3.1587e-08 0 3.159e-08 0.0007 3.1593e-08 0 3.1787e-08 0 3.179e-08 0.0007 3.1793e-08 0 3.1987e-08 0 3.199e-08 0.0007 3.1993e-08 0 3.2187e-08 0 3.219e-08 0.0007 3.2193e-08 0 3.2387e-08 0 3.239e-08 0.0007 3.2393e-08 0 3.2587e-08 0 3.259e-08 0.0007 3.2593e-08 0 3.2787e-08 0 3.279e-08 0.0007 3.2793e-08 0 3.2987e-08 0 3.299e-08 0.0007 3.2993e-08 0 3.3187e-08 0 3.319e-08 0.0007 3.3193e-08 0 3.3387e-08 0 3.339e-08 0.0007 3.3393e-08 0 3.3587e-08 0 3.359e-08 0.0007 3.3593e-08 0 3.3787e-08 0 3.379e-08 0.0007 3.3793e-08 0 3.3987e-08 0 3.399e-08 0.0007 3.3993e-08 0 3.4187e-08 0 3.419e-08 0.0007 3.4193e-08 0 3.4387e-08 0 3.439e-08 0.0007 3.4393e-08 0 3.4587e-08 0 3.459e-08 0.0007 3.4593e-08 0 3.4787e-08 0 3.479e-08 0.0007 3.4793e-08 0 3.4987e-08 0 3.499e-08 0.0007 3.4993e-08 0 3.5187e-08 0 3.519e-08 0.0007 3.5193e-08 0 3.5387e-08 0 3.539e-08 0.0007 3.5393e-08 0 3.5587e-08 0 3.559e-08 0.0007 3.5593e-08 0 3.5787e-08 0 3.579e-08 0.0007 3.5793e-08 0 3.5987e-08 0 3.599e-08 0.0007 3.5993e-08 0 3.6187e-08 0 3.619e-08 0.0007 3.6193e-08 0 3.6387e-08 0 3.639e-08 0.0007 3.6393e-08 0 3.6587e-08 0 3.659e-08 0.0007 3.6593e-08 0 3.6787e-08 0 3.679e-08 0.0007 3.6793e-08 0 3.6987e-08 0 3.699e-08 0.0007 3.6993e-08 0 3.7187e-08 0 3.719e-08 0.0007 3.7193e-08 0 3.7387e-08 0 3.739e-08 0.0007 3.7393e-08 0 3.7587e-08 0 3.759e-08 0.0007 3.7593e-08 0 3.7787e-08 0 3.779e-08 0.0007 3.7793e-08 0 3.7987e-08 0 3.799e-08 0.0007 3.7993e-08 0 3.8187e-08 0 3.819e-08 0.0007 3.8193e-08 0 3.8387e-08 0 3.839e-08 0.0007 3.8393e-08 0 3.8587e-08 0 3.859e-08 0.0007 3.8593e-08 0 3.8787e-08 0 3.879e-08 0.0007 3.8793e-08 0 3.8987e-08 0 3.899e-08 0.0007 3.8993e-08 0 3.9187e-08 0 3.919e-08 0.0007 3.9193e-08 0 3.9387e-08 0 3.939e-08 0.0007 3.9393e-08 0 3.9587e-08 0 3.959e-08 0.0007 3.9593e-08 0 3.9787e-08 0 3.979e-08 0.0007 3.9793e-08 0 3.9987e-08 0 3.999e-08 0.0007 3.9993e-08 0 4.0187e-08 0 4.019e-08 0.0007 4.0193e-08 0 4.0387e-08 0 4.039e-08 0.0007 4.0393e-08 0 4.0587e-08 0 4.059e-08 0.0007 4.0593e-08 0 4.0787e-08 0 4.079e-08 0.0007 4.0793e-08 0 4.0987e-08 0 4.099e-08 0.0007 4.0993e-08 0 4.1187e-08 0 4.119e-08 0.0007 4.1193e-08 0 4.1387e-08 0 4.139e-08 0.0007 4.1393e-08 0 4.1587e-08 0 4.159e-08 0.0007 4.1593e-08 0 4.1787e-08 0 4.179e-08 0.0007 4.1793e-08 0 4.1987e-08 0 4.199e-08 0.0007 4.1993e-08 0 4.2187e-08 0 4.219e-08 0.0007 4.2193e-08 0 4.2387e-08 0 4.239e-08 0.0007 4.2393e-08 0 4.2587e-08 0 4.259e-08 0.0007 4.2593e-08 0 4.2787e-08 0 4.279e-08 0.0007 4.2793e-08 0 4.2987e-08 0 4.299e-08 0.0007 4.2993e-08 0 4.3187e-08 0 4.319e-08 0.0007 4.3193e-08 0 4.3387e-08 0 4.339e-08 0.0007 4.3393e-08 0 4.3587e-08 0 4.359e-08 0.0007 4.3593e-08 0 4.3787e-08 0 4.379e-08 0.0007 4.3793e-08 0 4.3987e-08 0 4.399e-08 0.0007 4.3993e-08 0 4.4187e-08 0 4.419e-08 0.0007 4.4193e-08 0 4.4387e-08 0 4.439e-08 0.0007 4.4393e-08 0 4.4587e-08 0 4.459e-08 0.0007 4.4593e-08 0 4.4787e-08 0 4.479e-08 0.0007 4.4793e-08 0 4.4987e-08 0 4.499e-08 0.0007 4.4993e-08 0 4.5187e-08 0 4.519e-08 0.0007 4.5193e-08 0 4.5387e-08 0 4.539e-08 0.0007 4.5393e-08 0 4.5587e-08 0 4.559e-08 0.0007 4.5593e-08 0 4.5787e-08 0 4.579e-08 0.0007 4.5793e-08 0 4.5987e-08 0 4.599e-08 0.0007 4.5993e-08 0 4.6187e-08 0 4.619e-08 0.0007 4.6193e-08 0 4.6387e-08 0 4.639e-08 0.0007 4.6393e-08 0 4.6587e-08 0 4.659e-08 0.0007 4.6593e-08 0 4.6787e-08 0 4.679e-08 0.0007 4.6793e-08 0 4.6987e-08 0 4.699e-08 0.0007 4.6993e-08 0 4.7187e-08 0 4.719e-08 0.0007 4.7193e-08 0 4.7387e-08 0 4.739e-08 0.0007 4.7393e-08 0 4.7587e-08 0 4.759e-08 0.0007 4.7593e-08 0 4.7787e-08 0 4.779e-08 0.0007 4.7793e-08 0 4.7987e-08 0 4.799e-08 0.0007 4.7993e-08 0 4.8187e-08 0 4.819e-08 0.0007 4.8193e-08 0 4.8387e-08 0 4.839e-08 0.0007 4.8393e-08 0 4.8587e-08 0 4.859e-08 0.0007 4.8593e-08 0 4.8787e-08 0 4.879e-08 0.0007 4.8793e-08 0 4.8987e-08 0 4.899e-08 0.0007 4.8993e-08 0 4.9187e-08 0 4.919e-08 0.0007 4.9193e-08 0 4.9387e-08 0 4.939e-08 0.0007 4.9393e-08 0 4.9587e-08 0 4.959e-08 0.0007 4.9593e-08 0 4.9787e-08 0 4.979e-08 0.0007 4.9793e-08 0 4.9987e-08 0 4.999e-08 0.0007 4.9993e-08 0 5.0187e-08 0 5.019e-08 0.0007 5.0193e-08 0 5.0387e-08 0 5.039e-08 0.0007 5.0393e-08 0 5.0587e-08 0 5.059e-08 0.0007 5.0593e-08 0 5.0787e-08 0 5.079e-08 0.0007 5.0793e-08 0 5.0987e-08 0 5.099e-08 0.0007 5.0993e-08 0 5.1187e-08 0 5.119e-08 0.0007 5.1193e-08 0 5.1387e-08 0 5.139e-08 0.0007 5.1393e-08 0 5.1587e-08 0 5.159e-08 0.0007 5.1593e-08 0 5.1787e-08 0 5.179e-08 0.0007 5.1793e-08 0 5.1987e-08 0 5.199e-08 0.0007 5.1993e-08 0 5.2187e-08 0 5.219e-08 0.0007 5.2193e-08 0 5.2387e-08 0 5.239e-08 0.0007 5.2393e-08 0 5.2587e-08 0 5.259e-08 0.0007 5.2593e-08 0 5.2787e-08 0 5.279e-08 0.0007 5.2793e-08 0 5.2987e-08 0 5.299e-08 0.0007 5.2993e-08 0 5.3187e-08 0 5.319e-08 0.0007 5.3193e-08 0 5.3387e-08 0 5.339e-08 0.0007 5.3393e-08 0 5.3587e-08 0 5.359e-08 0.0007 5.3593e-08 0 5.3787e-08 0 5.379e-08 0.0007 5.3793e-08 0 5.3987e-08 0 5.399e-08 0.0007 5.3993e-08 0 5.4187e-08 0 5.419e-08 0.0007 5.4193e-08 0 5.4387e-08 0 5.439e-08 0.0007 5.4393e-08 0 5.4587e-08 0 5.459e-08 0.0007 5.4593e-08 0 5.4787e-08 0 5.479e-08 0.0007 5.4793e-08 0 5.4987e-08 0 5.499e-08 0.0007 5.4993e-08 0 5.5187e-08 0 5.519e-08 0.0007 5.5193e-08 0 5.5387e-08 0 5.539e-08 0.0007 5.5393e-08 0 5.5587e-08 0 5.559e-08 0.0007 5.5593e-08 0 5.5787e-08 0 5.579e-08 0.0007 5.5793e-08 0 5.5987e-08 0 5.599e-08 0.0007 5.5993e-08 0 5.6187e-08 0 5.619e-08 0.0007 5.6193e-08 0 5.6387e-08 0 5.639e-08 0.0007 5.6393e-08 0 5.6587e-08 0 5.659e-08 0.0007 5.6593e-08 0 5.6787e-08 0 5.679e-08 0.0007 5.6793e-08 0 5.6987e-08 0 5.699e-08 0.0007 5.6993e-08 0 5.7187e-08 0 5.719e-08 0.0007 5.7193e-08 0 5.7387e-08 0 5.739e-08 0.0007 5.7393e-08 0 5.7587e-08 0 5.759e-08 0.0007 5.7593e-08 0 5.7787e-08 0 5.779e-08 0.0007 5.7793e-08 0 5.7987e-08 0 5.799e-08 0.0007 5.7993e-08 0 5.8187e-08 0 5.819e-08 0.0007 5.8193e-08 0 5.8387e-08 0 5.839e-08 0.0007 5.8393e-08 0 5.8587e-08 0 5.859e-08 0.0007 5.8593e-08 0 5.8787e-08 0 5.879e-08 0.0007 5.8793e-08 0 5.8987e-08 0 5.899e-08 0.0007 5.8993e-08 0 5.9187e-08 0 5.919e-08 0.0007 5.9193e-08 0 5.9387e-08 0 5.939e-08 0.0007 5.9393e-08 0 5.9587e-08 0 5.959e-08 0.0007 5.9593e-08 0 5.9787e-08 0 5.979e-08 0.0007 5.9793e-08 0 5.9987e-08 0 5.999e-08 0.0007 5.9993e-08 0 6.0187e-08 0 6.019e-08 0.0007 6.0193e-08 0 6.0387e-08 0 6.039e-08 0.0007 6.0393e-08 0 6.0587e-08 0 6.059e-08 0.0007 6.0593e-08 0 6.0787e-08 0 6.079e-08 0.0007 6.0793e-08 0 6.0987e-08 0 6.099e-08 0.0007 6.0993e-08 0 6.1187e-08 0 6.119e-08 0.0007 6.1193e-08 0 6.1387e-08 0 6.139e-08 0.0007 6.1393e-08 0 6.1587e-08 0 6.159e-08 0.0007 6.1593e-08 0 6.1787e-08 0 6.179e-08 0.0007 6.1793e-08 0 6.1987e-08 0 6.199e-08 0.0007 6.1993e-08 0 6.2187e-08 0 6.219e-08 0.0007 6.2193e-08 0 6.2387e-08 0 6.239e-08 0.0007 6.2393e-08 0 6.2587e-08 0 6.259e-08 0.0007 6.2593e-08 0 6.2787e-08 0 6.279e-08 0.0007 6.2793e-08 0 6.2987e-08 0 6.299e-08 0.0007 6.2993e-08 0 6.3187e-08 0 6.319e-08 0.0007 6.3193e-08 0 6.3387e-08 0 6.339e-08 0.0007 6.3393e-08 0 6.3587e-08 0 6.359e-08 0.0007 6.3593e-08 0 6.3787e-08 0 6.379e-08 0.0007 6.3793e-08 0 6.3987e-08 0 6.399e-08 0.0007 6.3993e-08 0 6.4187e-08 0 6.419e-08 0.0007 6.4193e-08 0 6.4387e-08 0 6.439e-08 0.0007 6.4393e-08 0 6.4587e-08 0 6.459e-08 0.0007 6.4593e-08 0 6.4787e-08 0 6.479e-08 0.0007 6.4793e-08 0 6.4987e-08 0 6.499e-08 0.0007 6.4993e-08 0 6.5187e-08 0 6.519e-08 0.0007 6.5193e-08 0 6.5387e-08 0 6.539e-08 0.0007 6.5393e-08 0 6.5587e-08 0 6.559e-08 0.0007 6.5593e-08 0 6.5787e-08 0 6.579e-08 0.0007 6.5793e-08 0 6.5987e-08 0 6.599e-08 0.0007 6.5993e-08 0 6.6187e-08 0 6.619e-08 0.0007 6.6193e-08 0 6.6387e-08 0 6.639e-08 0.0007 6.6393e-08 0 6.6587e-08 0 6.659e-08 0.0007 6.6593e-08 0 6.6787e-08 0 6.679e-08 0.0007 6.6793e-08 0 6.6987e-08 0 6.699e-08 0.0007 6.6993e-08 0 6.7187e-08 0 6.719e-08 0.0007 6.7193e-08 0 6.7387e-08 0 6.739e-08 0.0007 6.7393e-08 0 6.7587e-08 0 6.759e-08 0.0007 6.7593e-08 0 6.7787e-08 0 6.779e-08 0.0007 6.7793e-08 0 6.7987e-08 0 6.799e-08 0.0007 6.7993e-08 0 6.8187e-08 0 6.819e-08 0.0007 6.8193e-08 0 6.8387e-08 0 6.839e-08 0.0007 6.8393e-08 0 6.8587e-08 0 6.859e-08 0.0007 6.8593e-08 0 6.8787e-08 0 6.879e-08 0.0007 6.8793e-08 0 6.8987e-08 0 6.899e-08 0.0007 6.8993e-08 0 6.9187e-08 0 6.919e-08 0.0007 6.9193e-08 0 6.9387e-08 0 6.939e-08 0.0007 6.9393e-08 0 6.9587e-08 0 6.959e-08 0.0007 6.9593e-08 0 6.9787e-08 0 6.979e-08 0.0007 6.9793e-08 0 6.9987e-08 0 6.999e-08 0.0007 6.9993e-08 0 7.0187e-08 0 7.019e-08 0.0007 7.0193e-08 0 7.0387e-08 0 7.039e-08 0.0007 7.0393e-08 0 7.0587e-08 0 7.059e-08 0.0007 7.0593e-08 0 7.0787e-08 0 7.079e-08 0.0007 7.0793e-08 0 7.0987e-08 0 7.099e-08 0.0007 7.0993e-08 0 7.1187e-08 0 7.119e-08 0.0007 7.1193e-08 0 7.1387e-08 0 7.139e-08 0.0007 7.1393e-08 0 7.1587e-08 0 7.159e-08 0.0007 7.1593e-08 0 7.1787e-08 0 7.179e-08 0.0007 7.1793e-08 0 7.1987e-08 0 7.199e-08 0.0007 7.1993e-08 0 7.2187e-08 0 7.219e-08 0.0007 7.2193e-08 0 7.2387e-08 0 7.239e-08 0.0007 7.2393e-08 0 7.2587e-08 0 7.259e-08 0.0007 7.2593e-08 0 7.2787e-08 0 7.279e-08 0.0007 7.2793e-08 0 7.2987e-08 0 7.299e-08 0.0007 7.2993e-08 0 7.3187e-08 0 7.319e-08 0.0007 7.3193e-08 0 7.3387e-08 0 7.339e-08 0.0007 7.3393e-08 0 7.3587e-08 0 7.359e-08 0.0007 7.3593e-08 0 7.3787e-08 0 7.379e-08 0.0007 7.3793e-08 0 7.3987e-08 0 7.399e-08 0.0007 7.3993e-08 0 7.4187e-08 0 7.419e-08 0.0007 7.4193e-08 0 7.4387e-08 0 7.439e-08 0.0007 7.4393e-08 0 7.4587e-08 0 7.459e-08 0.0007 7.4593e-08 0 7.4787e-08 0 7.479e-08 0.0007 7.4793e-08 0 7.4987e-08 0 7.499e-08 0.0007 7.4993e-08 0 7.5187e-08 0 7.519e-08 0.0007 7.5193e-08 0 7.5387e-08 0 7.539e-08 0.0007 7.5393e-08 0 7.5587e-08 0 7.559e-08 0.0007 7.5593e-08 0 7.5787e-08 0 7.579e-08 0.0007 7.5793e-08 0 7.5987e-08 0 7.599e-08 0.0007 7.5993e-08 0 7.6187e-08 0 7.619e-08 0.0007 7.6193e-08 0 7.6387e-08 0 7.639e-08 0.0007 7.6393e-08 0 7.6587e-08 0 7.659e-08 0.0007 7.6593e-08 0 7.6787e-08 0 7.679e-08 0.0007 7.6793e-08 0 7.6987e-08 0 7.699e-08 0.0007 7.6993e-08 0 7.7187e-08 0 7.719e-08 0.0007 7.7193e-08 0 7.7387e-08 0 7.739e-08 0.0007 7.7393e-08 0 7.7587e-08 0 7.759e-08 0.0007 7.7593e-08 0 7.7787e-08 0 7.779e-08 0.0007 7.7793e-08 0 7.7987e-08 0 7.799e-08 0.0007 7.7993e-08 0 7.8187e-08 0 7.819e-08 0.0007 7.8193e-08 0 7.8387e-08 0 7.839e-08 0.0007 7.8393e-08 0 7.8587e-08 0 7.859e-08 0.0007 7.8593e-08 0 7.8787e-08 0 7.879e-08 0.0007 7.8793e-08 0 7.8987e-08 0 7.899e-08 0.0007 7.8993e-08 0 7.9187e-08 0 7.919e-08 0.0007 7.9193e-08 0 7.9387e-08 0 7.939e-08 0.0007 7.9393e-08 0 7.9587e-08 0 7.959e-08 0.0007 7.9593e-08 0)
L_S8_45|1 S8_4 _S8_45|A1  2.067833848e-12
L_S8_45|2 _S8_45|A1 _S8_45|A2  4.135667696e-12
L_S8_45|3 _S8_45|A3 _S8_45|A4  8.271335392e-12
L_S8_45|T T58 _S8_45|T1  2.067833848e-12
L_S8_45|4 _S8_45|T1 _S8_45|T2  4.135667696e-12
L_S8_45|5 _S8_45|A4 _S8_45|Q1  4.135667696e-12
L_S8_45|6 _S8_45|Q1 S8_5_TX  2.067833848e-12
B_PTL_A0|_TX|1 _PTL_A0|_TX|1 _PTL_A0|_TX|2 JJMIT AREA=2.5
B_PTL_A0|_TX|2 _PTL_A0|_TX|4 _PTL_A0|_TX|5 JJMIT AREA=2.5
I_PTL_A0|_TX|B1 0 _PTL_A0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A0|_TX|B2 0 _PTL_A0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|3  1.684e-12
L_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|6  3.596e-12
L_PTL_A0|_TX|1 A0_TX _PTL_A0|_TX|1  2.063e-12
L_PTL_A0|_TX|2 _PTL_A0|_TX|1 _PTL_A0|_TX|4  4.123e-12
L_PTL_A0|_TX|3 _PTL_A0|_TX|4 _PTL_A0|_TX|7  2.193e-12
R_PTL_A0|_TX|D _PTL_A0|_TX|7 _PTL_A0|A_PTL  1.36
L_PTL_A0|_TX|P1 _PTL_A0|_TX|2 0  5.254e-13
L_PTL_A0|_TX|P2 _PTL_A0|_TX|5 0  5.141e-13
R_PTL_A0|_TX|B1 _PTL_A0|_TX|1 _PTL_A0|_TX|101  2.7439617672
R_PTL_A0|_TX|B2 _PTL_A0|_TX|4 _PTL_A0|_TX|104  2.7439617672
L_PTL_A0|_TX|RB1 _PTL_A0|_TX|101 0  1.550338398468e-12
L_PTL_A0|_TX|RB2 _PTL_A0|_TX|104 0  1.550338398468e-12
B_PTL_A0|_RX|1 _PTL_A0|_RX|1 _PTL_A0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A0|_RX|2 _PTL_A0|_RX|4 _PTL_A0|_RX|5 JJMIT AREA=2.0
B_PTL_A0|_RX|3 _PTL_A0|_RX|7 _PTL_A0|_RX|8 JJMIT AREA=2.5
I_PTL_A0|_RX|B1 0 _PTL_A0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|3  2.777e-12
I_PTL_A0|_RX|B2 0 _PTL_A0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|6  2.685e-12
I_PTL_A0|_RX|B3 0 _PTL_A0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|9  2.764e-12
L_PTL_A0|_RX|1 _PTL_A0|A_PTL _PTL_A0|_RX|1  1.346e-12
L_PTL_A0|_RX|2 _PTL_A0|_RX|1 _PTL_A0|_RX|4  6.348e-12
L_PTL_A0|_RX|3 _PTL_A0|_RX|4 _PTL_A0|_RX|7  5.197e-12
L_PTL_A0|_RX|4 _PTL_A0|_RX|7 _PTL_A0|A_PTL_RX  2.058e-12
L_PTL_A0|_RX|P1 _PTL_A0|_RX|2 0  4.795e-13
L_PTL_A0|_RX|P2 _PTL_A0|_RX|5 0  5.431e-13
L_PTL_A0|_RX|P3 _PTL_A0|_RX|8 0  5.339e-13
R_PTL_A0|_RX|B1 _PTL_A0|_RX|1 _PTL_A0|_RX|101  4.225701121488
R_PTL_A0|_RX|B2 _PTL_A0|_RX|4 _PTL_A0|_RX|104  3.429952209
R_PTL_A0|_RX|B3 _PTL_A0|_RX|7 _PTL_A0|_RX|107  2.7439617672
L_PTL_A0|_RX|RB1 _PTL_A0|_RX|101 0  2.38752113364072e-12
L_PTL_A0|_RX|RB2 _PTL_A0|_RX|104 0  1.937922998085e-12
L_PTL_A0|_RX|RB3 _PTL_A0|_RX|107 0  1.550338398468e-12
B_PTL_A0|_JTL|1 _PTL_A0|_JTL|1 _PTL_A0|_JTL|2 JJMIT AREA=2.5
B_PTL_A0|_JTL|2 _PTL_A0|_JTL|6 _PTL_A0|_JTL|7 JJMIT AREA=2.5
I_PTL_A0|_JTL|B1 0 _PTL_A0|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A0|_JTL|1 _PTL_A0|A_PTL_RX _PTL_A0|_JTL|1  2.067833848e-12
L_PTL_A0|_JTL|2 _PTL_A0|_JTL|1 _PTL_A0|_JTL|4  2.067833848e-12
L_PTL_A0|_JTL|3 _PTL_A0|_JTL|4 _PTL_A0|_JTL|6  2.067833848e-12
L_PTL_A0|_JTL|4 _PTL_A0|_JTL|6 A0_RX  2.067833848e-12
L_PTL_A0|_JTL|P1 _PTL_A0|_JTL|2 0  2e-13
L_PTL_A0|_JTL|P2 _PTL_A0|_JTL|7 0  2e-13
L_PTL_A0|_JTL|B1 _PTL_A0|_JTL|5 _PTL_A0|_JTL|4  2e-12
R_PTL_A0|_JTL|B1 _PTL_A0|_JTL|1 _PTL_A0|_JTL|3  2.7439617672
R_PTL_A0|_JTL|B2 _PTL_A0|_JTL|6 _PTL_A0|_JTL|8  2.7439617672
L_PTL_A0|_JTL|RB1 _PTL_A0|_JTL|3 0  1.750338398468e-12
L_PTL_A0|_JTL|RB2 _PTL_A0|_JTL|8 0  1.750338398468e-12
B_PTL_B0|_TX|1 _PTL_B0|_TX|1 _PTL_B0|_TX|2 JJMIT AREA=2.5
B_PTL_B0|_TX|2 _PTL_B0|_TX|4 _PTL_B0|_TX|5 JJMIT AREA=2.5
I_PTL_B0|_TX|B1 0 _PTL_B0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B0|_TX|B2 0 _PTL_B0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|3  1.684e-12
L_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|6  3.596e-12
L_PTL_B0|_TX|1 B0_TX _PTL_B0|_TX|1  2.063e-12
L_PTL_B0|_TX|2 _PTL_B0|_TX|1 _PTL_B0|_TX|4  4.123e-12
L_PTL_B0|_TX|3 _PTL_B0|_TX|4 _PTL_B0|_TX|7  2.193e-12
R_PTL_B0|_TX|D _PTL_B0|_TX|7 _PTL_B0|A_PTL  1.36
L_PTL_B0|_TX|P1 _PTL_B0|_TX|2 0  5.254e-13
L_PTL_B0|_TX|P2 _PTL_B0|_TX|5 0  5.141e-13
R_PTL_B0|_TX|B1 _PTL_B0|_TX|1 _PTL_B0|_TX|101  2.7439617672
R_PTL_B0|_TX|B2 _PTL_B0|_TX|4 _PTL_B0|_TX|104  2.7439617672
L_PTL_B0|_TX|RB1 _PTL_B0|_TX|101 0  1.550338398468e-12
L_PTL_B0|_TX|RB2 _PTL_B0|_TX|104 0  1.550338398468e-12
B_PTL_B0|_RX|1 _PTL_B0|_RX|1 _PTL_B0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B0|_RX|2 _PTL_B0|_RX|4 _PTL_B0|_RX|5 JJMIT AREA=2.0
B_PTL_B0|_RX|3 _PTL_B0|_RX|7 _PTL_B0|_RX|8 JJMIT AREA=2.5
I_PTL_B0|_RX|B1 0 _PTL_B0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|3  2.777e-12
I_PTL_B0|_RX|B2 0 _PTL_B0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|6  2.685e-12
I_PTL_B0|_RX|B3 0 _PTL_B0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|9  2.764e-12
L_PTL_B0|_RX|1 _PTL_B0|A_PTL _PTL_B0|_RX|1  1.346e-12
L_PTL_B0|_RX|2 _PTL_B0|_RX|1 _PTL_B0|_RX|4  6.348e-12
L_PTL_B0|_RX|3 _PTL_B0|_RX|4 _PTL_B0|_RX|7  5.197e-12
L_PTL_B0|_RX|4 _PTL_B0|_RX|7 _PTL_B0|A_PTL_RX  2.058e-12
L_PTL_B0|_RX|P1 _PTL_B0|_RX|2 0  4.795e-13
L_PTL_B0|_RX|P2 _PTL_B0|_RX|5 0  5.431e-13
L_PTL_B0|_RX|P3 _PTL_B0|_RX|8 0  5.339e-13
R_PTL_B0|_RX|B1 _PTL_B0|_RX|1 _PTL_B0|_RX|101  4.225701121488
R_PTL_B0|_RX|B2 _PTL_B0|_RX|4 _PTL_B0|_RX|104  3.429952209
R_PTL_B0|_RX|B3 _PTL_B0|_RX|7 _PTL_B0|_RX|107  2.7439617672
L_PTL_B0|_RX|RB1 _PTL_B0|_RX|101 0  2.38752113364072e-12
L_PTL_B0|_RX|RB2 _PTL_B0|_RX|104 0  1.937922998085e-12
L_PTL_B0|_RX|RB3 _PTL_B0|_RX|107 0  1.550338398468e-12
B_PTL_B0|_JTL|1 _PTL_B0|_JTL|1 _PTL_B0|_JTL|2 JJMIT AREA=2.5
B_PTL_B0|_JTL|2 _PTL_B0|_JTL|6 _PTL_B0|_JTL|7 JJMIT AREA=2.5
I_PTL_B0|_JTL|B1 0 _PTL_B0|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B0|_JTL|1 _PTL_B0|A_PTL_RX _PTL_B0|_JTL|1  2.067833848e-12
L_PTL_B0|_JTL|2 _PTL_B0|_JTL|1 _PTL_B0|_JTL|4  2.067833848e-12
L_PTL_B0|_JTL|3 _PTL_B0|_JTL|4 _PTL_B0|_JTL|6  2.067833848e-12
L_PTL_B0|_JTL|4 _PTL_B0|_JTL|6 B0_RX  2.067833848e-12
L_PTL_B0|_JTL|P1 _PTL_B0|_JTL|2 0  2e-13
L_PTL_B0|_JTL|P2 _PTL_B0|_JTL|7 0  2e-13
L_PTL_B0|_JTL|B1 _PTL_B0|_JTL|5 _PTL_B0|_JTL|4  2e-12
R_PTL_B0|_JTL|B1 _PTL_B0|_JTL|1 _PTL_B0|_JTL|3  2.7439617672
R_PTL_B0|_JTL|B2 _PTL_B0|_JTL|6 _PTL_B0|_JTL|8  2.7439617672
L_PTL_B0|_JTL|RB1 _PTL_B0|_JTL|3 0  1.750338398468e-12
L_PTL_B0|_JTL|RB2 _PTL_B0|_JTL|8 0  1.750338398468e-12
B_PTL_A1|_TX|1 _PTL_A1|_TX|1 _PTL_A1|_TX|2 JJMIT AREA=2.5
B_PTL_A1|_TX|2 _PTL_A1|_TX|4 _PTL_A1|_TX|5 JJMIT AREA=2.5
I_PTL_A1|_TX|B1 0 _PTL_A1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A1|_TX|B2 0 _PTL_A1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|3  1.684e-12
L_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|6  3.596e-12
L_PTL_A1|_TX|1 A1_TX _PTL_A1|_TX|1  2.063e-12
L_PTL_A1|_TX|2 _PTL_A1|_TX|1 _PTL_A1|_TX|4  4.123e-12
L_PTL_A1|_TX|3 _PTL_A1|_TX|4 _PTL_A1|_TX|7  2.193e-12
R_PTL_A1|_TX|D _PTL_A1|_TX|7 _PTL_A1|A_PTL  1.36
L_PTL_A1|_TX|P1 _PTL_A1|_TX|2 0  5.254e-13
L_PTL_A1|_TX|P2 _PTL_A1|_TX|5 0  5.141e-13
R_PTL_A1|_TX|B1 _PTL_A1|_TX|1 _PTL_A1|_TX|101  2.7439617672
R_PTL_A1|_TX|B2 _PTL_A1|_TX|4 _PTL_A1|_TX|104  2.7439617672
L_PTL_A1|_TX|RB1 _PTL_A1|_TX|101 0  1.550338398468e-12
L_PTL_A1|_TX|RB2 _PTL_A1|_TX|104 0  1.550338398468e-12
B_PTL_A1|_RX|1 _PTL_A1|_RX|1 _PTL_A1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A1|_RX|2 _PTL_A1|_RX|4 _PTL_A1|_RX|5 JJMIT AREA=2.0
B_PTL_A1|_RX|3 _PTL_A1|_RX|7 _PTL_A1|_RX|8 JJMIT AREA=2.5
I_PTL_A1|_RX|B1 0 _PTL_A1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|3  2.777e-12
I_PTL_A1|_RX|B2 0 _PTL_A1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|6  2.685e-12
I_PTL_A1|_RX|B3 0 _PTL_A1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|9  2.764e-12
L_PTL_A1|_RX|1 _PTL_A1|A_PTL _PTL_A1|_RX|1  1.346e-12
L_PTL_A1|_RX|2 _PTL_A1|_RX|1 _PTL_A1|_RX|4  6.348e-12
L_PTL_A1|_RX|3 _PTL_A1|_RX|4 _PTL_A1|_RX|7  5.197e-12
L_PTL_A1|_RX|4 _PTL_A1|_RX|7 _PTL_A1|A_PTL_RX  2.058e-12
L_PTL_A1|_RX|P1 _PTL_A1|_RX|2 0  4.795e-13
L_PTL_A1|_RX|P2 _PTL_A1|_RX|5 0  5.431e-13
L_PTL_A1|_RX|P3 _PTL_A1|_RX|8 0  5.339e-13
R_PTL_A1|_RX|B1 _PTL_A1|_RX|1 _PTL_A1|_RX|101  4.225701121488
R_PTL_A1|_RX|B2 _PTL_A1|_RX|4 _PTL_A1|_RX|104  3.429952209
R_PTL_A1|_RX|B3 _PTL_A1|_RX|7 _PTL_A1|_RX|107  2.7439617672
L_PTL_A1|_RX|RB1 _PTL_A1|_RX|101 0  2.38752113364072e-12
L_PTL_A1|_RX|RB2 _PTL_A1|_RX|104 0  1.937922998085e-12
L_PTL_A1|_RX|RB3 _PTL_A1|_RX|107 0  1.550338398468e-12
B_PTL_A1|_JTL|1 _PTL_A1|_JTL|1 _PTL_A1|_JTL|2 JJMIT AREA=2.5
B_PTL_A1|_JTL|2 _PTL_A1|_JTL|6 _PTL_A1|_JTL|7 JJMIT AREA=2.5
I_PTL_A1|_JTL|B1 0 _PTL_A1|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A1|_JTL|1 _PTL_A1|A_PTL_RX _PTL_A1|_JTL|1  2.067833848e-12
L_PTL_A1|_JTL|2 _PTL_A1|_JTL|1 _PTL_A1|_JTL|4  2.067833848e-12
L_PTL_A1|_JTL|3 _PTL_A1|_JTL|4 _PTL_A1|_JTL|6  2.067833848e-12
L_PTL_A1|_JTL|4 _PTL_A1|_JTL|6 A1_RX  2.067833848e-12
L_PTL_A1|_JTL|P1 _PTL_A1|_JTL|2 0  2e-13
L_PTL_A1|_JTL|P2 _PTL_A1|_JTL|7 0  2e-13
L_PTL_A1|_JTL|B1 _PTL_A1|_JTL|5 _PTL_A1|_JTL|4  2e-12
R_PTL_A1|_JTL|B1 _PTL_A1|_JTL|1 _PTL_A1|_JTL|3  2.7439617672
R_PTL_A1|_JTL|B2 _PTL_A1|_JTL|6 _PTL_A1|_JTL|8  2.7439617672
L_PTL_A1|_JTL|RB1 _PTL_A1|_JTL|3 0  1.750338398468e-12
L_PTL_A1|_JTL|RB2 _PTL_A1|_JTL|8 0  1.750338398468e-12
B_PTL_B1|_TX|1 _PTL_B1|_TX|1 _PTL_B1|_TX|2 JJMIT AREA=2.5
B_PTL_B1|_TX|2 _PTL_B1|_TX|4 _PTL_B1|_TX|5 JJMIT AREA=2.5
I_PTL_B1|_TX|B1 0 _PTL_B1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B1|_TX|B2 0 _PTL_B1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|3  1.684e-12
L_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|6  3.596e-12
L_PTL_B1|_TX|1 B1_TX _PTL_B1|_TX|1  2.063e-12
L_PTL_B1|_TX|2 _PTL_B1|_TX|1 _PTL_B1|_TX|4  4.123e-12
L_PTL_B1|_TX|3 _PTL_B1|_TX|4 _PTL_B1|_TX|7  2.193e-12
R_PTL_B1|_TX|D _PTL_B1|_TX|7 _PTL_B1|A_PTL  1.36
L_PTL_B1|_TX|P1 _PTL_B1|_TX|2 0  5.254e-13
L_PTL_B1|_TX|P2 _PTL_B1|_TX|5 0  5.141e-13
R_PTL_B1|_TX|B1 _PTL_B1|_TX|1 _PTL_B1|_TX|101  2.7439617672
R_PTL_B1|_TX|B2 _PTL_B1|_TX|4 _PTL_B1|_TX|104  2.7439617672
L_PTL_B1|_TX|RB1 _PTL_B1|_TX|101 0  1.550338398468e-12
L_PTL_B1|_TX|RB2 _PTL_B1|_TX|104 0  1.550338398468e-12
B_PTL_B1|_RX|1 _PTL_B1|_RX|1 _PTL_B1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B1|_RX|2 _PTL_B1|_RX|4 _PTL_B1|_RX|5 JJMIT AREA=2.0
B_PTL_B1|_RX|3 _PTL_B1|_RX|7 _PTL_B1|_RX|8 JJMIT AREA=2.5
I_PTL_B1|_RX|B1 0 _PTL_B1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|3  2.777e-12
I_PTL_B1|_RX|B2 0 _PTL_B1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|6  2.685e-12
I_PTL_B1|_RX|B3 0 _PTL_B1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|9  2.764e-12
L_PTL_B1|_RX|1 _PTL_B1|A_PTL _PTL_B1|_RX|1  1.346e-12
L_PTL_B1|_RX|2 _PTL_B1|_RX|1 _PTL_B1|_RX|4  6.348e-12
L_PTL_B1|_RX|3 _PTL_B1|_RX|4 _PTL_B1|_RX|7  5.197e-12
L_PTL_B1|_RX|4 _PTL_B1|_RX|7 _PTL_B1|A_PTL_RX  2.058e-12
L_PTL_B1|_RX|P1 _PTL_B1|_RX|2 0  4.795e-13
L_PTL_B1|_RX|P2 _PTL_B1|_RX|5 0  5.431e-13
L_PTL_B1|_RX|P3 _PTL_B1|_RX|8 0  5.339e-13
R_PTL_B1|_RX|B1 _PTL_B1|_RX|1 _PTL_B1|_RX|101  4.225701121488
R_PTL_B1|_RX|B2 _PTL_B1|_RX|4 _PTL_B1|_RX|104  3.429952209
R_PTL_B1|_RX|B3 _PTL_B1|_RX|7 _PTL_B1|_RX|107  2.7439617672
L_PTL_B1|_RX|RB1 _PTL_B1|_RX|101 0  2.38752113364072e-12
L_PTL_B1|_RX|RB2 _PTL_B1|_RX|104 0  1.937922998085e-12
L_PTL_B1|_RX|RB3 _PTL_B1|_RX|107 0  1.550338398468e-12
B_PTL_B1|_JTL|1 _PTL_B1|_JTL|1 _PTL_B1|_JTL|2 JJMIT AREA=2.5
B_PTL_B1|_JTL|2 _PTL_B1|_JTL|6 _PTL_B1|_JTL|7 JJMIT AREA=2.5
I_PTL_B1|_JTL|B1 0 _PTL_B1|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B1|_JTL|1 _PTL_B1|A_PTL_RX _PTL_B1|_JTL|1  2.067833848e-12
L_PTL_B1|_JTL|2 _PTL_B1|_JTL|1 _PTL_B1|_JTL|4  2.067833848e-12
L_PTL_B1|_JTL|3 _PTL_B1|_JTL|4 _PTL_B1|_JTL|6  2.067833848e-12
L_PTL_B1|_JTL|4 _PTL_B1|_JTL|6 B1_RX  2.067833848e-12
L_PTL_B1|_JTL|P1 _PTL_B1|_JTL|2 0  2e-13
L_PTL_B1|_JTL|P2 _PTL_B1|_JTL|7 0  2e-13
L_PTL_B1|_JTL|B1 _PTL_B1|_JTL|5 _PTL_B1|_JTL|4  2e-12
R_PTL_B1|_JTL|B1 _PTL_B1|_JTL|1 _PTL_B1|_JTL|3  2.7439617672
R_PTL_B1|_JTL|B2 _PTL_B1|_JTL|6 _PTL_B1|_JTL|8  2.7439617672
L_PTL_B1|_JTL|RB1 _PTL_B1|_JTL|3 0  1.750338398468e-12
L_PTL_B1|_JTL|RB2 _PTL_B1|_JTL|8 0  1.750338398468e-12
B_PTL_A2|_TX|1 _PTL_A2|_TX|1 _PTL_A2|_TX|2 JJMIT AREA=2.5
B_PTL_A2|_TX|2 _PTL_A2|_TX|4 _PTL_A2|_TX|5 JJMIT AREA=2.5
I_PTL_A2|_TX|B1 0 _PTL_A2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A2|_TX|B2 0 _PTL_A2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|3  1.684e-12
L_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|6  3.596e-12
L_PTL_A2|_TX|1 A2_TX _PTL_A2|_TX|1  2.063e-12
L_PTL_A2|_TX|2 _PTL_A2|_TX|1 _PTL_A2|_TX|4  4.123e-12
L_PTL_A2|_TX|3 _PTL_A2|_TX|4 _PTL_A2|_TX|7  2.193e-12
R_PTL_A2|_TX|D _PTL_A2|_TX|7 _PTL_A2|A_PTL  1.36
L_PTL_A2|_TX|P1 _PTL_A2|_TX|2 0  5.254e-13
L_PTL_A2|_TX|P2 _PTL_A2|_TX|5 0  5.141e-13
R_PTL_A2|_TX|B1 _PTL_A2|_TX|1 _PTL_A2|_TX|101  2.7439617672
R_PTL_A2|_TX|B2 _PTL_A2|_TX|4 _PTL_A2|_TX|104  2.7439617672
L_PTL_A2|_TX|RB1 _PTL_A2|_TX|101 0  1.550338398468e-12
L_PTL_A2|_TX|RB2 _PTL_A2|_TX|104 0  1.550338398468e-12
B_PTL_A2|_RX|1 _PTL_A2|_RX|1 _PTL_A2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A2|_RX|2 _PTL_A2|_RX|4 _PTL_A2|_RX|5 JJMIT AREA=2.0
B_PTL_A2|_RX|3 _PTL_A2|_RX|7 _PTL_A2|_RX|8 JJMIT AREA=2.5
I_PTL_A2|_RX|B1 0 _PTL_A2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|3  2.777e-12
I_PTL_A2|_RX|B2 0 _PTL_A2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|6  2.685e-12
I_PTL_A2|_RX|B3 0 _PTL_A2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|9  2.764e-12
L_PTL_A2|_RX|1 _PTL_A2|A_PTL _PTL_A2|_RX|1  1.346e-12
L_PTL_A2|_RX|2 _PTL_A2|_RX|1 _PTL_A2|_RX|4  6.348e-12
L_PTL_A2|_RX|3 _PTL_A2|_RX|4 _PTL_A2|_RX|7  5.197e-12
L_PTL_A2|_RX|4 _PTL_A2|_RX|7 _PTL_A2|A_PTL_RX  2.058e-12
L_PTL_A2|_RX|P1 _PTL_A2|_RX|2 0  4.795e-13
L_PTL_A2|_RX|P2 _PTL_A2|_RX|5 0  5.431e-13
L_PTL_A2|_RX|P3 _PTL_A2|_RX|8 0  5.339e-13
R_PTL_A2|_RX|B1 _PTL_A2|_RX|1 _PTL_A2|_RX|101  4.225701121488
R_PTL_A2|_RX|B2 _PTL_A2|_RX|4 _PTL_A2|_RX|104  3.429952209
R_PTL_A2|_RX|B3 _PTL_A2|_RX|7 _PTL_A2|_RX|107  2.7439617672
L_PTL_A2|_RX|RB1 _PTL_A2|_RX|101 0  2.38752113364072e-12
L_PTL_A2|_RX|RB2 _PTL_A2|_RX|104 0  1.937922998085e-12
L_PTL_A2|_RX|RB3 _PTL_A2|_RX|107 0  1.550338398468e-12
B_PTL_A2|_JTL|1 _PTL_A2|_JTL|1 _PTL_A2|_JTL|2 JJMIT AREA=2.5
B_PTL_A2|_JTL|2 _PTL_A2|_JTL|6 _PTL_A2|_JTL|7 JJMIT AREA=2.5
I_PTL_A2|_JTL|B1 0 _PTL_A2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A2|_JTL|1 _PTL_A2|A_PTL_RX _PTL_A2|_JTL|1  2.067833848e-12
L_PTL_A2|_JTL|2 _PTL_A2|_JTL|1 _PTL_A2|_JTL|4  2.067833848e-12
L_PTL_A2|_JTL|3 _PTL_A2|_JTL|4 _PTL_A2|_JTL|6  2.067833848e-12
L_PTL_A2|_JTL|4 _PTL_A2|_JTL|6 A2_RX  2.067833848e-12
L_PTL_A2|_JTL|P1 _PTL_A2|_JTL|2 0  2e-13
L_PTL_A2|_JTL|P2 _PTL_A2|_JTL|7 0  2e-13
L_PTL_A2|_JTL|B1 _PTL_A2|_JTL|5 _PTL_A2|_JTL|4  2e-12
R_PTL_A2|_JTL|B1 _PTL_A2|_JTL|1 _PTL_A2|_JTL|3  2.7439617672
R_PTL_A2|_JTL|B2 _PTL_A2|_JTL|6 _PTL_A2|_JTL|8  2.7439617672
L_PTL_A2|_JTL|RB1 _PTL_A2|_JTL|3 0  1.750338398468e-12
L_PTL_A2|_JTL|RB2 _PTL_A2|_JTL|8 0  1.750338398468e-12
B_PTL_B2|_TX|1 _PTL_B2|_TX|1 _PTL_B2|_TX|2 JJMIT AREA=2.5
B_PTL_B2|_TX|2 _PTL_B2|_TX|4 _PTL_B2|_TX|5 JJMIT AREA=2.5
I_PTL_B2|_TX|B1 0 _PTL_B2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B2|_TX|B2 0 _PTL_B2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|3  1.684e-12
L_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|6  3.596e-12
L_PTL_B2|_TX|1 B2_TX _PTL_B2|_TX|1  2.063e-12
L_PTL_B2|_TX|2 _PTL_B2|_TX|1 _PTL_B2|_TX|4  4.123e-12
L_PTL_B2|_TX|3 _PTL_B2|_TX|4 _PTL_B2|_TX|7  2.193e-12
R_PTL_B2|_TX|D _PTL_B2|_TX|7 _PTL_B2|A_PTL  1.36
L_PTL_B2|_TX|P1 _PTL_B2|_TX|2 0  5.254e-13
L_PTL_B2|_TX|P2 _PTL_B2|_TX|5 0  5.141e-13
R_PTL_B2|_TX|B1 _PTL_B2|_TX|1 _PTL_B2|_TX|101  2.7439617672
R_PTL_B2|_TX|B2 _PTL_B2|_TX|4 _PTL_B2|_TX|104  2.7439617672
L_PTL_B2|_TX|RB1 _PTL_B2|_TX|101 0  1.550338398468e-12
L_PTL_B2|_TX|RB2 _PTL_B2|_TX|104 0  1.550338398468e-12
B_PTL_B2|_RX|1 _PTL_B2|_RX|1 _PTL_B2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B2|_RX|2 _PTL_B2|_RX|4 _PTL_B2|_RX|5 JJMIT AREA=2.0
B_PTL_B2|_RX|3 _PTL_B2|_RX|7 _PTL_B2|_RX|8 JJMIT AREA=2.5
I_PTL_B2|_RX|B1 0 _PTL_B2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|3  2.777e-12
I_PTL_B2|_RX|B2 0 _PTL_B2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|6  2.685e-12
I_PTL_B2|_RX|B3 0 _PTL_B2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|9  2.764e-12
L_PTL_B2|_RX|1 _PTL_B2|A_PTL _PTL_B2|_RX|1  1.346e-12
L_PTL_B2|_RX|2 _PTL_B2|_RX|1 _PTL_B2|_RX|4  6.348e-12
L_PTL_B2|_RX|3 _PTL_B2|_RX|4 _PTL_B2|_RX|7  5.197e-12
L_PTL_B2|_RX|4 _PTL_B2|_RX|7 _PTL_B2|A_PTL_RX  2.058e-12
L_PTL_B2|_RX|P1 _PTL_B2|_RX|2 0  4.795e-13
L_PTL_B2|_RX|P2 _PTL_B2|_RX|5 0  5.431e-13
L_PTL_B2|_RX|P3 _PTL_B2|_RX|8 0  5.339e-13
R_PTL_B2|_RX|B1 _PTL_B2|_RX|1 _PTL_B2|_RX|101  4.225701121488
R_PTL_B2|_RX|B2 _PTL_B2|_RX|4 _PTL_B2|_RX|104  3.429952209
R_PTL_B2|_RX|B3 _PTL_B2|_RX|7 _PTL_B2|_RX|107  2.7439617672
L_PTL_B2|_RX|RB1 _PTL_B2|_RX|101 0  2.38752113364072e-12
L_PTL_B2|_RX|RB2 _PTL_B2|_RX|104 0  1.937922998085e-12
L_PTL_B2|_RX|RB3 _PTL_B2|_RX|107 0  1.550338398468e-12
B_PTL_B2|_JTL|1 _PTL_B2|_JTL|1 _PTL_B2|_JTL|2 JJMIT AREA=2.5
B_PTL_B2|_JTL|2 _PTL_B2|_JTL|6 _PTL_B2|_JTL|7 JJMIT AREA=2.5
I_PTL_B2|_JTL|B1 0 _PTL_B2|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B2|_JTL|1 _PTL_B2|A_PTL_RX _PTL_B2|_JTL|1  2.067833848e-12
L_PTL_B2|_JTL|2 _PTL_B2|_JTL|1 _PTL_B2|_JTL|4  2.067833848e-12
L_PTL_B2|_JTL|3 _PTL_B2|_JTL|4 _PTL_B2|_JTL|6  2.067833848e-12
L_PTL_B2|_JTL|4 _PTL_B2|_JTL|6 B2_RX  2.067833848e-12
L_PTL_B2|_JTL|P1 _PTL_B2|_JTL|2 0  2e-13
L_PTL_B2|_JTL|P2 _PTL_B2|_JTL|7 0  2e-13
L_PTL_B2|_JTL|B1 _PTL_B2|_JTL|5 _PTL_B2|_JTL|4  2e-12
R_PTL_B2|_JTL|B1 _PTL_B2|_JTL|1 _PTL_B2|_JTL|3  2.7439617672
R_PTL_B2|_JTL|B2 _PTL_B2|_JTL|6 _PTL_B2|_JTL|8  2.7439617672
L_PTL_B2|_JTL|RB1 _PTL_B2|_JTL|3 0  1.750338398468e-12
L_PTL_B2|_JTL|RB2 _PTL_B2|_JTL|8 0  1.750338398468e-12
B_PTL_A3|_TX|1 _PTL_A3|_TX|1 _PTL_A3|_TX|2 JJMIT AREA=2.5
B_PTL_A3|_TX|2 _PTL_A3|_TX|4 _PTL_A3|_TX|5 JJMIT AREA=2.5
I_PTL_A3|_TX|B1 0 _PTL_A3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A3|_TX|B2 0 _PTL_A3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|3  1.684e-12
L_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|6  3.596e-12
L_PTL_A3|_TX|1 A3_TX _PTL_A3|_TX|1  2.063e-12
L_PTL_A3|_TX|2 _PTL_A3|_TX|1 _PTL_A3|_TX|4  4.123e-12
L_PTL_A3|_TX|3 _PTL_A3|_TX|4 _PTL_A3|_TX|7  2.193e-12
R_PTL_A3|_TX|D _PTL_A3|_TX|7 _PTL_A3|A_PTL  1.36
L_PTL_A3|_TX|P1 _PTL_A3|_TX|2 0  5.254e-13
L_PTL_A3|_TX|P2 _PTL_A3|_TX|5 0  5.141e-13
R_PTL_A3|_TX|B1 _PTL_A3|_TX|1 _PTL_A3|_TX|101  2.7439617672
R_PTL_A3|_TX|B2 _PTL_A3|_TX|4 _PTL_A3|_TX|104  2.7439617672
L_PTL_A3|_TX|RB1 _PTL_A3|_TX|101 0  1.550338398468e-12
L_PTL_A3|_TX|RB2 _PTL_A3|_TX|104 0  1.550338398468e-12
B_PTL_A3|_RX|1 _PTL_A3|_RX|1 _PTL_A3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A3|_RX|2 _PTL_A3|_RX|4 _PTL_A3|_RX|5 JJMIT AREA=2.0
B_PTL_A3|_RX|3 _PTL_A3|_RX|7 _PTL_A3|_RX|8 JJMIT AREA=2.5
I_PTL_A3|_RX|B1 0 _PTL_A3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|3  2.777e-12
I_PTL_A3|_RX|B2 0 _PTL_A3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|6  2.685e-12
I_PTL_A3|_RX|B3 0 _PTL_A3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|9  2.764e-12
L_PTL_A3|_RX|1 _PTL_A3|A_PTL _PTL_A3|_RX|1  1.346e-12
L_PTL_A3|_RX|2 _PTL_A3|_RX|1 _PTL_A3|_RX|4  6.348e-12
L_PTL_A3|_RX|3 _PTL_A3|_RX|4 _PTL_A3|_RX|7  5.197e-12
L_PTL_A3|_RX|4 _PTL_A3|_RX|7 _PTL_A3|A_PTL_RX  2.058e-12
L_PTL_A3|_RX|P1 _PTL_A3|_RX|2 0  4.795e-13
L_PTL_A3|_RX|P2 _PTL_A3|_RX|5 0  5.431e-13
L_PTL_A3|_RX|P3 _PTL_A3|_RX|8 0  5.339e-13
R_PTL_A3|_RX|B1 _PTL_A3|_RX|1 _PTL_A3|_RX|101  4.225701121488
R_PTL_A3|_RX|B2 _PTL_A3|_RX|4 _PTL_A3|_RX|104  3.429952209
R_PTL_A3|_RX|B3 _PTL_A3|_RX|7 _PTL_A3|_RX|107  2.7439617672
L_PTL_A3|_RX|RB1 _PTL_A3|_RX|101 0  2.38752113364072e-12
L_PTL_A3|_RX|RB2 _PTL_A3|_RX|104 0  1.937922998085e-12
L_PTL_A3|_RX|RB3 _PTL_A3|_RX|107 0  1.550338398468e-12
B_PTL_A3|_JTL|1 _PTL_A3|_JTL|1 _PTL_A3|_JTL|2 JJMIT AREA=2.5
B_PTL_A3|_JTL|2 _PTL_A3|_JTL|6 _PTL_A3|_JTL|7 JJMIT AREA=2.5
I_PTL_A3|_JTL|B1 0 _PTL_A3|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A3|_JTL|1 _PTL_A3|A_PTL_RX _PTL_A3|_JTL|1  2.067833848e-12
L_PTL_A3|_JTL|2 _PTL_A3|_JTL|1 _PTL_A3|_JTL|4  2.067833848e-12
L_PTL_A3|_JTL|3 _PTL_A3|_JTL|4 _PTL_A3|_JTL|6  2.067833848e-12
L_PTL_A3|_JTL|4 _PTL_A3|_JTL|6 A3_RX  2.067833848e-12
L_PTL_A3|_JTL|P1 _PTL_A3|_JTL|2 0  2e-13
L_PTL_A3|_JTL|P2 _PTL_A3|_JTL|7 0  2e-13
L_PTL_A3|_JTL|B1 _PTL_A3|_JTL|5 _PTL_A3|_JTL|4  2e-12
R_PTL_A3|_JTL|B1 _PTL_A3|_JTL|1 _PTL_A3|_JTL|3  2.7439617672
R_PTL_A3|_JTL|B2 _PTL_A3|_JTL|6 _PTL_A3|_JTL|8  2.7439617672
L_PTL_A3|_JTL|RB1 _PTL_A3|_JTL|3 0  1.750338398468e-12
L_PTL_A3|_JTL|RB2 _PTL_A3|_JTL|8 0  1.750338398468e-12
B_PTL_B3|_TX|1 _PTL_B3|_TX|1 _PTL_B3|_TX|2 JJMIT AREA=2.5
B_PTL_B3|_TX|2 _PTL_B3|_TX|4 _PTL_B3|_TX|5 JJMIT AREA=2.5
I_PTL_B3|_TX|B1 0 _PTL_B3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B3|_TX|B2 0 _PTL_B3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|3  1.684e-12
L_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|6  3.596e-12
L_PTL_B3|_TX|1 B3_TX _PTL_B3|_TX|1  2.063e-12
L_PTL_B3|_TX|2 _PTL_B3|_TX|1 _PTL_B3|_TX|4  4.123e-12
L_PTL_B3|_TX|3 _PTL_B3|_TX|4 _PTL_B3|_TX|7  2.193e-12
R_PTL_B3|_TX|D _PTL_B3|_TX|7 _PTL_B3|A_PTL  1.36
L_PTL_B3|_TX|P1 _PTL_B3|_TX|2 0  5.254e-13
L_PTL_B3|_TX|P2 _PTL_B3|_TX|5 0  5.141e-13
R_PTL_B3|_TX|B1 _PTL_B3|_TX|1 _PTL_B3|_TX|101  2.7439617672
R_PTL_B3|_TX|B2 _PTL_B3|_TX|4 _PTL_B3|_TX|104  2.7439617672
L_PTL_B3|_TX|RB1 _PTL_B3|_TX|101 0  1.550338398468e-12
L_PTL_B3|_TX|RB2 _PTL_B3|_TX|104 0  1.550338398468e-12
B_PTL_B3|_RX|1 _PTL_B3|_RX|1 _PTL_B3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B3|_RX|2 _PTL_B3|_RX|4 _PTL_B3|_RX|5 JJMIT AREA=2.0
B_PTL_B3|_RX|3 _PTL_B3|_RX|7 _PTL_B3|_RX|8 JJMIT AREA=2.5
I_PTL_B3|_RX|B1 0 _PTL_B3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|3  2.777e-12
I_PTL_B3|_RX|B2 0 _PTL_B3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|6  2.685e-12
I_PTL_B3|_RX|B3 0 _PTL_B3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|9  2.764e-12
L_PTL_B3|_RX|1 _PTL_B3|A_PTL _PTL_B3|_RX|1  1.346e-12
L_PTL_B3|_RX|2 _PTL_B3|_RX|1 _PTL_B3|_RX|4  6.348e-12
L_PTL_B3|_RX|3 _PTL_B3|_RX|4 _PTL_B3|_RX|7  5.197e-12
L_PTL_B3|_RX|4 _PTL_B3|_RX|7 _PTL_B3|A_PTL_RX  2.058e-12
L_PTL_B3|_RX|P1 _PTL_B3|_RX|2 0  4.795e-13
L_PTL_B3|_RX|P2 _PTL_B3|_RX|5 0  5.431e-13
L_PTL_B3|_RX|P3 _PTL_B3|_RX|8 0  5.339e-13
R_PTL_B3|_RX|B1 _PTL_B3|_RX|1 _PTL_B3|_RX|101  4.225701121488
R_PTL_B3|_RX|B2 _PTL_B3|_RX|4 _PTL_B3|_RX|104  3.429952209
R_PTL_B3|_RX|B3 _PTL_B3|_RX|7 _PTL_B3|_RX|107  2.7439617672
L_PTL_B3|_RX|RB1 _PTL_B3|_RX|101 0  2.38752113364072e-12
L_PTL_B3|_RX|RB2 _PTL_B3|_RX|104 0  1.937922998085e-12
L_PTL_B3|_RX|RB3 _PTL_B3|_RX|107 0  1.550338398468e-12
B_PTL_B3|_JTL|1 _PTL_B3|_JTL|1 _PTL_B3|_JTL|2 JJMIT AREA=2.5
B_PTL_B3|_JTL|2 _PTL_B3|_JTL|6 _PTL_B3|_JTL|7 JJMIT AREA=2.5
I_PTL_B3|_JTL|B1 0 _PTL_B3|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B3|_JTL|1 _PTL_B3|A_PTL_RX _PTL_B3|_JTL|1  2.067833848e-12
L_PTL_B3|_JTL|2 _PTL_B3|_JTL|1 _PTL_B3|_JTL|4  2.067833848e-12
L_PTL_B3|_JTL|3 _PTL_B3|_JTL|4 _PTL_B3|_JTL|6  2.067833848e-12
L_PTL_B3|_JTL|4 _PTL_B3|_JTL|6 B3_RX  2.067833848e-12
L_PTL_B3|_JTL|P1 _PTL_B3|_JTL|2 0  2e-13
L_PTL_B3|_JTL|P2 _PTL_B3|_JTL|7 0  2e-13
L_PTL_B3|_JTL|B1 _PTL_B3|_JTL|5 _PTL_B3|_JTL|4  2e-12
R_PTL_B3|_JTL|B1 _PTL_B3|_JTL|1 _PTL_B3|_JTL|3  2.7439617672
R_PTL_B3|_JTL|B2 _PTL_B3|_JTL|6 _PTL_B3|_JTL|8  2.7439617672
L_PTL_B3|_JTL|RB1 _PTL_B3|_JTL|3 0  1.750338398468e-12
L_PTL_B3|_JTL|RB2 _PTL_B3|_JTL|8 0  1.750338398468e-12
B_PTL_A4|_TX|1 _PTL_A4|_TX|1 _PTL_A4|_TX|2 JJMIT AREA=2.5
B_PTL_A4|_TX|2 _PTL_A4|_TX|4 _PTL_A4|_TX|5 JJMIT AREA=2.5
I_PTL_A4|_TX|B1 0 _PTL_A4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A4|_TX|B2 0 _PTL_A4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A4|_TX|B1 _PTL_A4|_TX|1 _PTL_A4|_TX|3  1.684e-12
L_PTL_A4|_TX|B2 _PTL_A4|_TX|4 _PTL_A4|_TX|6  3.596e-12
L_PTL_A4|_TX|1 A4_TX _PTL_A4|_TX|1  2.063e-12
L_PTL_A4|_TX|2 _PTL_A4|_TX|1 _PTL_A4|_TX|4  4.123e-12
L_PTL_A4|_TX|3 _PTL_A4|_TX|4 _PTL_A4|_TX|7  2.193e-12
R_PTL_A4|_TX|D _PTL_A4|_TX|7 _PTL_A4|A_PTL  1.36
L_PTL_A4|_TX|P1 _PTL_A4|_TX|2 0  5.254e-13
L_PTL_A4|_TX|P2 _PTL_A4|_TX|5 0  5.141e-13
R_PTL_A4|_TX|B1 _PTL_A4|_TX|1 _PTL_A4|_TX|101  2.7439617672
R_PTL_A4|_TX|B2 _PTL_A4|_TX|4 _PTL_A4|_TX|104  2.7439617672
L_PTL_A4|_TX|RB1 _PTL_A4|_TX|101 0  1.550338398468e-12
L_PTL_A4|_TX|RB2 _PTL_A4|_TX|104 0  1.550338398468e-12
B_PTL_A4|_RX|1 _PTL_A4|_RX|1 _PTL_A4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A4|_RX|2 _PTL_A4|_RX|4 _PTL_A4|_RX|5 JJMIT AREA=2.0
B_PTL_A4|_RX|3 _PTL_A4|_RX|7 _PTL_A4|_RX|8 JJMIT AREA=2.5
I_PTL_A4|_RX|B1 0 _PTL_A4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A4|_RX|B1 _PTL_A4|_RX|1 _PTL_A4|_RX|3  2.777e-12
I_PTL_A4|_RX|B2 0 _PTL_A4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A4|_RX|B2 _PTL_A4|_RX|4 _PTL_A4|_RX|6  2.685e-12
I_PTL_A4|_RX|B3 0 _PTL_A4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A4|_RX|B3 _PTL_A4|_RX|7 _PTL_A4|_RX|9  2.764e-12
L_PTL_A4|_RX|1 _PTL_A4|A_PTL _PTL_A4|_RX|1  1.346e-12
L_PTL_A4|_RX|2 _PTL_A4|_RX|1 _PTL_A4|_RX|4  6.348e-12
L_PTL_A4|_RX|3 _PTL_A4|_RX|4 _PTL_A4|_RX|7  5.197e-12
L_PTL_A4|_RX|4 _PTL_A4|_RX|7 _PTL_A4|A_PTL_RX  2.058e-12
L_PTL_A4|_RX|P1 _PTL_A4|_RX|2 0  4.795e-13
L_PTL_A4|_RX|P2 _PTL_A4|_RX|5 0  5.431e-13
L_PTL_A4|_RX|P3 _PTL_A4|_RX|8 0  5.339e-13
R_PTL_A4|_RX|B1 _PTL_A4|_RX|1 _PTL_A4|_RX|101  4.225701121488
R_PTL_A4|_RX|B2 _PTL_A4|_RX|4 _PTL_A4|_RX|104  3.429952209
R_PTL_A4|_RX|B3 _PTL_A4|_RX|7 _PTL_A4|_RX|107  2.7439617672
L_PTL_A4|_RX|RB1 _PTL_A4|_RX|101 0  2.38752113364072e-12
L_PTL_A4|_RX|RB2 _PTL_A4|_RX|104 0  1.937922998085e-12
L_PTL_A4|_RX|RB3 _PTL_A4|_RX|107 0  1.550338398468e-12
B_PTL_A4|_JTL|1 _PTL_A4|_JTL|1 _PTL_A4|_JTL|2 JJMIT AREA=2.5
B_PTL_A4|_JTL|2 _PTL_A4|_JTL|6 _PTL_A4|_JTL|7 JJMIT AREA=2.5
I_PTL_A4|_JTL|B1 0 _PTL_A4|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A4|_JTL|1 _PTL_A4|A_PTL_RX _PTL_A4|_JTL|1  2.067833848e-12
L_PTL_A4|_JTL|2 _PTL_A4|_JTL|1 _PTL_A4|_JTL|4  2.067833848e-12
L_PTL_A4|_JTL|3 _PTL_A4|_JTL|4 _PTL_A4|_JTL|6  2.067833848e-12
L_PTL_A4|_JTL|4 _PTL_A4|_JTL|6 A4_RX  2.067833848e-12
L_PTL_A4|_JTL|P1 _PTL_A4|_JTL|2 0  2e-13
L_PTL_A4|_JTL|P2 _PTL_A4|_JTL|7 0  2e-13
L_PTL_A4|_JTL|B1 _PTL_A4|_JTL|5 _PTL_A4|_JTL|4  2e-12
R_PTL_A4|_JTL|B1 _PTL_A4|_JTL|1 _PTL_A4|_JTL|3  2.7439617672
R_PTL_A4|_JTL|B2 _PTL_A4|_JTL|6 _PTL_A4|_JTL|8  2.7439617672
L_PTL_A4|_JTL|RB1 _PTL_A4|_JTL|3 0  1.750338398468e-12
L_PTL_A4|_JTL|RB2 _PTL_A4|_JTL|8 0  1.750338398468e-12
B_PTL_B4|_TX|1 _PTL_B4|_TX|1 _PTL_B4|_TX|2 JJMIT AREA=2.5
B_PTL_B4|_TX|2 _PTL_B4|_TX|4 _PTL_B4|_TX|5 JJMIT AREA=2.5
I_PTL_B4|_TX|B1 0 _PTL_B4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B4|_TX|B2 0 _PTL_B4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B4|_TX|B1 _PTL_B4|_TX|1 _PTL_B4|_TX|3  1.684e-12
L_PTL_B4|_TX|B2 _PTL_B4|_TX|4 _PTL_B4|_TX|6  3.596e-12
L_PTL_B4|_TX|1 B4_TX _PTL_B4|_TX|1  2.063e-12
L_PTL_B4|_TX|2 _PTL_B4|_TX|1 _PTL_B4|_TX|4  4.123e-12
L_PTL_B4|_TX|3 _PTL_B4|_TX|4 _PTL_B4|_TX|7  2.193e-12
R_PTL_B4|_TX|D _PTL_B4|_TX|7 _PTL_B4|A_PTL  1.36
L_PTL_B4|_TX|P1 _PTL_B4|_TX|2 0  5.254e-13
L_PTL_B4|_TX|P2 _PTL_B4|_TX|5 0  5.141e-13
R_PTL_B4|_TX|B1 _PTL_B4|_TX|1 _PTL_B4|_TX|101  2.7439617672
R_PTL_B4|_TX|B2 _PTL_B4|_TX|4 _PTL_B4|_TX|104  2.7439617672
L_PTL_B4|_TX|RB1 _PTL_B4|_TX|101 0  1.550338398468e-12
L_PTL_B4|_TX|RB2 _PTL_B4|_TX|104 0  1.550338398468e-12
B_PTL_B4|_RX|1 _PTL_B4|_RX|1 _PTL_B4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B4|_RX|2 _PTL_B4|_RX|4 _PTL_B4|_RX|5 JJMIT AREA=2.0
B_PTL_B4|_RX|3 _PTL_B4|_RX|7 _PTL_B4|_RX|8 JJMIT AREA=2.5
I_PTL_B4|_RX|B1 0 _PTL_B4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B4|_RX|B1 _PTL_B4|_RX|1 _PTL_B4|_RX|3  2.777e-12
I_PTL_B4|_RX|B2 0 _PTL_B4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B4|_RX|B2 _PTL_B4|_RX|4 _PTL_B4|_RX|6  2.685e-12
I_PTL_B4|_RX|B3 0 _PTL_B4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B4|_RX|B3 _PTL_B4|_RX|7 _PTL_B4|_RX|9  2.764e-12
L_PTL_B4|_RX|1 _PTL_B4|A_PTL _PTL_B4|_RX|1  1.346e-12
L_PTL_B4|_RX|2 _PTL_B4|_RX|1 _PTL_B4|_RX|4  6.348e-12
L_PTL_B4|_RX|3 _PTL_B4|_RX|4 _PTL_B4|_RX|7  5.197e-12
L_PTL_B4|_RX|4 _PTL_B4|_RX|7 _PTL_B4|A_PTL_RX  2.058e-12
L_PTL_B4|_RX|P1 _PTL_B4|_RX|2 0  4.795e-13
L_PTL_B4|_RX|P2 _PTL_B4|_RX|5 0  5.431e-13
L_PTL_B4|_RX|P3 _PTL_B4|_RX|8 0  5.339e-13
R_PTL_B4|_RX|B1 _PTL_B4|_RX|1 _PTL_B4|_RX|101  4.225701121488
R_PTL_B4|_RX|B2 _PTL_B4|_RX|4 _PTL_B4|_RX|104  3.429952209
R_PTL_B4|_RX|B3 _PTL_B4|_RX|7 _PTL_B4|_RX|107  2.7439617672
L_PTL_B4|_RX|RB1 _PTL_B4|_RX|101 0  2.38752113364072e-12
L_PTL_B4|_RX|RB2 _PTL_B4|_RX|104 0  1.937922998085e-12
L_PTL_B4|_RX|RB3 _PTL_B4|_RX|107 0  1.550338398468e-12
B_PTL_B4|_JTL|1 _PTL_B4|_JTL|1 _PTL_B4|_JTL|2 JJMIT AREA=2.5
B_PTL_B4|_JTL|2 _PTL_B4|_JTL|6 _PTL_B4|_JTL|7 JJMIT AREA=2.5
I_PTL_B4|_JTL|B1 0 _PTL_B4|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B4|_JTL|1 _PTL_B4|A_PTL_RX _PTL_B4|_JTL|1  2.067833848e-12
L_PTL_B4|_JTL|2 _PTL_B4|_JTL|1 _PTL_B4|_JTL|4  2.067833848e-12
L_PTL_B4|_JTL|3 _PTL_B4|_JTL|4 _PTL_B4|_JTL|6  2.067833848e-12
L_PTL_B4|_JTL|4 _PTL_B4|_JTL|6 B4_RX  2.067833848e-12
L_PTL_B4|_JTL|P1 _PTL_B4|_JTL|2 0  2e-13
L_PTL_B4|_JTL|P2 _PTL_B4|_JTL|7 0  2e-13
L_PTL_B4|_JTL|B1 _PTL_B4|_JTL|5 _PTL_B4|_JTL|4  2e-12
R_PTL_B4|_JTL|B1 _PTL_B4|_JTL|1 _PTL_B4|_JTL|3  2.7439617672
R_PTL_B4|_JTL|B2 _PTL_B4|_JTL|6 _PTL_B4|_JTL|8  2.7439617672
L_PTL_B4|_JTL|RB1 _PTL_B4|_JTL|3 0  1.750338398468e-12
L_PTL_B4|_JTL|RB2 _PTL_B4|_JTL|8 0  1.750338398468e-12
B_PTL_A5|_TX|1 _PTL_A5|_TX|1 _PTL_A5|_TX|2 JJMIT AREA=2.5
B_PTL_A5|_TX|2 _PTL_A5|_TX|4 _PTL_A5|_TX|5 JJMIT AREA=2.5
I_PTL_A5|_TX|B1 0 _PTL_A5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A5|_TX|B2 0 _PTL_A5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A5|_TX|B1 _PTL_A5|_TX|1 _PTL_A5|_TX|3  1.684e-12
L_PTL_A5|_TX|B2 _PTL_A5|_TX|4 _PTL_A5|_TX|6  3.596e-12
L_PTL_A5|_TX|1 A5_TX _PTL_A5|_TX|1  2.063e-12
L_PTL_A5|_TX|2 _PTL_A5|_TX|1 _PTL_A5|_TX|4  4.123e-12
L_PTL_A5|_TX|3 _PTL_A5|_TX|4 _PTL_A5|_TX|7  2.193e-12
R_PTL_A5|_TX|D _PTL_A5|_TX|7 _PTL_A5|A_PTL  1.36
L_PTL_A5|_TX|P1 _PTL_A5|_TX|2 0  5.254e-13
L_PTL_A5|_TX|P2 _PTL_A5|_TX|5 0  5.141e-13
R_PTL_A5|_TX|B1 _PTL_A5|_TX|1 _PTL_A5|_TX|101  2.7439617672
R_PTL_A5|_TX|B2 _PTL_A5|_TX|4 _PTL_A5|_TX|104  2.7439617672
L_PTL_A5|_TX|RB1 _PTL_A5|_TX|101 0  1.550338398468e-12
L_PTL_A5|_TX|RB2 _PTL_A5|_TX|104 0  1.550338398468e-12
B_PTL_A5|_RX|1 _PTL_A5|_RX|1 _PTL_A5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A5|_RX|2 _PTL_A5|_RX|4 _PTL_A5|_RX|5 JJMIT AREA=2.0
B_PTL_A5|_RX|3 _PTL_A5|_RX|7 _PTL_A5|_RX|8 JJMIT AREA=2.5
I_PTL_A5|_RX|B1 0 _PTL_A5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A5|_RX|B1 _PTL_A5|_RX|1 _PTL_A5|_RX|3  2.777e-12
I_PTL_A5|_RX|B2 0 _PTL_A5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A5|_RX|B2 _PTL_A5|_RX|4 _PTL_A5|_RX|6  2.685e-12
I_PTL_A5|_RX|B3 0 _PTL_A5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A5|_RX|B3 _PTL_A5|_RX|7 _PTL_A5|_RX|9  2.764e-12
L_PTL_A5|_RX|1 _PTL_A5|A_PTL _PTL_A5|_RX|1  1.346e-12
L_PTL_A5|_RX|2 _PTL_A5|_RX|1 _PTL_A5|_RX|4  6.348e-12
L_PTL_A5|_RX|3 _PTL_A5|_RX|4 _PTL_A5|_RX|7  5.197e-12
L_PTL_A5|_RX|4 _PTL_A5|_RX|7 _PTL_A5|A_PTL_RX  2.058e-12
L_PTL_A5|_RX|P1 _PTL_A5|_RX|2 0  4.795e-13
L_PTL_A5|_RX|P2 _PTL_A5|_RX|5 0  5.431e-13
L_PTL_A5|_RX|P3 _PTL_A5|_RX|8 0  5.339e-13
R_PTL_A5|_RX|B1 _PTL_A5|_RX|1 _PTL_A5|_RX|101  4.225701121488
R_PTL_A5|_RX|B2 _PTL_A5|_RX|4 _PTL_A5|_RX|104  3.429952209
R_PTL_A5|_RX|B3 _PTL_A5|_RX|7 _PTL_A5|_RX|107  2.7439617672
L_PTL_A5|_RX|RB1 _PTL_A5|_RX|101 0  2.38752113364072e-12
L_PTL_A5|_RX|RB2 _PTL_A5|_RX|104 0  1.937922998085e-12
L_PTL_A5|_RX|RB3 _PTL_A5|_RX|107 0  1.550338398468e-12
B_PTL_A5|_JTL|1 _PTL_A5|_JTL|1 _PTL_A5|_JTL|2 JJMIT AREA=2.5
B_PTL_A5|_JTL|2 _PTL_A5|_JTL|6 _PTL_A5|_JTL|7 JJMIT AREA=2.5
I_PTL_A5|_JTL|B1 0 _PTL_A5|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A5|_JTL|1 _PTL_A5|A_PTL_RX _PTL_A5|_JTL|1  2.067833848e-12
L_PTL_A5|_JTL|2 _PTL_A5|_JTL|1 _PTL_A5|_JTL|4  2.067833848e-12
L_PTL_A5|_JTL|3 _PTL_A5|_JTL|4 _PTL_A5|_JTL|6  2.067833848e-12
L_PTL_A5|_JTL|4 _PTL_A5|_JTL|6 A5_RX  2.067833848e-12
L_PTL_A5|_JTL|P1 _PTL_A5|_JTL|2 0  2e-13
L_PTL_A5|_JTL|P2 _PTL_A5|_JTL|7 0  2e-13
L_PTL_A5|_JTL|B1 _PTL_A5|_JTL|5 _PTL_A5|_JTL|4  2e-12
R_PTL_A5|_JTL|B1 _PTL_A5|_JTL|1 _PTL_A5|_JTL|3  2.7439617672
R_PTL_A5|_JTL|B2 _PTL_A5|_JTL|6 _PTL_A5|_JTL|8  2.7439617672
L_PTL_A5|_JTL|RB1 _PTL_A5|_JTL|3 0  1.750338398468e-12
L_PTL_A5|_JTL|RB2 _PTL_A5|_JTL|8 0  1.750338398468e-12
B_PTL_B5|_TX|1 _PTL_B5|_TX|1 _PTL_B5|_TX|2 JJMIT AREA=2.5
B_PTL_B5|_TX|2 _PTL_B5|_TX|4 _PTL_B5|_TX|5 JJMIT AREA=2.5
I_PTL_B5|_TX|B1 0 _PTL_B5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B5|_TX|B2 0 _PTL_B5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B5|_TX|B1 _PTL_B5|_TX|1 _PTL_B5|_TX|3  1.684e-12
L_PTL_B5|_TX|B2 _PTL_B5|_TX|4 _PTL_B5|_TX|6  3.596e-12
L_PTL_B5|_TX|1 B5_TX _PTL_B5|_TX|1  2.063e-12
L_PTL_B5|_TX|2 _PTL_B5|_TX|1 _PTL_B5|_TX|4  4.123e-12
L_PTL_B5|_TX|3 _PTL_B5|_TX|4 _PTL_B5|_TX|7  2.193e-12
R_PTL_B5|_TX|D _PTL_B5|_TX|7 _PTL_B5|A_PTL  1.36
L_PTL_B5|_TX|P1 _PTL_B5|_TX|2 0  5.254e-13
L_PTL_B5|_TX|P2 _PTL_B5|_TX|5 0  5.141e-13
R_PTL_B5|_TX|B1 _PTL_B5|_TX|1 _PTL_B5|_TX|101  2.7439617672
R_PTL_B5|_TX|B2 _PTL_B5|_TX|4 _PTL_B5|_TX|104  2.7439617672
L_PTL_B5|_TX|RB1 _PTL_B5|_TX|101 0  1.550338398468e-12
L_PTL_B5|_TX|RB2 _PTL_B5|_TX|104 0  1.550338398468e-12
B_PTL_B5|_RX|1 _PTL_B5|_RX|1 _PTL_B5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B5|_RX|2 _PTL_B5|_RX|4 _PTL_B5|_RX|5 JJMIT AREA=2.0
B_PTL_B5|_RX|3 _PTL_B5|_RX|7 _PTL_B5|_RX|8 JJMIT AREA=2.5
I_PTL_B5|_RX|B1 0 _PTL_B5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B5|_RX|B1 _PTL_B5|_RX|1 _PTL_B5|_RX|3  2.777e-12
I_PTL_B5|_RX|B2 0 _PTL_B5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B5|_RX|B2 _PTL_B5|_RX|4 _PTL_B5|_RX|6  2.685e-12
I_PTL_B5|_RX|B3 0 _PTL_B5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B5|_RX|B3 _PTL_B5|_RX|7 _PTL_B5|_RX|9  2.764e-12
L_PTL_B5|_RX|1 _PTL_B5|A_PTL _PTL_B5|_RX|1  1.346e-12
L_PTL_B5|_RX|2 _PTL_B5|_RX|1 _PTL_B5|_RX|4  6.348e-12
L_PTL_B5|_RX|3 _PTL_B5|_RX|4 _PTL_B5|_RX|7  5.197e-12
L_PTL_B5|_RX|4 _PTL_B5|_RX|7 _PTL_B5|A_PTL_RX  2.058e-12
L_PTL_B5|_RX|P1 _PTL_B5|_RX|2 0  4.795e-13
L_PTL_B5|_RX|P2 _PTL_B5|_RX|5 0  5.431e-13
L_PTL_B5|_RX|P3 _PTL_B5|_RX|8 0  5.339e-13
R_PTL_B5|_RX|B1 _PTL_B5|_RX|1 _PTL_B5|_RX|101  4.225701121488
R_PTL_B5|_RX|B2 _PTL_B5|_RX|4 _PTL_B5|_RX|104  3.429952209
R_PTL_B5|_RX|B3 _PTL_B5|_RX|7 _PTL_B5|_RX|107  2.7439617672
L_PTL_B5|_RX|RB1 _PTL_B5|_RX|101 0  2.38752113364072e-12
L_PTL_B5|_RX|RB2 _PTL_B5|_RX|104 0  1.937922998085e-12
L_PTL_B5|_RX|RB3 _PTL_B5|_RX|107 0  1.550338398468e-12
B_PTL_B5|_JTL|1 _PTL_B5|_JTL|1 _PTL_B5|_JTL|2 JJMIT AREA=2.5
B_PTL_B5|_JTL|2 _PTL_B5|_JTL|6 _PTL_B5|_JTL|7 JJMIT AREA=2.5
I_PTL_B5|_JTL|B1 0 _PTL_B5|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B5|_JTL|1 _PTL_B5|A_PTL_RX _PTL_B5|_JTL|1  2.067833848e-12
L_PTL_B5|_JTL|2 _PTL_B5|_JTL|1 _PTL_B5|_JTL|4  2.067833848e-12
L_PTL_B5|_JTL|3 _PTL_B5|_JTL|4 _PTL_B5|_JTL|6  2.067833848e-12
L_PTL_B5|_JTL|4 _PTL_B5|_JTL|6 B5_RX  2.067833848e-12
L_PTL_B5|_JTL|P1 _PTL_B5|_JTL|2 0  2e-13
L_PTL_B5|_JTL|P2 _PTL_B5|_JTL|7 0  2e-13
L_PTL_B5|_JTL|B1 _PTL_B5|_JTL|5 _PTL_B5|_JTL|4  2e-12
R_PTL_B5|_JTL|B1 _PTL_B5|_JTL|1 _PTL_B5|_JTL|3  2.7439617672
R_PTL_B5|_JTL|B2 _PTL_B5|_JTL|6 _PTL_B5|_JTL|8  2.7439617672
L_PTL_B5|_JTL|RB1 _PTL_B5|_JTL|3 0  1.750338398468e-12
L_PTL_B5|_JTL|RB2 _PTL_B5|_JTL|8 0  1.750338398468e-12
B_PTL_A6|_TX|1 _PTL_A6|_TX|1 _PTL_A6|_TX|2 JJMIT AREA=2.5
B_PTL_A6|_TX|2 _PTL_A6|_TX|4 _PTL_A6|_TX|5 JJMIT AREA=2.5
I_PTL_A6|_TX|B1 0 _PTL_A6|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A6|_TX|B2 0 _PTL_A6|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A6|_TX|B1 _PTL_A6|_TX|1 _PTL_A6|_TX|3  1.684e-12
L_PTL_A6|_TX|B2 _PTL_A6|_TX|4 _PTL_A6|_TX|6  3.596e-12
L_PTL_A6|_TX|1 A6_TX _PTL_A6|_TX|1  2.063e-12
L_PTL_A6|_TX|2 _PTL_A6|_TX|1 _PTL_A6|_TX|4  4.123e-12
L_PTL_A6|_TX|3 _PTL_A6|_TX|4 _PTL_A6|_TX|7  2.193e-12
R_PTL_A6|_TX|D _PTL_A6|_TX|7 _PTL_A6|A_PTL  1.36
L_PTL_A6|_TX|P1 _PTL_A6|_TX|2 0  5.254e-13
L_PTL_A6|_TX|P2 _PTL_A6|_TX|5 0  5.141e-13
R_PTL_A6|_TX|B1 _PTL_A6|_TX|1 _PTL_A6|_TX|101  2.7439617672
R_PTL_A6|_TX|B2 _PTL_A6|_TX|4 _PTL_A6|_TX|104  2.7439617672
L_PTL_A6|_TX|RB1 _PTL_A6|_TX|101 0  1.550338398468e-12
L_PTL_A6|_TX|RB2 _PTL_A6|_TX|104 0  1.550338398468e-12
B_PTL_A6|_RX|1 _PTL_A6|_RX|1 _PTL_A6|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A6|_RX|2 _PTL_A6|_RX|4 _PTL_A6|_RX|5 JJMIT AREA=2.0
B_PTL_A6|_RX|3 _PTL_A6|_RX|7 _PTL_A6|_RX|8 JJMIT AREA=2.5
I_PTL_A6|_RX|B1 0 _PTL_A6|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A6|_RX|B1 _PTL_A6|_RX|1 _PTL_A6|_RX|3  2.777e-12
I_PTL_A6|_RX|B2 0 _PTL_A6|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A6|_RX|B2 _PTL_A6|_RX|4 _PTL_A6|_RX|6  2.685e-12
I_PTL_A6|_RX|B3 0 _PTL_A6|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A6|_RX|B3 _PTL_A6|_RX|7 _PTL_A6|_RX|9  2.764e-12
L_PTL_A6|_RX|1 _PTL_A6|A_PTL _PTL_A6|_RX|1  1.346e-12
L_PTL_A6|_RX|2 _PTL_A6|_RX|1 _PTL_A6|_RX|4  6.348e-12
L_PTL_A6|_RX|3 _PTL_A6|_RX|4 _PTL_A6|_RX|7  5.197e-12
L_PTL_A6|_RX|4 _PTL_A6|_RX|7 _PTL_A6|A_PTL_RX  2.058e-12
L_PTL_A6|_RX|P1 _PTL_A6|_RX|2 0  4.795e-13
L_PTL_A6|_RX|P2 _PTL_A6|_RX|5 0  5.431e-13
L_PTL_A6|_RX|P3 _PTL_A6|_RX|8 0  5.339e-13
R_PTL_A6|_RX|B1 _PTL_A6|_RX|1 _PTL_A6|_RX|101  4.225701121488
R_PTL_A6|_RX|B2 _PTL_A6|_RX|4 _PTL_A6|_RX|104  3.429952209
R_PTL_A6|_RX|B3 _PTL_A6|_RX|7 _PTL_A6|_RX|107  2.7439617672
L_PTL_A6|_RX|RB1 _PTL_A6|_RX|101 0  2.38752113364072e-12
L_PTL_A6|_RX|RB2 _PTL_A6|_RX|104 0  1.937922998085e-12
L_PTL_A6|_RX|RB3 _PTL_A6|_RX|107 0  1.550338398468e-12
B_PTL_A6|_JTL|1 _PTL_A6|_JTL|1 _PTL_A6|_JTL|2 JJMIT AREA=2.5
B_PTL_A6|_JTL|2 _PTL_A6|_JTL|6 _PTL_A6|_JTL|7 JJMIT AREA=2.5
I_PTL_A6|_JTL|B1 0 _PTL_A6|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A6|_JTL|1 _PTL_A6|A_PTL_RX _PTL_A6|_JTL|1  2.067833848e-12
L_PTL_A6|_JTL|2 _PTL_A6|_JTL|1 _PTL_A6|_JTL|4  2.067833848e-12
L_PTL_A6|_JTL|3 _PTL_A6|_JTL|4 _PTL_A6|_JTL|6  2.067833848e-12
L_PTL_A6|_JTL|4 _PTL_A6|_JTL|6 A6_RX  2.067833848e-12
L_PTL_A6|_JTL|P1 _PTL_A6|_JTL|2 0  2e-13
L_PTL_A6|_JTL|P2 _PTL_A6|_JTL|7 0  2e-13
L_PTL_A6|_JTL|B1 _PTL_A6|_JTL|5 _PTL_A6|_JTL|4  2e-12
R_PTL_A6|_JTL|B1 _PTL_A6|_JTL|1 _PTL_A6|_JTL|3  2.7439617672
R_PTL_A6|_JTL|B2 _PTL_A6|_JTL|6 _PTL_A6|_JTL|8  2.7439617672
L_PTL_A6|_JTL|RB1 _PTL_A6|_JTL|3 0  1.750338398468e-12
L_PTL_A6|_JTL|RB2 _PTL_A6|_JTL|8 0  1.750338398468e-12
B_PTL_B6|_TX|1 _PTL_B6|_TX|1 _PTL_B6|_TX|2 JJMIT AREA=2.5
B_PTL_B6|_TX|2 _PTL_B6|_TX|4 _PTL_B6|_TX|5 JJMIT AREA=2.5
I_PTL_B6|_TX|B1 0 _PTL_B6|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B6|_TX|B2 0 _PTL_B6|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B6|_TX|B1 _PTL_B6|_TX|1 _PTL_B6|_TX|3  1.684e-12
L_PTL_B6|_TX|B2 _PTL_B6|_TX|4 _PTL_B6|_TX|6  3.596e-12
L_PTL_B6|_TX|1 B6_TX _PTL_B6|_TX|1  2.063e-12
L_PTL_B6|_TX|2 _PTL_B6|_TX|1 _PTL_B6|_TX|4  4.123e-12
L_PTL_B6|_TX|3 _PTL_B6|_TX|4 _PTL_B6|_TX|7  2.193e-12
R_PTL_B6|_TX|D _PTL_B6|_TX|7 _PTL_B6|A_PTL  1.36
L_PTL_B6|_TX|P1 _PTL_B6|_TX|2 0  5.254e-13
L_PTL_B6|_TX|P2 _PTL_B6|_TX|5 0  5.141e-13
R_PTL_B6|_TX|B1 _PTL_B6|_TX|1 _PTL_B6|_TX|101  2.7439617672
R_PTL_B6|_TX|B2 _PTL_B6|_TX|4 _PTL_B6|_TX|104  2.7439617672
L_PTL_B6|_TX|RB1 _PTL_B6|_TX|101 0  1.550338398468e-12
L_PTL_B6|_TX|RB2 _PTL_B6|_TX|104 0  1.550338398468e-12
B_PTL_B6|_RX|1 _PTL_B6|_RX|1 _PTL_B6|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B6|_RX|2 _PTL_B6|_RX|4 _PTL_B6|_RX|5 JJMIT AREA=2.0
B_PTL_B6|_RX|3 _PTL_B6|_RX|7 _PTL_B6|_RX|8 JJMIT AREA=2.5
I_PTL_B6|_RX|B1 0 _PTL_B6|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B6|_RX|B1 _PTL_B6|_RX|1 _PTL_B6|_RX|3  2.777e-12
I_PTL_B6|_RX|B2 0 _PTL_B6|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B6|_RX|B2 _PTL_B6|_RX|4 _PTL_B6|_RX|6  2.685e-12
I_PTL_B6|_RX|B3 0 _PTL_B6|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B6|_RX|B3 _PTL_B6|_RX|7 _PTL_B6|_RX|9  2.764e-12
L_PTL_B6|_RX|1 _PTL_B6|A_PTL _PTL_B6|_RX|1  1.346e-12
L_PTL_B6|_RX|2 _PTL_B6|_RX|1 _PTL_B6|_RX|4  6.348e-12
L_PTL_B6|_RX|3 _PTL_B6|_RX|4 _PTL_B6|_RX|7  5.197e-12
L_PTL_B6|_RX|4 _PTL_B6|_RX|7 _PTL_B6|A_PTL_RX  2.058e-12
L_PTL_B6|_RX|P1 _PTL_B6|_RX|2 0  4.795e-13
L_PTL_B6|_RX|P2 _PTL_B6|_RX|5 0  5.431e-13
L_PTL_B6|_RX|P3 _PTL_B6|_RX|8 0  5.339e-13
R_PTL_B6|_RX|B1 _PTL_B6|_RX|1 _PTL_B6|_RX|101  4.225701121488
R_PTL_B6|_RX|B2 _PTL_B6|_RX|4 _PTL_B6|_RX|104  3.429952209
R_PTL_B6|_RX|B3 _PTL_B6|_RX|7 _PTL_B6|_RX|107  2.7439617672
L_PTL_B6|_RX|RB1 _PTL_B6|_RX|101 0  2.38752113364072e-12
L_PTL_B6|_RX|RB2 _PTL_B6|_RX|104 0  1.937922998085e-12
L_PTL_B6|_RX|RB3 _PTL_B6|_RX|107 0  1.550338398468e-12
B_PTL_B6|_JTL|1 _PTL_B6|_JTL|1 _PTL_B6|_JTL|2 JJMIT AREA=2.5
B_PTL_B6|_JTL|2 _PTL_B6|_JTL|6 _PTL_B6|_JTL|7 JJMIT AREA=2.5
I_PTL_B6|_JTL|B1 0 _PTL_B6|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B6|_JTL|1 _PTL_B6|A_PTL_RX _PTL_B6|_JTL|1  2.067833848e-12
L_PTL_B6|_JTL|2 _PTL_B6|_JTL|1 _PTL_B6|_JTL|4  2.067833848e-12
L_PTL_B6|_JTL|3 _PTL_B6|_JTL|4 _PTL_B6|_JTL|6  2.067833848e-12
L_PTL_B6|_JTL|4 _PTL_B6|_JTL|6 B6_RX  2.067833848e-12
L_PTL_B6|_JTL|P1 _PTL_B6|_JTL|2 0  2e-13
L_PTL_B6|_JTL|P2 _PTL_B6|_JTL|7 0  2e-13
L_PTL_B6|_JTL|B1 _PTL_B6|_JTL|5 _PTL_B6|_JTL|4  2e-12
R_PTL_B6|_JTL|B1 _PTL_B6|_JTL|1 _PTL_B6|_JTL|3  2.7439617672
R_PTL_B6|_JTL|B2 _PTL_B6|_JTL|6 _PTL_B6|_JTL|8  2.7439617672
L_PTL_B6|_JTL|RB1 _PTL_B6|_JTL|3 0  1.750338398468e-12
L_PTL_B6|_JTL|RB2 _PTL_B6|_JTL|8 0  1.750338398468e-12
B_PTL_A7|_TX|1 _PTL_A7|_TX|1 _PTL_A7|_TX|2 JJMIT AREA=2.5
B_PTL_A7|_TX|2 _PTL_A7|_TX|4 _PTL_A7|_TX|5 JJMIT AREA=2.5
I_PTL_A7|_TX|B1 0 _PTL_A7|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_A7|_TX|B2 0 _PTL_A7|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_A7|_TX|B1 _PTL_A7|_TX|1 _PTL_A7|_TX|3  1.684e-12
L_PTL_A7|_TX|B2 _PTL_A7|_TX|4 _PTL_A7|_TX|6  3.596e-12
L_PTL_A7|_TX|1 A7_TX _PTL_A7|_TX|1  2.063e-12
L_PTL_A7|_TX|2 _PTL_A7|_TX|1 _PTL_A7|_TX|4  4.123e-12
L_PTL_A7|_TX|3 _PTL_A7|_TX|4 _PTL_A7|_TX|7  2.193e-12
R_PTL_A7|_TX|D _PTL_A7|_TX|7 _PTL_A7|A_PTL  1.36
L_PTL_A7|_TX|P1 _PTL_A7|_TX|2 0  5.254e-13
L_PTL_A7|_TX|P2 _PTL_A7|_TX|5 0  5.141e-13
R_PTL_A7|_TX|B1 _PTL_A7|_TX|1 _PTL_A7|_TX|101  2.7439617672
R_PTL_A7|_TX|B2 _PTL_A7|_TX|4 _PTL_A7|_TX|104  2.7439617672
L_PTL_A7|_TX|RB1 _PTL_A7|_TX|101 0  1.550338398468e-12
L_PTL_A7|_TX|RB2 _PTL_A7|_TX|104 0  1.550338398468e-12
B_PTL_A7|_RX|1 _PTL_A7|_RX|1 _PTL_A7|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_A7|_RX|2 _PTL_A7|_RX|4 _PTL_A7|_RX|5 JJMIT AREA=2.0
B_PTL_A7|_RX|3 _PTL_A7|_RX|7 _PTL_A7|_RX|8 JJMIT AREA=2.5
I_PTL_A7|_RX|B1 0 _PTL_A7|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_A7|_RX|B1 _PTL_A7|_RX|1 _PTL_A7|_RX|3  2.777e-12
I_PTL_A7|_RX|B2 0 _PTL_A7|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_A7|_RX|B2 _PTL_A7|_RX|4 _PTL_A7|_RX|6  2.685e-12
I_PTL_A7|_RX|B3 0 _PTL_A7|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_A7|_RX|B3 _PTL_A7|_RX|7 _PTL_A7|_RX|9  2.764e-12
L_PTL_A7|_RX|1 _PTL_A7|A_PTL _PTL_A7|_RX|1  1.346e-12
L_PTL_A7|_RX|2 _PTL_A7|_RX|1 _PTL_A7|_RX|4  6.348e-12
L_PTL_A7|_RX|3 _PTL_A7|_RX|4 _PTL_A7|_RX|7  5.197e-12
L_PTL_A7|_RX|4 _PTL_A7|_RX|7 _PTL_A7|A_PTL_RX  2.058e-12
L_PTL_A7|_RX|P1 _PTL_A7|_RX|2 0  4.795e-13
L_PTL_A7|_RX|P2 _PTL_A7|_RX|5 0  5.431e-13
L_PTL_A7|_RX|P3 _PTL_A7|_RX|8 0  5.339e-13
R_PTL_A7|_RX|B1 _PTL_A7|_RX|1 _PTL_A7|_RX|101  4.225701121488
R_PTL_A7|_RX|B2 _PTL_A7|_RX|4 _PTL_A7|_RX|104  3.429952209
R_PTL_A7|_RX|B3 _PTL_A7|_RX|7 _PTL_A7|_RX|107  2.7439617672
L_PTL_A7|_RX|RB1 _PTL_A7|_RX|101 0  2.38752113364072e-12
L_PTL_A7|_RX|RB2 _PTL_A7|_RX|104 0  1.937922998085e-12
L_PTL_A7|_RX|RB3 _PTL_A7|_RX|107 0  1.550338398468e-12
B_PTL_A7|_JTL|1 _PTL_A7|_JTL|1 _PTL_A7|_JTL|2 JJMIT AREA=2.5
B_PTL_A7|_JTL|2 _PTL_A7|_JTL|6 _PTL_A7|_JTL|7 JJMIT AREA=2.5
I_PTL_A7|_JTL|B1 0 _PTL_A7|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_A7|_JTL|1 _PTL_A7|A_PTL_RX _PTL_A7|_JTL|1  2.067833848e-12
L_PTL_A7|_JTL|2 _PTL_A7|_JTL|1 _PTL_A7|_JTL|4  2.067833848e-12
L_PTL_A7|_JTL|3 _PTL_A7|_JTL|4 _PTL_A7|_JTL|6  2.067833848e-12
L_PTL_A7|_JTL|4 _PTL_A7|_JTL|6 A7_RX  2.067833848e-12
L_PTL_A7|_JTL|P1 _PTL_A7|_JTL|2 0  2e-13
L_PTL_A7|_JTL|P2 _PTL_A7|_JTL|7 0  2e-13
L_PTL_A7|_JTL|B1 _PTL_A7|_JTL|5 _PTL_A7|_JTL|4  2e-12
R_PTL_A7|_JTL|B1 _PTL_A7|_JTL|1 _PTL_A7|_JTL|3  2.7439617672
R_PTL_A7|_JTL|B2 _PTL_A7|_JTL|6 _PTL_A7|_JTL|8  2.7439617672
L_PTL_A7|_JTL|RB1 _PTL_A7|_JTL|3 0  1.750338398468e-12
L_PTL_A7|_JTL|RB2 _PTL_A7|_JTL|8 0  1.750338398468e-12
B_PTL_B7|_TX|1 _PTL_B7|_TX|1 _PTL_B7|_TX|2 JJMIT AREA=2.5
B_PTL_B7|_TX|2 _PTL_B7|_TX|4 _PTL_B7|_TX|5 JJMIT AREA=2.5
I_PTL_B7|_TX|B1 0 _PTL_B7|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_B7|_TX|B2 0 _PTL_B7|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_B7|_TX|B1 _PTL_B7|_TX|1 _PTL_B7|_TX|3  1.684e-12
L_PTL_B7|_TX|B2 _PTL_B7|_TX|4 _PTL_B7|_TX|6  3.596e-12
L_PTL_B7|_TX|1 B7_TX _PTL_B7|_TX|1  2.063e-12
L_PTL_B7|_TX|2 _PTL_B7|_TX|1 _PTL_B7|_TX|4  4.123e-12
L_PTL_B7|_TX|3 _PTL_B7|_TX|4 _PTL_B7|_TX|7  2.193e-12
R_PTL_B7|_TX|D _PTL_B7|_TX|7 _PTL_B7|A_PTL  1.36
L_PTL_B7|_TX|P1 _PTL_B7|_TX|2 0  5.254e-13
L_PTL_B7|_TX|P2 _PTL_B7|_TX|5 0  5.141e-13
R_PTL_B7|_TX|B1 _PTL_B7|_TX|1 _PTL_B7|_TX|101  2.7439617672
R_PTL_B7|_TX|B2 _PTL_B7|_TX|4 _PTL_B7|_TX|104  2.7439617672
L_PTL_B7|_TX|RB1 _PTL_B7|_TX|101 0  1.550338398468e-12
L_PTL_B7|_TX|RB2 _PTL_B7|_TX|104 0  1.550338398468e-12
B_PTL_B7|_RX|1 _PTL_B7|_RX|1 _PTL_B7|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_B7|_RX|2 _PTL_B7|_RX|4 _PTL_B7|_RX|5 JJMIT AREA=2.0
B_PTL_B7|_RX|3 _PTL_B7|_RX|7 _PTL_B7|_RX|8 JJMIT AREA=2.5
I_PTL_B7|_RX|B1 0 _PTL_B7|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_B7|_RX|B1 _PTL_B7|_RX|1 _PTL_B7|_RX|3  2.777e-12
I_PTL_B7|_RX|B2 0 _PTL_B7|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_B7|_RX|B2 _PTL_B7|_RX|4 _PTL_B7|_RX|6  2.685e-12
I_PTL_B7|_RX|B3 0 _PTL_B7|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_B7|_RX|B3 _PTL_B7|_RX|7 _PTL_B7|_RX|9  2.764e-12
L_PTL_B7|_RX|1 _PTL_B7|A_PTL _PTL_B7|_RX|1  1.346e-12
L_PTL_B7|_RX|2 _PTL_B7|_RX|1 _PTL_B7|_RX|4  6.348e-12
L_PTL_B7|_RX|3 _PTL_B7|_RX|4 _PTL_B7|_RX|7  5.197e-12
L_PTL_B7|_RX|4 _PTL_B7|_RX|7 _PTL_B7|A_PTL_RX  2.058e-12
L_PTL_B7|_RX|P1 _PTL_B7|_RX|2 0  4.795e-13
L_PTL_B7|_RX|P2 _PTL_B7|_RX|5 0  5.431e-13
L_PTL_B7|_RX|P3 _PTL_B7|_RX|8 0  5.339e-13
R_PTL_B7|_RX|B1 _PTL_B7|_RX|1 _PTL_B7|_RX|101  4.225701121488
R_PTL_B7|_RX|B2 _PTL_B7|_RX|4 _PTL_B7|_RX|104  3.429952209
R_PTL_B7|_RX|B3 _PTL_B7|_RX|7 _PTL_B7|_RX|107  2.7439617672
L_PTL_B7|_RX|RB1 _PTL_B7|_RX|101 0  2.38752113364072e-12
L_PTL_B7|_RX|RB2 _PTL_B7|_RX|104 0  1.937922998085e-12
L_PTL_B7|_RX|RB3 _PTL_B7|_RX|107 0  1.550338398468e-12
B_PTL_B7|_JTL|1 _PTL_B7|_JTL|1 _PTL_B7|_JTL|2 JJMIT AREA=2.5
B_PTL_B7|_JTL|2 _PTL_B7|_JTL|6 _PTL_B7|_JTL|7 JJMIT AREA=2.5
I_PTL_B7|_JTL|B1 0 _PTL_B7|_JTL|5  PWL(0 0 5e-12 0.00035)
L_PTL_B7|_JTL|1 _PTL_B7|A_PTL_RX _PTL_B7|_JTL|1  2.067833848e-12
L_PTL_B7|_JTL|2 _PTL_B7|_JTL|1 _PTL_B7|_JTL|4  2.067833848e-12
L_PTL_B7|_JTL|3 _PTL_B7|_JTL|4 _PTL_B7|_JTL|6  2.067833848e-12
L_PTL_B7|_JTL|4 _PTL_B7|_JTL|6 B7_RX  2.067833848e-12
L_PTL_B7|_JTL|P1 _PTL_B7|_JTL|2 0  2e-13
L_PTL_B7|_JTL|P2 _PTL_B7|_JTL|7 0  2e-13
L_PTL_B7|_JTL|B1 _PTL_B7|_JTL|5 _PTL_B7|_JTL|4  2e-12
R_PTL_B7|_JTL|B1 _PTL_B7|_JTL|1 _PTL_B7|_JTL|3  2.7439617672
R_PTL_B7|_JTL|B2 _PTL_B7|_JTL|6 _PTL_B7|_JTL|8  2.7439617672
L_PTL_B7|_JTL|RB1 _PTL_B7|_JTL|3 0  1.750338398468e-12
L_PTL_B7|_JTL|RB2 _PTL_B7|_JTL|8 0  1.750338398468e-12
LI0|_SPL_A|1 A0_RX I0|_SPL_A|D1  2e-12
LI0|_SPL_A|2 I0|_SPL_A|D1 I0|_SPL_A|D2  4.135667696e-12
LI0|_SPL_A|3 I0|_SPL_A|D2 I0|_SPL_A|JCT  9.84682784761905e-13
LI0|_SPL_A|4 I0|_SPL_A|JCT I0|_SPL_A|QA1  9.84682784761905e-13
LI0|_SPL_A|5 I0|_SPL_A|QA1 I0|A1  2e-12
LI0|_SPL_A|6 I0|_SPL_A|JCT I0|_SPL_A|QB1  9.84682784761905e-13
LI0|_SPL_A|7 I0|_SPL_A|QB1 I0|A2  2e-12
LI0|_SPL_B|1 B0_RX I0|_SPL_B|D1  2e-12
LI0|_SPL_B|2 I0|_SPL_B|D1 I0|_SPL_B|D2  4.135667696e-12
LI0|_SPL_B|3 I0|_SPL_B|D2 I0|_SPL_B|JCT  9.84682784761905e-13
LI0|_SPL_B|4 I0|_SPL_B|JCT I0|_SPL_B|QA1  9.84682784761905e-13
LI0|_SPL_B|5 I0|_SPL_B|QA1 I0|B1  2e-12
LI0|_SPL_B|6 I0|_SPL_B|JCT I0|_SPL_B|QB1  9.84682784761905e-13
LI0|_SPL_B|7 I0|_SPL_B|QB1 I0|B2  2e-12
LI0|_DFF_A|1 I0|A1 I0|_DFF_A|A1  2.067833848e-12
LI0|_DFF_A|2 I0|_DFF_A|A1 I0|_DFF_A|A2  4.135667696e-12
LI0|_DFF_A|3 I0|_DFF_A|A3 I0|_DFF_A|A4  8.271335392e-12
LI0|_DFF_A|T T00 I0|_DFF_A|T1  2.067833848e-12
LI0|_DFF_A|4 I0|_DFF_A|T1 I0|_DFF_A|T2  4.135667696e-12
LI0|_DFF_A|5 I0|_DFF_A|A4 I0|_DFF_A|Q1  4.135667696e-12
LI0|_DFF_A|6 I0|_DFF_A|Q1 I0|A1_SYNC  2.067833848e-12
LI0|_DFF_B|1 I0|B1 I0|_DFF_B|A1  2.067833848e-12
LI0|_DFF_B|2 I0|_DFF_B|A1 I0|_DFF_B|A2  4.135667696e-12
LI0|_DFF_B|3 I0|_DFF_B|A3 I0|_DFF_B|A4  8.271335392e-12
LI0|_DFF_B|T T00 I0|_DFF_B|T1  2.067833848e-12
LI0|_DFF_B|4 I0|_DFF_B|T1 I0|_DFF_B|T2  4.135667696e-12
LI0|_DFF_B|5 I0|_DFF_B|A4 I0|_DFF_B|Q1  4.135667696e-12
LI0|_DFF_B|6 I0|_DFF_B|Q1 I0|B1_SYNC  2.067833848e-12
LI0|_XOR|A1 I0|A2 I0|_XOR|A1  2.067833848e-12
LI0|_XOR|A2 I0|_XOR|A1 I0|_XOR|A2  4.135667696e-12
LI0|_XOR|A3 I0|_XOR|A3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|B1 I0|B2 I0|_XOR|B1  2.067833848e-12
LI0|_XOR|B2 I0|_XOR|B1 I0|_XOR|B2  4.135667696e-12
LI0|_XOR|B3 I0|_XOR|B3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|T1 T00 I0|_XOR|T1  2.067833848e-12
LI0|_XOR|T2 I0|_XOR|T1 I0|_XOR|T2  4.135667696e-12
LI0|_XOR|Q2 I0|_XOR|ABTQ I0|_XOR|Q1  4.135667696e-12
LI0|_XOR|Q1 I0|_XOR|Q1 IP0_0  2.067833848e-12
LI0|_AND|A1 I0|A1_SYNC I0|_AND|A1  2.067833848e-12
LI0|_AND|A2 I0|_AND|A1 I0|_AND|A2  4.135667696e-12
LI0|_AND|A3 I0|_AND|A3 I0|_AND|Q3  1.2e-12
LI0|_AND|B1 I0|B1_SYNC I0|_AND|B1  2.067833848e-12
LI0|_AND|B2 I0|_AND|B1 I0|_AND|B2  4.135667696e-12
LI0|_AND|B3 I0|_AND|B3 I0|_AND|Q3  1.2e-12
LI0|_AND|Q3 I0|_AND|Q3 I0|_AND|Q2  4.135667696e-12
LI0|_AND|Q2 I0|_AND|Q2 I0|_AND|Q1  4.135667696e-12
LI0|_AND|Q1 I0|_AND|Q1 IG0_0  2.067833848e-12
LI1|_SPL_A|1 A1_RX I1|_SPL_A|D1  2e-12
LI1|_SPL_A|2 I1|_SPL_A|D1 I1|_SPL_A|D2  4.135667696e-12
LI1|_SPL_A|3 I1|_SPL_A|D2 I1|_SPL_A|JCT  9.84682784761905e-13
LI1|_SPL_A|4 I1|_SPL_A|JCT I1|_SPL_A|QA1  9.84682784761905e-13
LI1|_SPL_A|5 I1|_SPL_A|QA1 I1|A1  2e-12
LI1|_SPL_A|6 I1|_SPL_A|JCT I1|_SPL_A|QB1  9.84682784761905e-13
LI1|_SPL_A|7 I1|_SPL_A|QB1 I1|A2  2e-12
LI1|_SPL_B|1 B1_RX I1|_SPL_B|D1  2e-12
LI1|_SPL_B|2 I1|_SPL_B|D1 I1|_SPL_B|D2  4.135667696e-12
LI1|_SPL_B|3 I1|_SPL_B|D2 I1|_SPL_B|JCT  9.84682784761905e-13
LI1|_SPL_B|4 I1|_SPL_B|JCT I1|_SPL_B|QA1  9.84682784761905e-13
LI1|_SPL_B|5 I1|_SPL_B|QA1 I1|B1  2e-12
LI1|_SPL_B|6 I1|_SPL_B|JCT I1|_SPL_B|QB1  9.84682784761905e-13
LI1|_SPL_B|7 I1|_SPL_B|QB1 I1|B2  2e-12
LI1|_DFF_A|1 I1|A1 I1|_DFF_A|A1  2.067833848e-12
LI1|_DFF_A|2 I1|_DFF_A|A1 I1|_DFF_A|A2  4.135667696e-12
LI1|_DFF_A|3 I1|_DFF_A|A3 I1|_DFF_A|A4  8.271335392e-12
LI1|_DFF_A|T T01 I1|_DFF_A|T1  2.067833848e-12
LI1|_DFF_A|4 I1|_DFF_A|T1 I1|_DFF_A|T2  4.135667696e-12
LI1|_DFF_A|5 I1|_DFF_A|A4 I1|_DFF_A|Q1  4.135667696e-12
LI1|_DFF_A|6 I1|_DFF_A|Q1 I1|A1_SYNC  2.067833848e-12
LI1|_DFF_B|1 I1|B1 I1|_DFF_B|A1  2.067833848e-12
LI1|_DFF_B|2 I1|_DFF_B|A1 I1|_DFF_B|A2  4.135667696e-12
LI1|_DFF_B|3 I1|_DFF_B|A3 I1|_DFF_B|A4  8.271335392e-12
LI1|_DFF_B|T T01 I1|_DFF_B|T1  2.067833848e-12
LI1|_DFF_B|4 I1|_DFF_B|T1 I1|_DFF_B|T2  4.135667696e-12
LI1|_DFF_B|5 I1|_DFF_B|A4 I1|_DFF_B|Q1  4.135667696e-12
LI1|_DFF_B|6 I1|_DFF_B|Q1 I1|B1_SYNC  2.067833848e-12
LI1|_XOR|A1 I1|A2 I1|_XOR|A1  2.067833848e-12
LI1|_XOR|A2 I1|_XOR|A1 I1|_XOR|A2  4.135667696e-12
LI1|_XOR|A3 I1|_XOR|A3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|B1 I1|B2 I1|_XOR|B1  2.067833848e-12
LI1|_XOR|B2 I1|_XOR|B1 I1|_XOR|B2  4.135667696e-12
LI1|_XOR|B3 I1|_XOR|B3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|T1 T01 I1|_XOR|T1  2.067833848e-12
LI1|_XOR|T2 I1|_XOR|T1 I1|_XOR|T2  4.135667696e-12
LI1|_XOR|Q2 I1|_XOR|ABTQ I1|_XOR|Q1  4.135667696e-12
LI1|_XOR|Q1 I1|_XOR|Q1 IP1_0  2.067833848e-12
LI1|_AND|A1 I1|A1_SYNC I1|_AND|A1  2.067833848e-12
LI1|_AND|A2 I1|_AND|A1 I1|_AND|A2  4.135667696e-12
LI1|_AND|A3 I1|_AND|A3 I1|_AND|Q3  1.2e-12
LI1|_AND|B1 I1|B1_SYNC I1|_AND|B1  2.067833848e-12
LI1|_AND|B2 I1|_AND|B1 I1|_AND|B2  4.135667696e-12
LI1|_AND|B3 I1|_AND|B3 I1|_AND|Q3  1.2e-12
LI1|_AND|Q3 I1|_AND|Q3 I1|_AND|Q2  4.135667696e-12
LI1|_AND|Q2 I1|_AND|Q2 I1|_AND|Q1  4.135667696e-12
LI1|_AND|Q1 I1|_AND|Q1 IG1_0  2.067833848e-12
LI2|_SPL_A|1 A2_RX I2|_SPL_A|D1  2e-12
LI2|_SPL_A|2 I2|_SPL_A|D1 I2|_SPL_A|D2  4.135667696e-12
LI2|_SPL_A|3 I2|_SPL_A|D2 I2|_SPL_A|JCT  9.84682784761905e-13
LI2|_SPL_A|4 I2|_SPL_A|JCT I2|_SPL_A|QA1  9.84682784761905e-13
LI2|_SPL_A|5 I2|_SPL_A|QA1 I2|A1  2e-12
LI2|_SPL_A|6 I2|_SPL_A|JCT I2|_SPL_A|QB1  9.84682784761905e-13
LI2|_SPL_A|7 I2|_SPL_A|QB1 I2|A2  2e-12
LI2|_SPL_B|1 B2_RX I2|_SPL_B|D1  2e-12
LI2|_SPL_B|2 I2|_SPL_B|D1 I2|_SPL_B|D2  4.135667696e-12
LI2|_SPL_B|3 I2|_SPL_B|D2 I2|_SPL_B|JCT  9.84682784761905e-13
LI2|_SPL_B|4 I2|_SPL_B|JCT I2|_SPL_B|QA1  9.84682784761905e-13
LI2|_SPL_B|5 I2|_SPL_B|QA1 I2|B1  2e-12
LI2|_SPL_B|6 I2|_SPL_B|JCT I2|_SPL_B|QB1  9.84682784761905e-13
LI2|_SPL_B|7 I2|_SPL_B|QB1 I2|B2  2e-12
LI2|_DFF_A|1 I2|A1 I2|_DFF_A|A1  2.067833848e-12
LI2|_DFF_A|2 I2|_DFF_A|A1 I2|_DFF_A|A2  4.135667696e-12
LI2|_DFF_A|3 I2|_DFF_A|A3 I2|_DFF_A|A4  8.271335392e-12
LI2|_DFF_A|T T02 I2|_DFF_A|T1  2.067833848e-12
LI2|_DFF_A|4 I2|_DFF_A|T1 I2|_DFF_A|T2  4.135667696e-12
LI2|_DFF_A|5 I2|_DFF_A|A4 I2|_DFF_A|Q1  4.135667696e-12
LI2|_DFF_A|6 I2|_DFF_A|Q1 I2|A1_SYNC  2.067833848e-12
LI2|_DFF_B|1 I2|B1 I2|_DFF_B|A1  2.067833848e-12
LI2|_DFF_B|2 I2|_DFF_B|A1 I2|_DFF_B|A2  4.135667696e-12
LI2|_DFF_B|3 I2|_DFF_B|A3 I2|_DFF_B|A4  8.271335392e-12
LI2|_DFF_B|T T02 I2|_DFF_B|T1  2.067833848e-12
LI2|_DFF_B|4 I2|_DFF_B|T1 I2|_DFF_B|T2  4.135667696e-12
LI2|_DFF_B|5 I2|_DFF_B|A4 I2|_DFF_B|Q1  4.135667696e-12
LI2|_DFF_B|6 I2|_DFF_B|Q1 I2|B1_SYNC  2.067833848e-12
LI2|_XOR|A1 I2|A2 I2|_XOR|A1  2.067833848e-12
LI2|_XOR|A2 I2|_XOR|A1 I2|_XOR|A2  4.135667696e-12
LI2|_XOR|A3 I2|_XOR|A3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|B1 I2|B2 I2|_XOR|B1  2.067833848e-12
LI2|_XOR|B2 I2|_XOR|B1 I2|_XOR|B2  4.135667696e-12
LI2|_XOR|B3 I2|_XOR|B3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|T1 T02 I2|_XOR|T1  2.067833848e-12
LI2|_XOR|T2 I2|_XOR|T1 I2|_XOR|T2  4.135667696e-12
LI2|_XOR|Q2 I2|_XOR|ABTQ I2|_XOR|Q1  4.135667696e-12
LI2|_XOR|Q1 I2|_XOR|Q1 IP2_0  2.067833848e-12
LI2|_AND|A1 I2|A1_SYNC I2|_AND|A1  2.067833848e-12
LI2|_AND|A2 I2|_AND|A1 I2|_AND|A2  4.135667696e-12
LI2|_AND|A3 I2|_AND|A3 I2|_AND|Q3  1.2e-12
LI2|_AND|B1 I2|B1_SYNC I2|_AND|B1  2.067833848e-12
LI2|_AND|B2 I2|_AND|B1 I2|_AND|B2  4.135667696e-12
LI2|_AND|B3 I2|_AND|B3 I2|_AND|Q3  1.2e-12
LI2|_AND|Q3 I2|_AND|Q3 I2|_AND|Q2  4.135667696e-12
LI2|_AND|Q2 I2|_AND|Q2 I2|_AND|Q1  4.135667696e-12
LI2|_AND|Q1 I2|_AND|Q1 IG2_0  2.067833848e-12
LI3|_SPL_A|1 A3_RX I3|_SPL_A|D1  2e-12
LI3|_SPL_A|2 I3|_SPL_A|D1 I3|_SPL_A|D2  4.135667696e-12
LI3|_SPL_A|3 I3|_SPL_A|D2 I3|_SPL_A|JCT  9.84682784761905e-13
LI3|_SPL_A|4 I3|_SPL_A|JCT I3|_SPL_A|QA1  9.84682784761905e-13
LI3|_SPL_A|5 I3|_SPL_A|QA1 I3|A1  2e-12
LI3|_SPL_A|6 I3|_SPL_A|JCT I3|_SPL_A|QB1  9.84682784761905e-13
LI3|_SPL_A|7 I3|_SPL_A|QB1 I3|A2  2e-12
LI3|_SPL_B|1 B3_RX I3|_SPL_B|D1  2e-12
LI3|_SPL_B|2 I3|_SPL_B|D1 I3|_SPL_B|D2  4.135667696e-12
LI3|_SPL_B|3 I3|_SPL_B|D2 I3|_SPL_B|JCT  9.84682784761905e-13
LI3|_SPL_B|4 I3|_SPL_B|JCT I3|_SPL_B|QA1  9.84682784761905e-13
LI3|_SPL_B|5 I3|_SPL_B|QA1 I3|B1  2e-12
LI3|_SPL_B|6 I3|_SPL_B|JCT I3|_SPL_B|QB1  9.84682784761905e-13
LI3|_SPL_B|7 I3|_SPL_B|QB1 I3|B2  2e-12
LI3|_DFF_A|1 I3|A1 I3|_DFF_A|A1  2.067833848e-12
LI3|_DFF_A|2 I3|_DFF_A|A1 I3|_DFF_A|A2  4.135667696e-12
LI3|_DFF_A|3 I3|_DFF_A|A3 I3|_DFF_A|A4  8.271335392e-12
LI3|_DFF_A|T T03 I3|_DFF_A|T1  2.067833848e-12
LI3|_DFF_A|4 I3|_DFF_A|T1 I3|_DFF_A|T2  4.135667696e-12
LI3|_DFF_A|5 I3|_DFF_A|A4 I3|_DFF_A|Q1  4.135667696e-12
LI3|_DFF_A|6 I3|_DFF_A|Q1 I3|A1_SYNC  2.067833848e-12
LI3|_DFF_B|1 I3|B1 I3|_DFF_B|A1  2.067833848e-12
LI3|_DFF_B|2 I3|_DFF_B|A1 I3|_DFF_B|A2  4.135667696e-12
LI3|_DFF_B|3 I3|_DFF_B|A3 I3|_DFF_B|A4  8.271335392e-12
LI3|_DFF_B|T T03 I3|_DFF_B|T1  2.067833848e-12
LI3|_DFF_B|4 I3|_DFF_B|T1 I3|_DFF_B|T2  4.135667696e-12
LI3|_DFF_B|5 I3|_DFF_B|A4 I3|_DFF_B|Q1  4.135667696e-12
LI3|_DFF_B|6 I3|_DFF_B|Q1 I3|B1_SYNC  2.067833848e-12
LI3|_XOR|A1 I3|A2 I3|_XOR|A1  2.067833848e-12
LI3|_XOR|A2 I3|_XOR|A1 I3|_XOR|A2  4.135667696e-12
LI3|_XOR|A3 I3|_XOR|A3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|B1 I3|B2 I3|_XOR|B1  2.067833848e-12
LI3|_XOR|B2 I3|_XOR|B1 I3|_XOR|B2  4.135667696e-12
LI3|_XOR|B3 I3|_XOR|B3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|T1 T03 I3|_XOR|T1  2.067833848e-12
LI3|_XOR|T2 I3|_XOR|T1 I3|_XOR|T2  4.135667696e-12
LI3|_XOR|Q2 I3|_XOR|ABTQ I3|_XOR|Q1  4.135667696e-12
LI3|_XOR|Q1 I3|_XOR|Q1 IP3_0  2.067833848e-12
LI3|_AND|A1 I3|A1_SYNC I3|_AND|A1  2.067833848e-12
LI3|_AND|A2 I3|_AND|A1 I3|_AND|A2  4.135667696e-12
LI3|_AND|A3 I3|_AND|A3 I3|_AND|Q3  1.2e-12
LI3|_AND|B1 I3|B1_SYNC I3|_AND|B1  2.067833848e-12
LI3|_AND|B2 I3|_AND|B1 I3|_AND|B2  4.135667696e-12
LI3|_AND|B3 I3|_AND|B3 I3|_AND|Q3  1.2e-12
LI3|_AND|Q3 I3|_AND|Q3 I3|_AND|Q2  4.135667696e-12
LI3|_AND|Q2 I3|_AND|Q2 I3|_AND|Q1  4.135667696e-12
LI3|_AND|Q1 I3|_AND|Q1 IG3_0  2.067833848e-12
LI4|_SPL_A|1 A4_RX I4|_SPL_A|D1  2e-12
LI4|_SPL_A|2 I4|_SPL_A|D1 I4|_SPL_A|D2  4.135667696e-12
LI4|_SPL_A|3 I4|_SPL_A|D2 I4|_SPL_A|JCT  9.84682784761905e-13
LI4|_SPL_A|4 I4|_SPL_A|JCT I4|_SPL_A|QA1  9.84682784761905e-13
LI4|_SPL_A|5 I4|_SPL_A|QA1 I4|A1  2e-12
LI4|_SPL_A|6 I4|_SPL_A|JCT I4|_SPL_A|QB1  9.84682784761905e-13
LI4|_SPL_A|7 I4|_SPL_A|QB1 I4|A2  2e-12
LI4|_SPL_B|1 B4_RX I4|_SPL_B|D1  2e-12
LI4|_SPL_B|2 I4|_SPL_B|D1 I4|_SPL_B|D2  4.135667696e-12
LI4|_SPL_B|3 I4|_SPL_B|D2 I4|_SPL_B|JCT  9.84682784761905e-13
LI4|_SPL_B|4 I4|_SPL_B|JCT I4|_SPL_B|QA1  9.84682784761905e-13
LI4|_SPL_B|5 I4|_SPL_B|QA1 I4|B1  2e-12
LI4|_SPL_B|6 I4|_SPL_B|JCT I4|_SPL_B|QB1  9.84682784761905e-13
LI4|_SPL_B|7 I4|_SPL_B|QB1 I4|B2  2e-12
LI4|_DFF_A|1 I4|A1 I4|_DFF_A|A1  2.067833848e-12
LI4|_DFF_A|2 I4|_DFF_A|A1 I4|_DFF_A|A2  4.135667696e-12
LI4|_DFF_A|3 I4|_DFF_A|A3 I4|_DFF_A|A4  8.271335392e-12
LI4|_DFF_A|T T04 I4|_DFF_A|T1  2.067833848e-12
LI4|_DFF_A|4 I4|_DFF_A|T1 I4|_DFF_A|T2  4.135667696e-12
LI4|_DFF_A|5 I4|_DFF_A|A4 I4|_DFF_A|Q1  4.135667696e-12
LI4|_DFF_A|6 I4|_DFF_A|Q1 I4|A1_SYNC  2.067833848e-12
LI4|_DFF_B|1 I4|B1 I4|_DFF_B|A1  2.067833848e-12
LI4|_DFF_B|2 I4|_DFF_B|A1 I4|_DFF_B|A2  4.135667696e-12
LI4|_DFF_B|3 I4|_DFF_B|A3 I4|_DFF_B|A4  8.271335392e-12
LI4|_DFF_B|T T04 I4|_DFF_B|T1  2.067833848e-12
LI4|_DFF_B|4 I4|_DFF_B|T1 I4|_DFF_B|T2  4.135667696e-12
LI4|_DFF_B|5 I4|_DFF_B|A4 I4|_DFF_B|Q1  4.135667696e-12
LI4|_DFF_B|6 I4|_DFF_B|Q1 I4|B1_SYNC  2.067833848e-12
LI4|_XOR|A1 I4|A2 I4|_XOR|A1  2.067833848e-12
LI4|_XOR|A2 I4|_XOR|A1 I4|_XOR|A2  4.135667696e-12
LI4|_XOR|A3 I4|_XOR|A3 I4|_XOR|AB  8.271335392e-12
LI4|_XOR|B1 I4|B2 I4|_XOR|B1  2.067833848e-12
LI4|_XOR|B2 I4|_XOR|B1 I4|_XOR|B2  4.135667696e-12
LI4|_XOR|B3 I4|_XOR|B3 I4|_XOR|AB  8.271335392e-12
LI4|_XOR|T1 T04 I4|_XOR|T1  2.067833848e-12
LI4|_XOR|T2 I4|_XOR|T1 I4|_XOR|T2  4.135667696e-12
LI4|_XOR|Q2 I4|_XOR|ABTQ I4|_XOR|Q1  4.135667696e-12
LI4|_XOR|Q1 I4|_XOR|Q1 IP4_0  2.067833848e-12
LI4|_AND|A1 I4|A1_SYNC I4|_AND|A1  2.067833848e-12
LI4|_AND|A2 I4|_AND|A1 I4|_AND|A2  4.135667696e-12
LI4|_AND|A3 I4|_AND|A3 I4|_AND|Q3  1.2e-12
LI4|_AND|B1 I4|B1_SYNC I4|_AND|B1  2.067833848e-12
LI4|_AND|B2 I4|_AND|B1 I4|_AND|B2  4.135667696e-12
LI4|_AND|B3 I4|_AND|B3 I4|_AND|Q3  1.2e-12
LI4|_AND|Q3 I4|_AND|Q3 I4|_AND|Q2  4.135667696e-12
LI4|_AND|Q2 I4|_AND|Q2 I4|_AND|Q1  4.135667696e-12
LI4|_AND|Q1 I4|_AND|Q1 IG4_0  2.067833848e-12
LI5|_SPL_A|1 A5_RX I5|_SPL_A|D1  2e-12
LI5|_SPL_A|2 I5|_SPL_A|D1 I5|_SPL_A|D2  4.135667696e-12
LI5|_SPL_A|3 I5|_SPL_A|D2 I5|_SPL_A|JCT  9.84682784761905e-13
LI5|_SPL_A|4 I5|_SPL_A|JCT I5|_SPL_A|QA1  9.84682784761905e-13
LI5|_SPL_A|5 I5|_SPL_A|QA1 I5|A1  2e-12
LI5|_SPL_A|6 I5|_SPL_A|JCT I5|_SPL_A|QB1  9.84682784761905e-13
LI5|_SPL_A|7 I5|_SPL_A|QB1 I5|A2  2e-12
LI5|_SPL_B|1 B5_RX I5|_SPL_B|D1  2e-12
LI5|_SPL_B|2 I5|_SPL_B|D1 I5|_SPL_B|D2  4.135667696e-12
LI5|_SPL_B|3 I5|_SPL_B|D2 I5|_SPL_B|JCT  9.84682784761905e-13
LI5|_SPL_B|4 I5|_SPL_B|JCT I5|_SPL_B|QA1  9.84682784761905e-13
LI5|_SPL_B|5 I5|_SPL_B|QA1 I5|B1  2e-12
LI5|_SPL_B|6 I5|_SPL_B|JCT I5|_SPL_B|QB1  9.84682784761905e-13
LI5|_SPL_B|7 I5|_SPL_B|QB1 I5|B2  2e-12
LI5|_DFF_A|1 I5|A1 I5|_DFF_A|A1  2.067833848e-12
LI5|_DFF_A|2 I5|_DFF_A|A1 I5|_DFF_A|A2  4.135667696e-12
LI5|_DFF_A|3 I5|_DFF_A|A3 I5|_DFF_A|A4  8.271335392e-12
LI5|_DFF_A|T T05 I5|_DFF_A|T1  2.067833848e-12
LI5|_DFF_A|4 I5|_DFF_A|T1 I5|_DFF_A|T2  4.135667696e-12
LI5|_DFF_A|5 I5|_DFF_A|A4 I5|_DFF_A|Q1  4.135667696e-12
LI5|_DFF_A|6 I5|_DFF_A|Q1 I5|A1_SYNC  2.067833848e-12
LI5|_DFF_B|1 I5|B1 I5|_DFF_B|A1  2.067833848e-12
LI5|_DFF_B|2 I5|_DFF_B|A1 I5|_DFF_B|A2  4.135667696e-12
LI5|_DFF_B|3 I5|_DFF_B|A3 I5|_DFF_B|A4  8.271335392e-12
LI5|_DFF_B|T T05 I5|_DFF_B|T1  2.067833848e-12
LI5|_DFF_B|4 I5|_DFF_B|T1 I5|_DFF_B|T2  4.135667696e-12
LI5|_DFF_B|5 I5|_DFF_B|A4 I5|_DFF_B|Q1  4.135667696e-12
LI5|_DFF_B|6 I5|_DFF_B|Q1 I5|B1_SYNC  2.067833848e-12
LI5|_XOR|A1 I5|A2 I5|_XOR|A1  2.067833848e-12
LI5|_XOR|A2 I5|_XOR|A1 I5|_XOR|A2  4.135667696e-12
LI5|_XOR|A3 I5|_XOR|A3 I5|_XOR|AB  8.271335392e-12
LI5|_XOR|B1 I5|B2 I5|_XOR|B1  2.067833848e-12
LI5|_XOR|B2 I5|_XOR|B1 I5|_XOR|B2  4.135667696e-12
LI5|_XOR|B3 I5|_XOR|B3 I5|_XOR|AB  8.271335392e-12
LI5|_XOR|T1 T05 I5|_XOR|T1  2.067833848e-12
LI5|_XOR|T2 I5|_XOR|T1 I5|_XOR|T2  4.135667696e-12
LI5|_XOR|Q2 I5|_XOR|ABTQ I5|_XOR|Q1  4.135667696e-12
LI5|_XOR|Q1 I5|_XOR|Q1 IP5_0  2.067833848e-12
LI5|_AND|A1 I5|A1_SYNC I5|_AND|A1  2.067833848e-12
LI5|_AND|A2 I5|_AND|A1 I5|_AND|A2  4.135667696e-12
LI5|_AND|A3 I5|_AND|A3 I5|_AND|Q3  1.2e-12
LI5|_AND|B1 I5|B1_SYNC I5|_AND|B1  2.067833848e-12
LI5|_AND|B2 I5|_AND|B1 I5|_AND|B2  4.135667696e-12
LI5|_AND|B3 I5|_AND|B3 I5|_AND|Q3  1.2e-12
LI5|_AND|Q3 I5|_AND|Q3 I5|_AND|Q2  4.135667696e-12
LI5|_AND|Q2 I5|_AND|Q2 I5|_AND|Q1  4.135667696e-12
LI5|_AND|Q1 I5|_AND|Q1 IG5_0  2.067833848e-12
LI6|_SPL_A|1 A6_RX I6|_SPL_A|D1  2e-12
LI6|_SPL_A|2 I6|_SPL_A|D1 I6|_SPL_A|D2  4.135667696e-12
LI6|_SPL_A|3 I6|_SPL_A|D2 I6|_SPL_A|JCT  9.84682784761905e-13
LI6|_SPL_A|4 I6|_SPL_A|JCT I6|_SPL_A|QA1  9.84682784761905e-13
LI6|_SPL_A|5 I6|_SPL_A|QA1 I6|A1  2e-12
LI6|_SPL_A|6 I6|_SPL_A|JCT I6|_SPL_A|QB1  9.84682784761905e-13
LI6|_SPL_A|7 I6|_SPL_A|QB1 I6|A2  2e-12
LI6|_SPL_B|1 B6_RX I6|_SPL_B|D1  2e-12
LI6|_SPL_B|2 I6|_SPL_B|D1 I6|_SPL_B|D2  4.135667696e-12
LI6|_SPL_B|3 I6|_SPL_B|D2 I6|_SPL_B|JCT  9.84682784761905e-13
LI6|_SPL_B|4 I6|_SPL_B|JCT I6|_SPL_B|QA1  9.84682784761905e-13
LI6|_SPL_B|5 I6|_SPL_B|QA1 I6|B1  2e-12
LI6|_SPL_B|6 I6|_SPL_B|JCT I6|_SPL_B|QB1  9.84682784761905e-13
LI6|_SPL_B|7 I6|_SPL_B|QB1 I6|B2  2e-12
LI6|_DFF_A|1 I6|A1 I6|_DFF_A|A1  2.067833848e-12
LI6|_DFF_A|2 I6|_DFF_A|A1 I6|_DFF_A|A2  4.135667696e-12
LI6|_DFF_A|3 I6|_DFF_A|A3 I6|_DFF_A|A4  8.271335392e-12
LI6|_DFF_A|T T06 I6|_DFF_A|T1  2.067833848e-12
LI6|_DFF_A|4 I6|_DFF_A|T1 I6|_DFF_A|T2  4.135667696e-12
LI6|_DFF_A|5 I6|_DFF_A|A4 I6|_DFF_A|Q1  4.135667696e-12
LI6|_DFF_A|6 I6|_DFF_A|Q1 I6|A1_SYNC  2.067833848e-12
LI6|_DFF_B|1 I6|B1 I6|_DFF_B|A1  2.067833848e-12
LI6|_DFF_B|2 I6|_DFF_B|A1 I6|_DFF_B|A2  4.135667696e-12
LI6|_DFF_B|3 I6|_DFF_B|A3 I6|_DFF_B|A4  8.271335392e-12
LI6|_DFF_B|T T06 I6|_DFF_B|T1  2.067833848e-12
LI6|_DFF_B|4 I6|_DFF_B|T1 I6|_DFF_B|T2  4.135667696e-12
LI6|_DFF_B|5 I6|_DFF_B|A4 I6|_DFF_B|Q1  4.135667696e-12
LI6|_DFF_B|6 I6|_DFF_B|Q1 I6|B1_SYNC  2.067833848e-12
LI6|_XOR|A1 I6|A2 I6|_XOR|A1  2.067833848e-12
LI6|_XOR|A2 I6|_XOR|A1 I6|_XOR|A2  4.135667696e-12
LI6|_XOR|A3 I6|_XOR|A3 I6|_XOR|AB  8.271335392e-12
LI6|_XOR|B1 I6|B2 I6|_XOR|B1  2.067833848e-12
LI6|_XOR|B2 I6|_XOR|B1 I6|_XOR|B2  4.135667696e-12
LI6|_XOR|B3 I6|_XOR|B3 I6|_XOR|AB  8.271335392e-12
LI6|_XOR|T1 T06 I6|_XOR|T1  2.067833848e-12
LI6|_XOR|T2 I6|_XOR|T1 I6|_XOR|T2  4.135667696e-12
LI6|_XOR|Q2 I6|_XOR|ABTQ I6|_XOR|Q1  4.135667696e-12
LI6|_XOR|Q1 I6|_XOR|Q1 IP6_0  2.067833848e-12
LI6|_AND|A1 I6|A1_SYNC I6|_AND|A1  2.067833848e-12
LI6|_AND|A2 I6|_AND|A1 I6|_AND|A2  4.135667696e-12
LI6|_AND|A3 I6|_AND|A3 I6|_AND|Q3  1.2e-12
LI6|_AND|B1 I6|B1_SYNC I6|_AND|B1  2.067833848e-12
LI6|_AND|B2 I6|_AND|B1 I6|_AND|B2  4.135667696e-12
LI6|_AND|B3 I6|_AND|B3 I6|_AND|Q3  1.2e-12
LI6|_AND|Q3 I6|_AND|Q3 I6|_AND|Q2  4.135667696e-12
LI6|_AND|Q2 I6|_AND|Q2 I6|_AND|Q1  4.135667696e-12
LI6|_AND|Q1 I6|_AND|Q1 IG6_0  2.067833848e-12
LI7|_SPL_A|1 A7_RX I7|_SPL_A|D1  2e-12
LI7|_SPL_A|2 I7|_SPL_A|D1 I7|_SPL_A|D2  4.135667696e-12
LI7|_SPL_A|3 I7|_SPL_A|D2 I7|_SPL_A|JCT  9.84682784761905e-13
LI7|_SPL_A|4 I7|_SPL_A|JCT I7|_SPL_A|QA1  9.84682784761905e-13
LI7|_SPL_A|5 I7|_SPL_A|QA1 I7|A1  2e-12
LI7|_SPL_A|6 I7|_SPL_A|JCT I7|_SPL_A|QB1  9.84682784761905e-13
LI7|_SPL_A|7 I7|_SPL_A|QB1 I7|A2  2e-12
LI7|_SPL_B|1 B7_RX I7|_SPL_B|D1  2e-12
LI7|_SPL_B|2 I7|_SPL_B|D1 I7|_SPL_B|D2  4.135667696e-12
LI7|_SPL_B|3 I7|_SPL_B|D2 I7|_SPL_B|JCT  9.84682784761905e-13
LI7|_SPL_B|4 I7|_SPL_B|JCT I7|_SPL_B|QA1  9.84682784761905e-13
LI7|_SPL_B|5 I7|_SPL_B|QA1 I7|B1  2e-12
LI7|_SPL_B|6 I7|_SPL_B|JCT I7|_SPL_B|QB1  9.84682784761905e-13
LI7|_SPL_B|7 I7|_SPL_B|QB1 I7|B2  2e-12
LI7|_DFF_A|1 I7|A1 I7|_DFF_A|A1  2.067833848e-12
LI7|_DFF_A|2 I7|_DFF_A|A1 I7|_DFF_A|A2  4.135667696e-12
LI7|_DFF_A|3 I7|_DFF_A|A3 I7|_DFF_A|A4  8.271335392e-12
LI7|_DFF_A|T T07 I7|_DFF_A|T1  2.067833848e-12
LI7|_DFF_A|4 I7|_DFF_A|T1 I7|_DFF_A|T2  4.135667696e-12
LI7|_DFF_A|5 I7|_DFF_A|A4 I7|_DFF_A|Q1  4.135667696e-12
LI7|_DFF_A|6 I7|_DFF_A|Q1 I7|A1_SYNC  2.067833848e-12
LI7|_DFF_B|1 I7|B1 I7|_DFF_B|A1  2.067833848e-12
LI7|_DFF_B|2 I7|_DFF_B|A1 I7|_DFF_B|A2  4.135667696e-12
LI7|_DFF_B|3 I7|_DFF_B|A3 I7|_DFF_B|A4  8.271335392e-12
LI7|_DFF_B|T T07 I7|_DFF_B|T1  2.067833848e-12
LI7|_DFF_B|4 I7|_DFF_B|T1 I7|_DFF_B|T2  4.135667696e-12
LI7|_DFF_B|5 I7|_DFF_B|A4 I7|_DFF_B|Q1  4.135667696e-12
LI7|_DFF_B|6 I7|_DFF_B|Q1 I7|B1_SYNC  2.067833848e-12
LI7|_XOR|A1 I7|A2 I7|_XOR|A1  2.067833848e-12
LI7|_XOR|A2 I7|_XOR|A1 I7|_XOR|A2  4.135667696e-12
LI7|_XOR|A3 I7|_XOR|A3 I7|_XOR|AB  8.271335392e-12
LI7|_XOR|B1 I7|B2 I7|_XOR|B1  2.067833848e-12
LI7|_XOR|B2 I7|_XOR|B1 I7|_XOR|B2  4.135667696e-12
LI7|_XOR|B3 I7|_XOR|B3 I7|_XOR|AB  8.271335392e-12
LI7|_XOR|T1 T07 I7|_XOR|T1  2.067833848e-12
LI7|_XOR|T2 I7|_XOR|T1 I7|_XOR|T2  4.135667696e-12
LI7|_XOR|Q2 I7|_XOR|ABTQ I7|_XOR|Q1  4.135667696e-12
LI7|_XOR|Q1 I7|_XOR|Q1 IP7_0  2.067833848e-12
LI7|_AND|A1 I7|A1_SYNC I7|_AND|A1  2.067833848e-12
LI7|_AND|A2 I7|_AND|A1 I7|_AND|A2  4.135667696e-12
LI7|_AND|A3 I7|_AND|A3 I7|_AND|Q3  1.2e-12
LI7|_AND|B1 I7|B1_SYNC I7|_AND|B1  2.067833848e-12
LI7|_AND|B2 I7|_AND|B1 I7|_AND|B2  4.135667696e-12
LI7|_AND|B3 I7|_AND|B3 I7|_AND|Q3  1.2e-12
LI7|_AND|Q3 I7|_AND|Q3 I7|_AND|Q2  4.135667696e-12
LI7|_AND|Q2 I7|_AND|Q2 I7|_AND|Q1  4.135667696e-12
LI7|_AND|Q1 I7|_AND|Q1 IG7_0  2.067833848e-12
B_PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP0_0|_TX|B1 0 _PTL_IP0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP0_0|_TX|B2 0 _PTL_IP0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|3  1.684e-12
L_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|6  3.596e-12
L_PTL_IP0_0|_TX|1 IP0_0 _PTL_IP0_0|_TX|1  2.063e-12
L_PTL_IP0_0|_TX|2 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|4  4.123e-12
L_PTL_IP0_0|_TX|3 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|7  2.193e-12
R_PTL_IP0_0|_TX|D _PTL_IP0_0|_TX|7 _PTL_IP0_0|A_PTL  1.36
L_PTL_IP0_0|_TX|P1 _PTL_IP0_0|_TX|2 0  5.254e-13
L_PTL_IP0_0|_TX|P2 _PTL_IP0_0|_TX|5 0  5.141e-13
R_PTL_IP0_0|_TX|B1 _PTL_IP0_0|_TX|1 _PTL_IP0_0|_TX|101  2.7439617672
R_PTL_IP0_0|_TX|B2 _PTL_IP0_0|_TX|4 _PTL_IP0_0|_TX|104  2.7439617672
L_PTL_IP0_0|_TX|RB1 _PTL_IP0_0|_TX|101 0  1.550338398468e-12
L_PTL_IP0_0|_TX|RB2 _PTL_IP0_0|_TX|104 0  1.550338398468e-12
B_PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP0_0|_RX|B1 0 _PTL_IP0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|3  2.777e-12
I_PTL_IP0_0|_RX|B2 0 _PTL_IP0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|6  2.685e-12
I_PTL_IP0_0|_RX|B3 0 _PTL_IP0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|9  2.764e-12
L_PTL_IP0_0|_RX|1 _PTL_IP0_0|A_PTL _PTL_IP0_0|_RX|1  1.346e-12
L_PTL_IP0_0|_RX|2 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|4  6.348e-12
L_PTL_IP0_0|_RX|3 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7  5.197e-12
L_PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|7 _PTL_IP0_0|D  2.058e-12
L_PTL_IP0_0|_RX|P1 _PTL_IP0_0|_RX|2 0  4.795e-13
L_PTL_IP0_0|_RX|P2 _PTL_IP0_0|_RX|5 0  5.431e-13
L_PTL_IP0_0|_RX|P3 _PTL_IP0_0|_RX|8 0  5.339e-13
R_PTL_IP0_0|_RX|B1 _PTL_IP0_0|_RX|1 _PTL_IP0_0|_RX|101  4.225701121488
R_PTL_IP0_0|_RX|B2 _PTL_IP0_0|_RX|4 _PTL_IP0_0|_RX|104  3.429952209
R_PTL_IP0_0|_RX|B3 _PTL_IP0_0|_RX|7 _PTL_IP0_0|_RX|107  2.7439617672
L_PTL_IP0_0|_RX|RB1 _PTL_IP0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP0_0|_RX|RB2 _PTL_IP0_0|_RX|104 0  1.937922998085e-12
L_PTL_IP0_0|_RX|RB3 _PTL_IP0_0|_RX|107 0  1.550338398468e-12
L_PTL_IP0_0|_SPL|1 _PTL_IP0_0|D _PTL_IP0_0|_SPL|D1  2e-12
L_PTL_IP0_0|_SPL|2 _PTL_IP0_0|_SPL|D1 _PTL_IP0_0|_SPL|D2  4.135667696e-12
L_PTL_IP0_0|_SPL|3 _PTL_IP0_0|_SPL|D2 _PTL_IP0_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP0_0|_SPL|4 _PTL_IP0_0|_SPL|JCT _PTL_IP0_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP0_0|_SPL|5 _PTL_IP0_0|_SPL|QA1 IP0_0_TO1  2e-12
L_PTL_IP0_0|_SPL|6 _PTL_IP0_0|_SPL|JCT _PTL_IP0_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP0_0|_SPL|7 _PTL_IP0_0|_SPL|QB1 S0_0  2e-12
B_PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG0_0|_TX|B1 0 _PTL_IG0_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG0_0|_TX|B2 0 _PTL_IG0_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|3  1.684e-12
L_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|6  3.596e-12
L_PTL_IG0_0|_TX|1 IG0_0 _PTL_IG0_0|_TX|1  2.063e-12
L_PTL_IG0_0|_TX|2 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|4  4.123e-12
L_PTL_IG0_0|_TX|3 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|7  2.193e-12
R_PTL_IG0_0|_TX|D _PTL_IG0_0|_TX|7 _PTL_IG0_0|A_PTL  1.36
L_PTL_IG0_0|_TX|P1 _PTL_IG0_0|_TX|2 0  5.254e-13
L_PTL_IG0_0|_TX|P2 _PTL_IG0_0|_TX|5 0  5.141e-13
R_PTL_IG0_0|_TX|B1 _PTL_IG0_0|_TX|1 _PTL_IG0_0|_TX|101  2.7439617672
R_PTL_IG0_0|_TX|B2 _PTL_IG0_0|_TX|4 _PTL_IG0_0|_TX|104  2.7439617672
L_PTL_IG0_0|_TX|RB1 _PTL_IG0_0|_TX|101 0  1.550338398468e-12
L_PTL_IG0_0|_TX|RB2 _PTL_IG0_0|_TX|104 0  1.550338398468e-12
B_PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG0_0|_RX|B1 0 _PTL_IG0_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|3  2.777e-12
I_PTL_IG0_0|_RX|B2 0 _PTL_IG0_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|6  2.685e-12
I_PTL_IG0_0|_RX|B3 0 _PTL_IG0_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|9  2.764e-12
L_PTL_IG0_0|_RX|1 _PTL_IG0_0|A_PTL _PTL_IG0_0|_RX|1  1.346e-12
L_PTL_IG0_0|_RX|2 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|4  6.348e-12
L_PTL_IG0_0|_RX|3 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7  5.197e-12
L_PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|7 _PTL_IG0_0|D  2.058e-12
L_PTL_IG0_0|_RX|P1 _PTL_IG0_0|_RX|2 0  4.795e-13
L_PTL_IG0_0|_RX|P2 _PTL_IG0_0|_RX|5 0  5.431e-13
L_PTL_IG0_0|_RX|P3 _PTL_IG0_0|_RX|8 0  5.339e-13
R_PTL_IG0_0|_RX|B1 _PTL_IG0_0|_RX|1 _PTL_IG0_0|_RX|101  4.225701121488
R_PTL_IG0_0|_RX|B2 _PTL_IG0_0|_RX|4 _PTL_IG0_0|_RX|104  3.429952209
R_PTL_IG0_0|_RX|B3 _PTL_IG0_0|_RX|7 _PTL_IG0_0|_RX|107  2.7439617672
L_PTL_IG0_0|_RX|RB1 _PTL_IG0_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG0_0|_RX|RB2 _PTL_IG0_0|_RX|104 0  1.937922998085e-12
L_PTL_IG0_0|_RX|RB3 _PTL_IG0_0|_RX|107 0  1.550338398468e-12
L_PTL_IG0_0|_SPL|1 _PTL_IG0_0|D _PTL_IG0_0|_SPL|D1  2e-12
L_PTL_IG0_0|_SPL|2 _PTL_IG0_0|_SPL|D1 _PTL_IG0_0|_SPL|D2  4.135667696e-12
L_PTL_IG0_0|_SPL|3 _PTL_IG0_0|_SPL|D2 _PTL_IG0_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IG0_0|_SPL|4 _PTL_IG0_0|_SPL|JCT _PTL_IG0_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IG0_0|_SPL|5 _PTL_IG0_0|_SPL|QA1 IG0_0_TO0  2e-12
L_PTL_IG0_0|_SPL|6 _PTL_IG0_0|_SPL|JCT _PTL_IG0_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IG0_0|_SPL|7 _PTL_IG0_0|_SPL|QB1 IG0_0_TO1  2e-12
B_PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP1_0|_TX|B1 0 _PTL_IP1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP1_0|_TX|B2 0 _PTL_IP1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|3  1.684e-12
L_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|6  3.596e-12
L_PTL_IP1_0|_TX|1 IP1_0 _PTL_IP1_0|_TX|1  2.063e-12
L_PTL_IP1_0|_TX|2 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|4  4.123e-12
L_PTL_IP1_0|_TX|3 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|7  2.193e-12
R_PTL_IP1_0|_TX|D _PTL_IP1_0|_TX|7 _PTL_IP1_0|A_PTL  1.36
L_PTL_IP1_0|_TX|P1 _PTL_IP1_0|_TX|2 0  5.254e-13
L_PTL_IP1_0|_TX|P2 _PTL_IP1_0|_TX|5 0  5.141e-13
R_PTL_IP1_0|_TX|B1 _PTL_IP1_0|_TX|1 _PTL_IP1_0|_TX|101  2.7439617672
R_PTL_IP1_0|_TX|B2 _PTL_IP1_0|_TX|4 _PTL_IP1_0|_TX|104  2.7439617672
L_PTL_IP1_0|_TX|RB1 _PTL_IP1_0|_TX|101 0  1.550338398468e-12
L_PTL_IP1_0|_TX|RB2 _PTL_IP1_0|_TX|104 0  1.550338398468e-12
B_PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP1_0|_RX|B1 0 _PTL_IP1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|3  2.777e-12
I_PTL_IP1_0|_RX|B2 0 _PTL_IP1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|6  2.685e-12
I_PTL_IP1_0|_RX|B3 0 _PTL_IP1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|9  2.764e-12
L_PTL_IP1_0|_RX|1 _PTL_IP1_0|A_PTL _PTL_IP1_0|_RX|1  1.346e-12
L_PTL_IP1_0|_RX|2 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|4  6.348e-12
L_PTL_IP1_0|_RX|3 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7  5.197e-12
L_PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|7 _PTL_IP1_0|D  2.058e-12
L_PTL_IP1_0|_RX|P1 _PTL_IP1_0|_RX|2 0  4.795e-13
L_PTL_IP1_0|_RX|P2 _PTL_IP1_0|_RX|5 0  5.431e-13
L_PTL_IP1_0|_RX|P3 _PTL_IP1_0|_RX|8 0  5.339e-13
R_PTL_IP1_0|_RX|B1 _PTL_IP1_0|_RX|1 _PTL_IP1_0|_RX|101  4.225701121488
R_PTL_IP1_0|_RX|B2 _PTL_IP1_0|_RX|4 _PTL_IP1_0|_RX|104  3.429952209
R_PTL_IP1_0|_RX|B3 _PTL_IP1_0|_RX|7 _PTL_IP1_0|_RX|107  2.7439617672
L_PTL_IP1_0|_RX|RB1 _PTL_IP1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP1_0|_RX|RB2 _PTL_IP1_0|_RX|104 0  1.937922998085e-12
L_PTL_IP1_0|_RX|RB3 _PTL_IP1_0|_RX|107 0  1.550338398468e-12
L_PTL_IP1_0|_SPL|1 _PTL_IP1_0|D _PTL_IP1_0|_SPL|D1  2e-12
L_PTL_IP1_0|_SPL|2 _PTL_IP1_0|_SPL|D1 _PTL_IP1_0|_SPL|D2  4.135667696e-12
L_PTL_IP1_0|_SPL|3 _PTL_IP1_0|_SPL|D2 _PTL_IP1_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP1_0|_SPL|4 _PTL_IP1_0|_SPL|JCT _PTL_IP1_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP1_0|_SPL|5 _PTL_IP1_0|_SPL|QA1 IP1_0_TO1  2e-12
L_PTL_IP1_0|_SPL|6 _PTL_IP1_0|_SPL|JCT _PTL_IP1_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP1_0|_SPL|7 _PTL_IP1_0|_SPL|QB1 IP1_0_OUT  2e-12
B_PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG1_0|_TX|B1 0 _PTL_IG1_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG1_0|_TX|B2 0 _PTL_IG1_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|3  1.684e-12
L_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|6  3.596e-12
L_PTL_IG1_0|_TX|1 IG1_0 _PTL_IG1_0|_TX|1  2.063e-12
L_PTL_IG1_0|_TX|2 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|4  4.123e-12
L_PTL_IG1_0|_TX|3 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|7  2.193e-12
R_PTL_IG1_0|_TX|D _PTL_IG1_0|_TX|7 _PTL_IG1_0|A_PTL  1.36
L_PTL_IG1_0|_TX|P1 _PTL_IG1_0|_TX|2 0  5.254e-13
L_PTL_IG1_0|_TX|P2 _PTL_IG1_0|_TX|5 0  5.141e-13
R_PTL_IG1_0|_TX|B1 _PTL_IG1_0|_TX|1 _PTL_IG1_0|_TX|101  2.7439617672
R_PTL_IG1_0|_TX|B2 _PTL_IG1_0|_TX|4 _PTL_IG1_0|_TX|104  2.7439617672
L_PTL_IG1_0|_TX|RB1 _PTL_IG1_0|_TX|101 0  1.550338398468e-12
L_PTL_IG1_0|_TX|RB2 _PTL_IG1_0|_TX|104 0  1.550338398468e-12
B_PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG1_0|_RX|B1 0 _PTL_IG1_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|3  2.777e-12
I_PTL_IG1_0|_RX|B2 0 _PTL_IG1_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|6  2.685e-12
I_PTL_IG1_0|_RX|B3 0 _PTL_IG1_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|9  2.764e-12
L_PTL_IG1_0|_RX|1 _PTL_IG1_0|A_PTL _PTL_IG1_0|_RX|1  1.346e-12
L_PTL_IG1_0|_RX|2 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|4  6.348e-12
L_PTL_IG1_0|_RX|3 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7  5.197e-12
L_PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|7 IG1_0_TO1  2.058e-12
L_PTL_IG1_0|_RX|P1 _PTL_IG1_0|_RX|2 0  4.795e-13
L_PTL_IG1_0|_RX|P2 _PTL_IG1_0|_RX|5 0  5.431e-13
L_PTL_IG1_0|_RX|P3 _PTL_IG1_0|_RX|8 0  5.339e-13
R_PTL_IG1_0|_RX|B1 _PTL_IG1_0|_RX|1 _PTL_IG1_0|_RX|101  4.225701121488
R_PTL_IG1_0|_RX|B2 _PTL_IG1_0|_RX|4 _PTL_IG1_0|_RX|104  3.429952209
R_PTL_IG1_0|_RX|B3 _PTL_IG1_0|_RX|7 _PTL_IG1_0|_RX|107  2.7439617672
L_PTL_IG1_0|_RX|RB1 _PTL_IG1_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG1_0|_RX|RB2 _PTL_IG1_0|_RX|104 0  1.937922998085e-12
L_PTL_IG1_0|_RX|RB3 _PTL_IG1_0|_RX|107 0  1.550338398468e-12
B_PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP2_0|_TX|B1 0 _PTL_IP2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP2_0|_TX|B2 0 _PTL_IP2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|3  1.684e-12
L_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|6  3.596e-12
L_PTL_IP2_0|_TX|1 IP2_0 _PTL_IP2_0|_TX|1  2.063e-12
L_PTL_IP2_0|_TX|2 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|4  4.123e-12
L_PTL_IP2_0|_TX|3 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|7  2.193e-12
R_PTL_IP2_0|_TX|D _PTL_IP2_0|_TX|7 _PTL_IP2_0|A_PTL  1.36
L_PTL_IP2_0|_TX|P1 _PTL_IP2_0|_TX|2 0  5.254e-13
L_PTL_IP2_0|_TX|P2 _PTL_IP2_0|_TX|5 0  5.141e-13
R_PTL_IP2_0|_TX|B1 _PTL_IP2_0|_TX|1 _PTL_IP2_0|_TX|101  2.7439617672
R_PTL_IP2_0|_TX|B2 _PTL_IP2_0|_TX|4 _PTL_IP2_0|_TX|104  2.7439617672
L_PTL_IP2_0|_TX|RB1 _PTL_IP2_0|_TX|101 0  1.550338398468e-12
L_PTL_IP2_0|_TX|RB2 _PTL_IP2_0|_TX|104 0  1.550338398468e-12
B_PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP2_0|_RX|B1 0 _PTL_IP2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|3  2.777e-12
I_PTL_IP2_0|_RX|B2 0 _PTL_IP2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|6  2.685e-12
I_PTL_IP2_0|_RX|B3 0 _PTL_IP2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|9  2.764e-12
L_PTL_IP2_0|_RX|1 _PTL_IP2_0|A_PTL _PTL_IP2_0|_RX|1  1.346e-12
L_PTL_IP2_0|_RX|2 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|4  6.348e-12
L_PTL_IP2_0|_RX|3 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7  5.197e-12
L_PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|7 _PTL_IP2_0|D  2.058e-12
L_PTL_IP2_0|_RX|P1 _PTL_IP2_0|_RX|2 0  4.795e-13
L_PTL_IP2_0|_RX|P2 _PTL_IP2_0|_RX|5 0  5.431e-13
L_PTL_IP2_0|_RX|P3 _PTL_IP2_0|_RX|8 0  5.339e-13
R_PTL_IP2_0|_RX|B1 _PTL_IP2_0|_RX|1 _PTL_IP2_0|_RX|101  4.225701121488
R_PTL_IP2_0|_RX|B2 _PTL_IP2_0|_RX|4 _PTL_IP2_0|_RX|104  3.429952209
R_PTL_IP2_0|_RX|B3 _PTL_IP2_0|_RX|7 _PTL_IP2_0|_RX|107  2.7439617672
L_PTL_IP2_0|_RX|RB1 _PTL_IP2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP2_0|_RX|RB2 _PTL_IP2_0|_RX|104 0  1.937922998085e-12
L_PTL_IP2_0|_RX|RB3 _PTL_IP2_0|_RX|107 0  1.550338398468e-12
L_PTL_IP2_0|_SPL|1 _PTL_IP2_0|D _PTL_IP2_0|_SPL|D1  2e-12
L_PTL_IP2_0|_SPL|2 _PTL_IP2_0|_SPL|D1 _PTL_IP2_0|_SPL|D2  4.135667696e-12
L_PTL_IP2_0|_SPL|3 _PTL_IP2_0|_SPL|D2 _PTL_IP2_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP2_0|_SPL|4 _PTL_IP2_0|_SPL|JCT _PTL_IP2_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP2_0|_SPL|5 _PTL_IP2_0|_SPL|QA1 IP2_0_TO2  2e-12
L_PTL_IP2_0|_SPL|6 _PTL_IP2_0|_SPL|JCT _PTL_IP2_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP2_0|_SPL|7 _PTL_IP2_0|_SPL|QB1 IP2_0_TO3  2e-12
B_PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG2_0|_TX|B1 0 _PTL_IG2_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG2_0|_TX|B2 0 _PTL_IG2_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|3  1.684e-12
L_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|6  3.596e-12
L_PTL_IG2_0|_TX|1 IG2_0 _PTL_IG2_0|_TX|1  2.063e-12
L_PTL_IG2_0|_TX|2 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|4  4.123e-12
L_PTL_IG2_0|_TX|3 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|7  2.193e-12
R_PTL_IG2_0|_TX|D _PTL_IG2_0|_TX|7 _PTL_IG2_0|A_PTL  1.36
L_PTL_IG2_0|_TX|P1 _PTL_IG2_0|_TX|2 0  5.254e-13
L_PTL_IG2_0|_TX|P2 _PTL_IG2_0|_TX|5 0  5.141e-13
R_PTL_IG2_0|_TX|B1 _PTL_IG2_0|_TX|1 _PTL_IG2_0|_TX|101  2.7439617672
R_PTL_IG2_0|_TX|B2 _PTL_IG2_0|_TX|4 _PTL_IG2_0|_TX|104  2.7439617672
L_PTL_IG2_0|_TX|RB1 _PTL_IG2_0|_TX|101 0  1.550338398468e-12
L_PTL_IG2_0|_TX|RB2 _PTL_IG2_0|_TX|104 0  1.550338398468e-12
B_PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG2_0|_RX|B1 0 _PTL_IG2_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|3  2.777e-12
I_PTL_IG2_0|_RX|B2 0 _PTL_IG2_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|6  2.685e-12
I_PTL_IG2_0|_RX|B3 0 _PTL_IG2_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|9  2.764e-12
L_PTL_IG2_0|_RX|1 _PTL_IG2_0|A_PTL _PTL_IG2_0|_RX|1  1.346e-12
L_PTL_IG2_0|_RX|2 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|4  6.348e-12
L_PTL_IG2_0|_RX|3 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7  5.197e-12
L_PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|7 _PTL_IG2_0|D  2.058e-12
L_PTL_IG2_0|_RX|P1 _PTL_IG2_0|_RX|2 0  4.795e-13
L_PTL_IG2_0|_RX|P2 _PTL_IG2_0|_RX|5 0  5.431e-13
L_PTL_IG2_0|_RX|P3 _PTL_IG2_0|_RX|8 0  5.339e-13
R_PTL_IG2_0|_RX|B1 _PTL_IG2_0|_RX|1 _PTL_IG2_0|_RX|101  4.225701121488
R_PTL_IG2_0|_RX|B2 _PTL_IG2_0|_RX|4 _PTL_IG2_0|_RX|104  3.429952209
R_PTL_IG2_0|_RX|B3 _PTL_IG2_0|_RX|7 _PTL_IG2_0|_RX|107  2.7439617672
L_PTL_IG2_0|_RX|RB1 _PTL_IG2_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG2_0|_RX|RB2 _PTL_IG2_0|_RX|104 0  1.937922998085e-12
L_PTL_IG2_0|_RX|RB3 _PTL_IG2_0|_RX|107 0  1.550338398468e-12
L_PTL_IG2_0|_SPL|1 _PTL_IG2_0|D _PTL_IG2_0|_SPL|D1  2e-12
L_PTL_IG2_0|_SPL|2 _PTL_IG2_0|_SPL|D1 _PTL_IG2_0|_SPL|D2  4.135667696e-12
L_PTL_IG2_0|_SPL|3 _PTL_IG2_0|_SPL|D2 _PTL_IG2_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IG2_0|_SPL|4 _PTL_IG2_0|_SPL|JCT _PTL_IG2_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IG2_0|_SPL|5 _PTL_IG2_0|_SPL|QA1 IG2_0_TO2  2e-12
L_PTL_IG2_0|_SPL|6 _PTL_IG2_0|_SPL|JCT _PTL_IG2_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IG2_0|_SPL|7 _PTL_IG2_0|_SPL|QB1 IG2_0_TO3  2e-12
B_PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_0|_TX|B1 0 _PTL_IP3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_0|_TX|B2 0 _PTL_IP3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|3  1.684e-12
L_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|6  3.596e-12
L_PTL_IP3_0|_TX|1 IP3_0 _PTL_IP3_0|_TX|1  2.063e-12
L_PTL_IP3_0|_TX|2 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|4  4.123e-12
L_PTL_IP3_0|_TX|3 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|7  2.193e-12
R_PTL_IP3_0|_TX|D _PTL_IP3_0|_TX|7 _PTL_IP3_0|A_PTL  1.36
L_PTL_IP3_0|_TX|P1 _PTL_IP3_0|_TX|2 0  5.254e-13
L_PTL_IP3_0|_TX|P2 _PTL_IP3_0|_TX|5 0  5.141e-13
R_PTL_IP3_0|_TX|B1 _PTL_IP3_0|_TX|1 _PTL_IP3_0|_TX|101  2.7439617672
R_PTL_IP3_0|_TX|B2 _PTL_IP3_0|_TX|4 _PTL_IP3_0|_TX|104  2.7439617672
L_PTL_IP3_0|_TX|RB1 _PTL_IP3_0|_TX|101 0  1.550338398468e-12
L_PTL_IP3_0|_TX|RB2 _PTL_IP3_0|_TX|104 0  1.550338398468e-12
B_PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_0|_RX|B1 0 _PTL_IP3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|3  2.777e-12
I_PTL_IP3_0|_RX|B2 0 _PTL_IP3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|6  2.685e-12
I_PTL_IP3_0|_RX|B3 0 _PTL_IP3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|9  2.764e-12
L_PTL_IP3_0|_RX|1 _PTL_IP3_0|A_PTL _PTL_IP3_0|_RX|1  1.346e-12
L_PTL_IP3_0|_RX|2 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|4  6.348e-12
L_PTL_IP3_0|_RX|3 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7  5.197e-12
L_PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|7 _PTL_IP3_0|D  2.058e-12
L_PTL_IP3_0|_RX|P1 _PTL_IP3_0|_RX|2 0  4.795e-13
L_PTL_IP3_0|_RX|P2 _PTL_IP3_0|_RX|5 0  5.431e-13
L_PTL_IP3_0|_RX|P3 _PTL_IP3_0|_RX|8 0  5.339e-13
R_PTL_IP3_0|_RX|B1 _PTL_IP3_0|_RX|1 _PTL_IP3_0|_RX|101  4.225701121488
R_PTL_IP3_0|_RX|B2 _PTL_IP3_0|_RX|4 _PTL_IP3_0|_RX|104  3.429952209
R_PTL_IP3_0|_RX|B3 _PTL_IP3_0|_RX|7 _PTL_IP3_0|_RX|107  2.7439617672
L_PTL_IP3_0|_RX|RB1 _PTL_IP3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_0|_RX|RB2 _PTL_IP3_0|_RX|104 0  1.937922998085e-12
L_PTL_IP3_0|_RX|RB3 _PTL_IP3_0|_RX|107 0  1.550338398468e-12
L_PTL_IP3_0|_SPL|1 _PTL_IP3_0|D _PTL_IP3_0|_SPL|D1  2e-12
L_PTL_IP3_0|_SPL|2 _PTL_IP3_0|_SPL|D1 _PTL_IP3_0|_SPL|D2  4.135667696e-12
L_PTL_IP3_0|_SPL|3 _PTL_IP3_0|_SPL|D2 _PTL_IP3_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP3_0|_SPL|4 _PTL_IP3_0|_SPL|JCT _PTL_IP3_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP3_0|_SPL|5 _PTL_IP3_0|_SPL|QA1 IP3_0_TO3  2e-12
L_PTL_IP3_0|_SPL|6 _PTL_IP3_0|_SPL|JCT _PTL_IP3_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP3_0|_SPL|7 _PTL_IP3_0|_SPL|QB1 IP3_0_OUT  2e-12
B_PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG3_0|_TX|B1 0 _PTL_IG3_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG3_0|_TX|B2 0 _PTL_IG3_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|3  1.684e-12
L_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|6  3.596e-12
L_PTL_IG3_0|_TX|1 IG3_0 _PTL_IG3_0|_TX|1  2.063e-12
L_PTL_IG3_0|_TX|2 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|4  4.123e-12
L_PTL_IG3_0|_TX|3 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|7  2.193e-12
R_PTL_IG3_0|_TX|D _PTL_IG3_0|_TX|7 _PTL_IG3_0|A_PTL  1.36
L_PTL_IG3_0|_TX|P1 _PTL_IG3_0|_TX|2 0  5.254e-13
L_PTL_IG3_0|_TX|P2 _PTL_IG3_0|_TX|5 0  5.141e-13
R_PTL_IG3_0|_TX|B1 _PTL_IG3_0|_TX|1 _PTL_IG3_0|_TX|101  2.7439617672
R_PTL_IG3_0|_TX|B2 _PTL_IG3_0|_TX|4 _PTL_IG3_0|_TX|104  2.7439617672
L_PTL_IG3_0|_TX|RB1 _PTL_IG3_0|_TX|101 0  1.550338398468e-12
L_PTL_IG3_0|_TX|RB2 _PTL_IG3_0|_TX|104 0  1.550338398468e-12
B_PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG3_0|_RX|B1 0 _PTL_IG3_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|3  2.777e-12
I_PTL_IG3_0|_RX|B2 0 _PTL_IG3_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|6  2.685e-12
I_PTL_IG3_0|_RX|B3 0 _PTL_IG3_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|9  2.764e-12
L_PTL_IG3_0|_RX|1 _PTL_IG3_0|A_PTL _PTL_IG3_0|_RX|1  1.346e-12
L_PTL_IG3_0|_RX|2 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|4  6.348e-12
L_PTL_IG3_0|_RX|3 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7  5.197e-12
L_PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|7 IG3_0_TO3  2.058e-12
L_PTL_IG3_0|_RX|P1 _PTL_IG3_0|_RX|2 0  4.795e-13
L_PTL_IG3_0|_RX|P2 _PTL_IG3_0|_RX|5 0  5.431e-13
L_PTL_IG3_0|_RX|P3 _PTL_IG3_0|_RX|8 0  5.339e-13
R_PTL_IG3_0|_RX|B1 _PTL_IG3_0|_RX|1 _PTL_IG3_0|_RX|101  4.225701121488
R_PTL_IG3_0|_RX|B2 _PTL_IG3_0|_RX|4 _PTL_IG3_0|_RX|104  3.429952209
R_PTL_IG3_0|_RX|B3 _PTL_IG3_0|_RX|7 _PTL_IG3_0|_RX|107  2.7439617672
L_PTL_IG3_0|_RX|RB1 _PTL_IG3_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG3_0|_RX|RB2 _PTL_IG3_0|_RX|104 0  1.937922998085e-12
L_PTL_IG3_0|_RX|RB3 _PTL_IG3_0|_RX|107 0  1.550338398468e-12
B_PTL_IP4_0|_TX|1 _PTL_IP4_0|_TX|1 _PTL_IP4_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP4_0|_TX|2 _PTL_IP4_0|_TX|4 _PTL_IP4_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP4_0|_TX|B1 0 _PTL_IP4_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP4_0|_TX|B2 0 _PTL_IP4_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP4_0|_TX|B1 _PTL_IP4_0|_TX|1 _PTL_IP4_0|_TX|3  1.684e-12
L_PTL_IP4_0|_TX|B2 _PTL_IP4_0|_TX|4 _PTL_IP4_0|_TX|6  3.596e-12
L_PTL_IP4_0|_TX|1 IP4_0 _PTL_IP4_0|_TX|1  2.063e-12
L_PTL_IP4_0|_TX|2 _PTL_IP4_0|_TX|1 _PTL_IP4_0|_TX|4  4.123e-12
L_PTL_IP4_0|_TX|3 _PTL_IP4_0|_TX|4 _PTL_IP4_0|_TX|7  2.193e-12
R_PTL_IP4_0|_TX|D _PTL_IP4_0|_TX|7 _PTL_IP4_0|A_PTL  1.36
L_PTL_IP4_0|_TX|P1 _PTL_IP4_0|_TX|2 0  5.254e-13
L_PTL_IP4_0|_TX|P2 _PTL_IP4_0|_TX|5 0  5.141e-13
R_PTL_IP4_0|_TX|B1 _PTL_IP4_0|_TX|1 _PTL_IP4_0|_TX|101  2.7439617672
R_PTL_IP4_0|_TX|B2 _PTL_IP4_0|_TX|4 _PTL_IP4_0|_TX|104  2.7439617672
L_PTL_IP4_0|_TX|RB1 _PTL_IP4_0|_TX|101 0  1.550338398468e-12
L_PTL_IP4_0|_TX|RB2 _PTL_IP4_0|_TX|104 0  1.550338398468e-12
B_PTL_IP4_0|_RX|1 _PTL_IP4_0|_RX|1 _PTL_IP4_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP4_0|_RX|2 _PTL_IP4_0|_RX|4 _PTL_IP4_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP4_0|_RX|3 _PTL_IP4_0|_RX|7 _PTL_IP4_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP4_0|_RX|B1 0 _PTL_IP4_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP4_0|_RX|B1 _PTL_IP4_0|_RX|1 _PTL_IP4_0|_RX|3  2.777e-12
I_PTL_IP4_0|_RX|B2 0 _PTL_IP4_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP4_0|_RX|B2 _PTL_IP4_0|_RX|4 _PTL_IP4_0|_RX|6  2.685e-12
I_PTL_IP4_0|_RX|B3 0 _PTL_IP4_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP4_0|_RX|B3 _PTL_IP4_0|_RX|7 _PTL_IP4_0|_RX|9  2.764e-12
L_PTL_IP4_0|_RX|1 _PTL_IP4_0|A_PTL _PTL_IP4_0|_RX|1  1.346e-12
L_PTL_IP4_0|_RX|2 _PTL_IP4_0|_RX|1 _PTL_IP4_0|_RX|4  6.348e-12
L_PTL_IP4_0|_RX|3 _PTL_IP4_0|_RX|4 _PTL_IP4_0|_RX|7  5.197e-12
L_PTL_IP4_0|_RX|4 _PTL_IP4_0|_RX|7 _PTL_IP4_0|D  2.058e-12
L_PTL_IP4_0|_RX|P1 _PTL_IP4_0|_RX|2 0  4.795e-13
L_PTL_IP4_0|_RX|P2 _PTL_IP4_0|_RX|5 0  5.431e-13
L_PTL_IP4_0|_RX|P3 _PTL_IP4_0|_RX|8 0  5.339e-13
R_PTL_IP4_0|_RX|B1 _PTL_IP4_0|_RX|1 _PTL_IP4_0|_RX|101  4.225701121488
R_PTL_IP4_0|_RX|B2 _PTL_IP4_0|_RX|4 _PTL_IP4_0|_RX|104  3.429952209
R_PTL_IP4_0|_RX|B3 _PTL_IP4_0|_RX|7 _PTL_IP4_0|_RX|107  2.7439617672
L_PTL_IP4_0|_RX|RB1 _PTL_IP4_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP4_0|_RX|RB2 _PTL_IP4_0|_RX|104 0  1.937922998085e-12
L_PTL_IP4_0|_RX|RB3 _PTL_IP4_0|_RX|107 0  1.550338398468e-12
L_PTL_IP4_0|_SPL|1 _PTL_IP4_0|D _PTL_IP4_0|_SPL|D1  2e-12
L_PTL_IP4_0|_SPL|2 _PTL_IP4_0|_SPL|D1 _PTL_IP4_0|_SPL|D2  4.135667696e-12
L_PTL_IP4_0|_SPL|3 _PTL_IP4_0|_SPL|D2 _PTL_IP4_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP4_0|_SPL|4 _PTL_IP4_0|_SPL|JCT _PTL_IP4_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP4_0|_SPL|5 _PTL_IP4_0|_SPL|QA1 IP4_0_TO4  2e-12
L_PTL_IP4_0|_SPL|6 _PTL_IP4_0|_SPL|JCT _PTL_IP4_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP4_0|_SPL|7 _PTL_IP4_0|_SPL|QB1 IP4_0_TO5  2e-12
B_PTL_IG4_0|_TX|1 _PTL_IG4_0|_TX|1 _PTL_IG4_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG4_0|_TX|2 _PTL_IG4_0|_TX|4 _PTL_IG4_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG4_0|_TX|B1 0 _PTL_IG4_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG4_0|_TX|B2 0 _PTL_IG4_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG4_0|_TX|B1 _PTL_IG4_0|_TX|1 _PTL_IG4_0|_TX|3  1.684e-12
L_PTL_IG4_0|_TX|B2 _PTL_IG4_0|_TX|4 _PTL_IG4_0|_TX|6  3.596e-12
L_PTL_IG4_0|_TX|1 IG4_0 _PTL_IG4_0|_TX|1  2.063e-12
L_PTL_IG4_0|_TX|2 _PTL_IG4_0|_TX|1 _PTL_IG4_0|_TX|4  4.123e-12
L_PTL_IG4_0|_TX|3 _PTL_IG4_0|_TX|4 _PTL_IG4_0|_TX|7  2.193e-12
R_PTL_IG4_0|_TX|D _PTL_IG4_0|_TX|7 _PTL_IG4_0|A_PTL  1.36
L_PTL_IG4_0|_TX|P1 _PTL_IG4_0|_TX|2 0  5.254e-13
L_PTL_IG4_0|_TX|P2 _PTL_IG4_0|_TX|5 0  5.141e-13
R_PTL_IG4_0|_TX|B1 _PTL_IG4_0|_TX|1 _PTL_IG4_0|_TX|101  2.7439617672
R_PTL_IG4_0|_TX|B2 _PTL_IG4_0|_TX|4 _PTL_IG4_0|_TX|104  2.7439617672
L_PTL_IG4_0|_TX|RB1 _PTL_IG4_0|_TX|101 0  1.550338398468e-12
L_PTL_IG4_0|_TX|RB2 _PTL_IG4_0|_TX|104 0  1.550338398468e-12
B_PTL_IG4_0|_RX|1 _PTL_IG4_0|_RX|1 _PTL_IG4_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG4_0|_RX|2 _PTL_IG4_0|_RX|4 _PTL_IG4_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG4_0|_RX|3 _PTL_IG4_0|_RX|7 _PTL_IG4_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG4_0|_RX|B1 0 _PTL_IG4_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG4_0|_RX|B1 _PTL_IG4_0|_RX|1 _PTL_IG4_0|_RX|3  2.777e-12
I_PTL_IG4_0|_RX|B2 0 _PTL_IG4_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG4_0|_RX|B2 _PTL_IG4_0|_RX|4 _PTL_IG4_0|_RX|6  2.685e-12
I_PTL_IG4_0|_RX|B3 0 _PTL_IG4_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG4_0|_RX|B3 _PTL_IG4_0|_RX|7 _PTL_IG4_0|_RX|9  2.764e-12
L_PTL_IG4_0|_RX|1 _PTL_IG4_0|A_PTL _PTL_IG4_0|_RX|1  1.346e-12
L_PTL_IG4_0|_RX|2 _PTL_IG4_0|_RX|1 _PTL_IG4_0|_RX|4  6.348e-12
L_PTL_IG4_0|_RX|3 _PTL_IG4_0|_RX|4 _PTL_IG4_0|_RX|7  5.197e-12
L_PTL_IG4_0|_RX|4 _PTL_IG4_0|_RX|7 _PTL_IG4_0|D  2.058e-12
L_PTL_IG4_0|_RX|P1 _PTL_IG4_0|_RX|2 0  4.795e-13
L_PTL_IG4_0|_RX|P2 _PTL_IG4_0|_RX|5 0  5.431e-13
L_PTL_IG4_0|_RX|P3 _PTL_IG4_0|_RX|8 0  5.339e-13
R_PTL_IG4_0|_RX|B1 _PTL_IG4_0|_RX|1 _PTL_IG4_0|_RX|101  4.225701121488
R_PTL_IG4_0|_RX|B2 _PTL_IG4_0|_RX|4 _PTL_IG4_0|_RX|104  3.429952209
R_PTL_IG4_0|_RX|B3 _PTL_IG4_0|_RX|7 _PTL_IG4_0|_RX|107  2.7439617672
L_PTL_IG4_0|_RX|RB1 _PTL_IG4_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG4_0|_RX|RB2 _PTL_IG4_0|_RX|104 0  1.937922998085e-12
L_PTL_IG4_0|_RX|RB3 _PTL_IG4_0|_RX|107 0  1.550338398468e-12
L_PTL_IG4_0|_SPL|1 _PTL_IG4_0|D _PTL_IG4_0|_SPL|D1  2e-12
L_PTL_IG4_0|_SPL|2 _PTL_IG4_0|_SPL|D1 _PTL_IG4_0|_SPL|D2  4.135667696e-12
L_PTL_IG4_0|_SPL|3 _PTL_IG4_0|_SPL|D2 _PTL_IG4_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IG4_0|_SPL|4 _PTL_IG4_0|_SPL|JCT _PTL_IG4_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IG4_0|_SPL|5 _PTL_IG4_0|_SPL|QA1 IG4_0_TO4  2e-12
L_PTL_IG4_0|_SPL|6 _PTL_IG4_0|_SPL|JCT _PTL_IG4_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IG4_0|_SPL|7 _PTL_IG4_0|_SPL|QB1 IG4_0_TO5  2e-12
B_PTL_IP5_0|_TX|1 _PTL_IP5_0|_TX|1 _PTL_IP5_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP5_0|_TX|2 _PTL_IP5_0|_TX|4 _PTL_IP5_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP5_0|_TX|B1 0 _PTL_IP5_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP5_0|_TX|B2 0 _PTL_IP5_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_0|_TX|B1 _PTL_IP5_0|_TX|1 _PTL_IP5_0|_TX|3  1.684e-12
L_PTL_IP5_0|_TX|B2 _PTL_IP5_0|_TX|4 _PTL_IP5_0|_TX|6  3.596e-12
L_PTL_IP5_0|_TX|1 IP5_0 _PTL_IP5_0|_TX|1  2.063e-12
L_PTL_IP5_0|_TX|2 _PTL_IP5_0|_TX|1 _PTL_IP5_0|_TX|4  4.123e-12
L_PTL_IP5_0|_TX|3 _PTL_IP5_0|_TX|4 _PTL_IP5_0|_TX|7  2.193e-12
R_PTL_IP5_0|_TX|D _PTL_IP5_0|_TX|7 _PTL_IP5_0|A_PTL  1.36
L_PTL_IP5_0|_TX|P1 _PTL_IP5_0|_TX|2 0  5.254e-13
L_PTL_IP5_0|_TX|P2 _PTL_IP5_0|_TX|5 0  5.141e-13
R_PTL_IP5_0|_TX|B1 _PTL_IP5_0|_TX|1 _PTL_IP5_0|_TX|101  2.7439617672
R_PTL_IP5_0|_TX|B2 _PTL_IP5_0|_TX|4 _PTL_IP5_0|_TX|104  2.7439617672
L_PTL_IP5_0|_TX|RB1 _PTL_IP5_0|_TX|101 0  1.550338398468e-12
L_PTL_IP5_0|_TX|RB2 _PTL_IP5_0|_TX|104 0  1.550338398468e-12
B_PTL_IP5_0|_RX|1 _PTL_IP5_0|_RX|1 _PTL_IP5_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP5_0|_RX|2 _PTL_IP5_0|_RX|4 _PTL_IP5_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP5_0|_RX|3 _PTL_IP5_0|_RX|7 _PTL_IP5_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP5_0|_RX|B1 0 _PTL_IP5_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP5_0|_RX|B1 _PTL_IP5_0|_RX|1 _PTL_IP5_0|_RX|3  2.777e-12
I_PTL_IP5_0|_RX|B2 0 _PTL_IP5_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP5_0|_RX|B2 _PTL_IP5_0|_RX|4 _PTL_IP5_0|_RX|6  2.685e-12
I_PTL_IP5_0|_RX|B3 0 _PTL_IP5_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_0|_RX|B3 _PTL_IP5_0|_RX|7 _PTL_IP5_0|_RX|9  2.764e-12
L_PTL_IP5_0|_RX|1 _PTL_IP5_0|A_PTL _PTL_IP5_0|_RX|1  1.346e-12
L_PTL_IP5_0|_RX|2 _PTL_IP5_0|_RX|1 _PTL_IP5_0|_RX|4  6.348e-12
L_PTL_IP5_0|_RX|3 _PTL_IP5_0|_RX|4 _PTL_IP5_0|_RX|7  5.197e-12
L_PTL_IP5_0|_RX|4 _PTL_IP5_0|_RX|7 _PTL_IP5_0|D  2.058e-12
L_PTL_IP5_0|_RX|P1 _PTL_IP5_0|_RX|2 0  4.795e-13
L_PTL_IP5_0|_RX|P2 _PTL_IP5_0|_RX|5 0  5.431e-13
L_PTL_IP5_0|_RX|P3 _PTL_IP5_0|_RX|8 0  5.339e-13
R_PTL_IP5_0|_RX|B1 _PTL_IP5_0|_RX|1 _PTL_IP5_0|_RX|101  4.225701121488
R_PTL_IP5_0|_RX|B2 _PTL_IP5_0|_RX|4 _PTL_IP5_0|_RX|104  3.429952209
R_PTL_IP5_0|_RX|B3 _PTL_IP5_0|_RX|7 _PTL_IP5_0|_RX|107  2.7439617672
L_PTL_IP5_0|_RX|RB1 _PTL_IP5_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP5_0|_RX|RB2 _PTL_IP5_0|_RX|104 0  1.937922998085e-12
L_PTL_IP5_0|_RX|RB3 _PTL_IP5_0|_RX|107 0  1.550338398468e-12
L_PTL_IP5_0|_SPL|1 _PTL_IP5_0|D _PTL_IP5_0|_SPL|D1  2e-12
L_PTL_IP5_0|_SPL|2 _PTL_IP5_0|_SPL|D1 _PTL_IP5_0|_SPL|D2  4.135667696e-12
L_PTL_IP5_0|_SPL|3 _PTL_IP5_0|_SPL|D2 _PTL_IP5_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP5_0|_SPL|4 _PTL_IP5_0|_SPL|JCT _PTL_IP5_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP5_0|_SPL|5 _PTL_IP5_0|_SPL|QA1 IP5_0_TO5  2e-12
L_PTL_IP5_0|_SPL|6 _PTL_IP5_0|_SPL|JCT _PTL_IP5_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP5_0|_SPL|7 _PTL_IP5_0|_SPL|QB1 IP5_0_OUT  2e-12
B_PTL_IG5_0|_TX|1 _PTL_IG5_0|_TX|1 _PTL_IG5_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG5_0|_TX|2 _PTL_IG5_0|_TX|4 _PTL_IG5_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG5_0|_TX|B1 0 _PTL_IG5_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG5_0|_TX|B2 0 _PTL_IG5_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG5_0|_TX|B1 _PTL_IG5_0|_TX|1 _PTL_IG5_0|_TX|3  1.684e-12
L_PTL_IG5_0|_TX|B2 _PTL_IG5_0|_TX|4 _PTL_IG5_0|_TX|6  3.596e-12
L_PTL_IG5_0|_TX|1 IG5_0 _PTL_IG5_0|_TX|1  2.063e-12
L_PTL_IG5_0|_TX|2 _PTL_IG5_0|_TX|1 _PTL_IG5_0|_TX|4  4.123e-12
L_PTL_IG5_0|_TX|3 _PTL_IG5_0|_TX|4 _PTL_IG5_0|_TX|7  2.193e-12
R_PTL_IG5_0|_TX|D _PTL_IG5_0|_TX|7 _PTL_IG5_0|A_PTL  1.36
L_PTL_IG5_0|_TX|P1 _PTL_IG5_0|_TX|2 0  5.254e-13
L_PTL_IG5_0|_TX|P2 _PTL_IG5_0|_TX|5 0  5.141e-13
R_PTL_IG5_0|_TX|B1 _PTL_IG5_0|_TX|1 _PTL_IG5_0|_TX|101  2.7439617672
R_PTL_IG5_0|_TX|B2 _PTL_IG5_0|_TX|4 _PTL_IG5_0|_TX|104  2.7439617672
L_PTL_IG5_0|_TX|RB1 _PTL_IG5_0|_TX|101 0  1.550338398468e-12
L_PTL_IG5_0|_TX|RB2 _PTL_IG5_0|_TX|104 0  1.550338398468e-12
B_PTL_IG5_0|_RX|1 _PTL_IG5_0|_RX|1 _PTL_IG5_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG5_0|_RX|2 _PTL_IG5_0|_RX|4 _PTL_IG5_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG5_0|_RX|3 _PTL_IG5_0|_RX|7 _PTL_IG5_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG5_0|_RX|B1 0 _PTL_IG5_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG5_0|_RX|B1 _PTL_IG5_0|_RX|1 _PTL_IG5_0|_RX|3  2.777e-12
I_PTL_IG5_0|_RX|B2 0 _PTL_IG5_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG5_0|_RX|B2 _PTL_IG5_0|_RX|4 _PTL_IG5_0|_RX|6  2.685e-12
I_PTL_IG5_0|_RX|B3 0 _PTL_IG5_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG5_0|_RX|B3 _PTL_IG5_0|_RX|7 _PTL_IG5_0|_RX|9  2.764e-12
L_PTL_IG5_0|_RX|1 _PTL_IG5_0|A_PTL _PTL_IG5_0|_RX|1  1.346e-12
L_PTL_IG5_0|_RX|2 _PTL_IG5_0|_RX|1 _PTL_IG5_0|_RX|4  6.348e-12
L_PTL_IG5_0|_RX|3 _PTL_IG5_0|_RX|4 _PTL_IG5_0|_RX|7  5.197e-12
L_PTL_IG5_0|_RX|4 _PTL_IG5_0|_RX|7 IG5_0_TO5  2.058e-12
L_PTL_IG5_0|_RX|P1 _PTL_IG5_0|_RX|2 0  4.795e-13
L_PTL_IG5_0|_RX|P2 _PTL_IG5_0|_RX|5 0  5.431e-13
L_PTL_IG5_0|_RX|P3 _PTL_IG5_0|_RX|8 0  5.339e-13
R_PTL_IG5_0|_RX|B1 _PTL_IG5_0|_RX|1 _PTL_IG5_0|_RX|101  4.225701121488
R_PTL_IG5_0|_RX|B2 _PTL_IG5_0|_RX|4 _PTL_IG5_0|_RX|104  3.429952209
R_PTL_IG5_0|_RX|B3 _PTL_IG5_0|_RX|7 _PTL_IG5_0|_RX|107  2.7439617672
L_PTL_IG5_0|_RX|RB1 _PTL_IG5_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG5_0|_RX|RB2 _PTL_IG5_0|_RX|104 0  1.937922998085e-12
L_PTL_IG5_0|_RX|RB3 _PTL_IG5_0|_RX|107 0  1.550338398468e-12
B_PTL_IP6_0|_TX|1 _PTL_IP6_0|_TX|1 _PTL_IP6_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP6_0|_TX|2 _PTL_IP6_0|_TX|4 _PTL_IP6_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP6_0|_TX|B1 0 _PTL_IP6_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP6_0|_TX|B2 0 _PTL_IP6_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP6_0|_TX|B1 _PTL_IP6_0|_TX|1 _PTL_IP6_0|_TX|3  1.684e-12
L_PTL_IP6_0|_TX|B2 _PTL_IP6_0|_TX|4 _PTL_IP6_0|_TX|6  3.596e-12
L_PTL_IP6_0|_TX|1 IP6_0 _PTL_IP6_0|_TX|1  2.063e-12
L_PTL_IP6_0|_TX|2 _PTL_IP6_0|_TX|1 _PTL_IP6_0|_TX|4  4.123e-12
L_PTL_IP6_0|_TX|3 _PTL_IP6_0|_TX|4 _PTL_IP6_0|_TX|7  2.193e-12
R_PTL_IP6_0|_TX|D _PTL_IP6_0|_TX|7 _PTL_IP6_0|A_PTL  1.36
L_PTL_IP6_0|_TX|P1 _PTL_IP6_0|_TX|2 0  5.254e-13
L_PTL_IP6_0|_TX|P2 _PTL_IP6_0|_TX|5 0  5.141e-13
R_PTL_IP6_0|_TX|B1 _PTL_IP6_0|_TX|1 _PTL_IP6_0|_TX|101  2.7439617672
R_PTL_IP6_0|_TX|B2 _PTL_IP6_0|_TX|4 _PTL_IP6_0|_TX|104  2.7439617672
L_PTL_IP6_0|_TX|RB1 _PTL_IP6_0|_TX|101 0  1.550338398468e-12
L_PTL_IP6_0|_TX|RB2 _PTL_IP6_0|_TX|104 0  1.550338398468e-12
B_PTL_IP6_0|_RX|1 _PTL_IP6_0|_RX|1 _PTL_IP6_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP6_0|_RX|2 _PTL_IP6_0|_RX|4 _PTL_IP6_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP6_0|_RX|3 _PTL_IP6_0|_RX|7 _PTL_IP6_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP6_0|_RX|B1 0 _PTL_IP6_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP6_0|_RX|B1 _PTL_IP6_0|_RX|1 _PTL_IP6_0|_RX|3  2.777e-12
I_PTL_IP6_0|_RX|B2 0 _PTL_IP6_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP6_0|_RX|B2 _PTL_IP6_0|_RX|4 _PTL_IP6_0|_RX|6  2.685e-12
I_PTL_IP6_0|_RX|B3 0 _PTL_IP6_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP6_0|_RX|B3 _PTL_IP6_0|_RX|7 _PTL_IP6_0|_RX|9  2.764e-12
L_PTL_IP6_0|_RX|1 _PTL_IP6_0|A_PTL _PTL_IP6_0|_RX|1  1.346e-12
L_PTL_IP6_0|_RX|2 _PTL_IP6_0|_RX|1 _PTL_IP6_0|_RX|4  6.348e-12
L_PTL_IP6_0|_RX|3 _PTL_IP6_0|_RX|4 _PTL_IP6_0|_RX|7  5.197e-12
L_PTL_IP6_0|_RX|4 _PTL_IP6_0|_RX|7 _PTL_IP6_0|D  2.058e-12
L_PTL_IP6_0|_RX|P1 _PTL_IP6_0|_RX|2 0  4.795e-13
L_PTL_IP6_0|_RX|P2 _PTL_IP6_0|_RX|5 0  5.431e-13
L_PTL_IP6_0|_RX|P3 _PTL_IP6_0|_RX|8 0  5.339e-13
R_PTL_IP6_0|_RX|B1 _PTL_IP6_0|_RX|1 _PTL_IP6_0|_RX|101  4.225701121488
R_PTL_IP6_0|_RX|B2 _PTL_IP6_0|_RX|4 _PTL_IP6_0|_RX|104  3.429952209
R_PTL_IP6_0|_RX|B3 _PTL_IP6_0|_RX|7 _PTL_IP6_0|_RX|107  2.7439617672
L_PTL_IP6_0|_RX|RB1 _PTL_IP6_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP6_0|_RX|RB2 _PTL_IP6_0|_RX|104 0  1.937922998085e-12
L_PTL_IP6_0|_RX|RB3 _PTL_IP6_0|_RX|107 0  1.550338398468e-12
L_PTL_IP6_0|_SPL|1 _PTL_IP6_0|D _PTL_IP6_0|_SPL|D1  2e-12
L_PTL_IP6_0|_SPL|2 _PTL_IP6_0|_SPL|D1 _PTL_IP6_0|_SPL|D2  4.135667696e-12
L_PTL_IP6_0|_SPL|3 _PTL_IP6_0|_SPL|D2 _PTL_IP6_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP6_0|_SPL|4 _PTL_IP6_0|_SPL|JCT _PTL_IP6_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP6_0|_SPL|5 _PTL_IP6_0|_SPL|QA1 IP6_0_TO6  2e-12
L_PTL_IP6_0|_SPL|6 _PTL_IP6_0|_SPL|JCT _PTL_IP6_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP6_0|_SPL|7 _PTL_IP6_0|_SPL|QB1 IP6_0_TO7  2e-12
B_PTL_IG6_0|_TX|1 _PTL_IG6_0|_TX|1 _PTL_IG6_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG6_0|_TX|2 _PTL_IG6_0|_TX|4 _PTL_IG6_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG6_0|_TX|B1 0 _PTL_IG6_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG6_0|_TX|B2 0 _PTL_IG6_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG6_0|_TX|B1 _PTL_IG6_0|_TX|1 _PTL_IG6_0|_TX|3  1.684e-12
L_PTL_IG6_0|_TX|B2 _PTL_IG6_0|_TX|4 _PTL_IG6_0|_TX|6  3.596e-12
L_PTL_IG6_0|_TX|1 IG6_0 _PTL_IG6_0|_TX|1  2.063e-12
L_PTL_IG6_0|_TX|2 _PTL_IG6_0|_TX|1 _PTL_IG6_0|_TX|4  4.123e-12
L_PTL_IG6_0|_TX|3 _PTL_IG6_0|_TX|4 _PTL_IG6_0|_TX|7  2.193e-12
R_PTL_IG6_0|_TX|D _PTL_IG6_0|_TX|7 _PTL_IG6_0|A_PTL  1.36
L_PTL_IG6_0|_TX|P1 _PTL_IG6_0|_TX|2 0  5.254e-13
L_PTL_IG6_0|_TX|P2 _PTL_IG6_0|_TX|5 0  5.141e-13
R_PTL_IG6_0|_TX|B1 _PTL_IG6_0|_TX|1 _PTL_IG6_0|_TX|101  2.7439617672
R_PTL_IG6_0|_TX|B2 _PTL_IG6_0|_TX|4 _PTL_IG6_0|_TX|104  2.7439617672
L_PTL_IG6_0|_TX|RB1 _PTL_IG6_0|_TX|101 0  1.550338398468e-12
L_PTL_IG6_0|_TX|RB2 _PTL_IG6_0|_TX|104 0  1.550338398468e-12
B_PTL_IG6_0|_RX|1 _PTL_IG6_0|_RX|1 _PTL_IG6_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG6_0|_RX|2 _PTL_IG6_0|_RX|4 _PTL_IG6_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG6_0|_RX|3 _PTL_IG6_0|_RX|7 _PTL_IG6_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG6_0|_RX|B1 0 _PTL_IG6_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG6_0|_RX|B1 _PTL_IG6_0|_RX|1 _PTL_IG6_0|_RX|3  2.777e-12
I_PTL_IG6_0|_RX|B2 0 _PTL_IG6_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG6_0|_RX|B2 _PTL_IG6_0|_RX|4 _PTL_IG6_0|_RX|6  2.685e-12
I_PTL_IG6_0|_RX|B3 0 _PTL_IG6_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG6_0|_RX|B3 _PTL_IG6_0|_RX|7 _PTL_IG6_0|_RX|9  2.764e-12
L_PTL_IG6_0|_RX|1 _PTL_IG6_0|A_PTL _PTL_IG6_0|_RX|1  1.346e-12
L_PTL_IG6_0|_RX|2 _PTL_IG6_0|_RX|1 _PTL_IG6_0|_RX|4  6.348e-12
L_PTL_IG6_0|_RX|3 _PTL_IG6_0|_RX|4 _PTL_IG6_0|_RX|7  5.197e-12
L_PTL_IG6_0|_RX|4 _PTL_IG6_0|_RX|7 _PTL_IG6_0|D  2.058e-12
L_PTL_IG6_0|_RX|P1 _PTL_IG6_0|_RX|2 0  4.795e-13
L_PTL_IG6_0|_RX|P2 _PTL_IG6_0|_RX|5 0  5.431e-13
L_PTL_IG6_0|_RX|P3 _PTL_IG6_0|_RX|8 0  5.339e-13
R_PTL_IG6_0|_RX|B1 _PTL_IG6_0|_RX|1 _PTL_IG6_0|_RX|101  4.225701121488
R_PTL_IG6_0|_RX|B2 _PTL_IG6_0|_RX|4 _PTL_IG6_0|_RX|104  3.429952209
R_PTL_IG6_0|_RX|B3 _PTL_IG6_0|_RX|7 _PTL_IG6_0|_RX|107  2.7439617672
L_PTL_IG6_0|_RX|RB1 _PTL_IG6_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG6_0|_RX|RB2 _PTL_IG6_0|_RX|104 0  1.937922998085e-12
L_PTL_IG6_0|_RX|RB3 _PTL_IG6_0|_RX|107 0  1.550338398468e-12
L_PTL_IG6_0|_SPL|1 _PTL_IG6_0|D _PTL_IG6_0|_SPL|D1  2e-12
L_PTL_IG6_0|_SPL|2 _PTL_IG6_0|_SPL|D1 _PTL_IG6_0|_SPL|D2  4.135667696e-12
L_PTL_IG6_0|_SPL|3 _PTL_IG6_0|_SPL|D2 _PTL_IG6_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IG6_0|_SPL|4 _PTL_IG6_0|_SPL|JCT _PTL_IG6_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IG6_0|_SPL|5 _PTL_IG6_0|_SPL|QA1 IG6_0_TO6  2e-12
L_PTL_IG6_0|_SPL|6 _PTL_IG6_0|_SPL|JCT _PTL_IG6_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IG6_0|_SPL|7 _PTL_IG6_0|_SPL|QB1 IG6_0_TO7  2e-12
B_PTL_IP7_0|_TX|1 _PTL_IP7_0|_TX|1 _PTL_IP7_0|_TX|2 JJMIT AREA=2.5
B_PTL_IP7_0|_TX|2 _PTL_IP7_0|_TX|4 _PTL_IP7_0|_TX|5 JJMIT AREA=2.5
I_PTL_IP7_0|_TX|B1 0 _PTL_IP7_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP7_0|_TX|B2 0 _PTL_IP7_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_0|_TX|B1 _PTL_IP7_0|_TX|1 _PTL_IP7_0|_TX|3  1.684e-12
L_PTL_IP7_0|_TX|B2 _PTL_IP7_0|_TX|4 _PTL_IP7_0|_TX|6  3.596e-12
L_PTL_IP7_0|_TX|1 IP7_0 _PTL_IP7_0|_TX|1  2.063e-12
L_PTL_IP7_0|_TX|2 _PTL_IP7_0|_TX|1 _PTL_IP7_0|_TX|4  4.123e-12
L_PTL_IP7_0|_TX|3 _PTL_IP7_0|_TX|4 _PTL_IP7_0|_TX|7  2.193e-12
R_PTL_IP7_0|_TX|D _PTL_IP7_0|_TX|7 _PTL_IP7_0|A_PTL  1.36
L_PTL_IP7_0|_TX|P1 _PTL_IP7_0|_TX|2 0  5.254e-13
L_PTL_IP7_0|_TX|P2 _PTL_IP7_0|_TX|5 0  5.141e-13
R_PTL_IP7_0|_TX|B1 _PTL_IP7_0|_TX|1 _PTL_IP7_0|_TX|101  2.7439617672
R_PTL_IP7_0|_TX|B2 _PTL_IP7_0|_TX|4 _PTL_IP7_0|_TX|104  2.7439617672
L_PTL_IP7_0|_TX|RB1 _PTL_IP7_0|_TX|101 0  1.550338398468e-12
L_PTL_IP7_0|_TX|RB2 _PTL_IP7_0|_TX|104 0  1.550338398468e-12
B_PTL_IP7_0|_RX|1 _PTL_IP7_0|_RX|1 _PTL_IP7_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP7_0|_RX|2 _PTL_IP7_0|_RX|4 _PTL_IP7_0|_RX|5 JJMIT AREA=2.0
B_PTL_IP7_0|_RX|3 _PTL_IP7_0|_RX|7 _PTL_IP7_0|_RX|8 JJMIT AREA=2.5
I_PTL_IP7_0|_RX|B1 0 _PTL_IP7_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP7_0|_RX|B1 _PTL_IP7_0|_RX|1 _PTL_IP7_0|_RX|3  2.777e-12
I_PTL_IP7_0|_RX|B2 0 _PTL_IP7_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP7_0|_RX|B2 _PTL_IP7_0|_RX|4 _PTL_IP7_0|_RX|6  2.685e-12
I_PTL_IP7_0|_RX|B3 0 _PTL_IP7_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_0|_RX|B3 _PTL_IP7_0|_RX|7 _PTL_IP7_0|_RX|9  2.764e-12
L_PTL_IP7_0|_RX|1 _PTL_IP7_0|A_PTL _PTL_IP7_0|_RX|1  1.346e-12
L_PTL_IP7_0|_RX|2 _PTL_IP7_0|_RX|1 _PTL_IP7_0|_RX|4  6.348e-12
L_PTL_IP7_0|_RX|3 _PTL_IP7_0|_RX|4 _PTL_IP7_0|_RX|7  5.197e-12
L_PTL_IP7_0|_RX|4 _PTL_IP7_0|_RX|7 _PTL_IP7_0|D  2.058e-12
L_PTL_IP7_0|_RX|P1 _PTL_IP7_0|_RX|2 0  4.795e-13
L_PTL_IP7_0|_RX|P2 _PTL_IP7_0|_RX|5 0  5.431e-13
L_PTL_IP7_0|_RX|P3 _PTL_IP7_0|_RX|8 0  5.339e-13
R_PTL_IP7_0|_RX|B1 _PTL_IP7_0|_RX|1 _PTL_IP7_0|_RX|101  4.225701121488
R_PTL_IP7_0|_RX|B2 _PTL_IP7_0|_RX|4 _PTL_IP7_0|_RX|104  3.429952209
R_PTL_IP7_0|_RX|B3 _PTL_IP7_0|_RX|7 _PTL_IP7_0|_RX|107  2.7439617672
L_PTL_IP7_0|_RX|RB1 _PTL_IP7_0|_RX|101 0  2.38752113364072e-12
L_PTL_IP7_0|_RX|RB2 _PTL_IP7_0|_RX|104 0  1.937922998085e-12
L_PTL_IP7_0|_RX|RB3 _PTL_IP7_0|_RX|107 0  1.550338398468e-12
L_PTL_IP7_0|_SPL|1 _PTL_IP7_0|D _PTL_IP7_0|_SPL|D1  2e-12
L_PTL_IP7_0|_SPL|2 _PTL_IP7_0|_SPL|D1 _PTL_IP7_0|_SPL|D2  4.135667696e-12
L_PTL_IP7_0|_SPL|3 _PTL_IP7_0|_SPL|D2 _PTL_IP7_0|_SPL|JCT  9.84682784761905e-13
L_PTL_IP7_0|_SPL|4 _PTL_IP7_0|_SPL|JCT _PTL_IP7_0|_SPL|QA1  9.84682784761905e-13
L_PTL_IP7_0|_SPL|5 _PTL_IP7_0|_SPL|QA1 IP7_0_TO7  2e-12
L_PTL_IP7_0|_SPL|6 _PTL_IP7_0|_SPL|JCT _PTL_IP7_0|_SPL|QB1  9.84682784761905e-13
L_PTL_IP7_0|_SPL|7 _PTL_IP7_0|_SPL|QB1 IP7_0_OUT  2e-12
B_PTL_IG7_0|_TX|1 _PTL_IG7_0|_TX|1 _PTL_IG7_0|_TX|2 JJMIT AREA=2.5
B_PTL_IG7_0|_TX|2 _PTL_IG7_0|_TX|4 _PTL_IG7_0|_TX|5 JJMIT AREA=2.5
I_PTL_IG7_0|_TX|B1 0 _PTL_IG7_0|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IG7_0|_TX|B2 0 _PTL_IG7_0|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IG7_0|_TX|B1 _PTL_IG7_0|_TX|1 _PTL_IG7_0|_TX|3  1.684e-12
L_PTL_IG7_0|_TX|B2 _PTL_IG7_0|_TX|4 _PTL_IG7_0|_TX|6  3.596e-12
L_PTL_IG7_0|_TX|1 IG7_0 _PTL_IG7_0|_TX|1  2.063e-12
L_PTL_IG7_0|_TX|2 _PTL_IG7_0|_TX|1 _PTL_IG7_0|_TX|4  4.123e-12
L_PTL_IG7_0|_TX|3 _PTL_IG7_0|_TX|4 _PTL_IG7_0|_TX|7  2.193e-12
R_PTL_IG7_0|_TX|D _PTL_IG7_0|_TX|7 _PTL_IG7_0|A_PTL  1.36
L_PTL_IG7_0|_TX|P1 _PTL_IG7_0|_TX|2 0  5.254e-13
L_PTL_IG7_0|_TX|P2 _PTL_IG7_0|_TX|5 0  5.141e-13
R_PTL_IG7_0|_TX|B1 _PTL_IG7_0|_TX|1 _PTL_IG7_0|_TX|101  2.7439617672
R_PTL_IG7_0|_TX|B2 _PTL_IG7_0|_TX|4 _PTL_IG7_0|_TX|104  2.7439617672
L_PTL_IG7_0|_TX|RB1 _PTL_IG7_0|_TX|101 0  1.550338398468e-12
L_PTL_IG7_0|_TX|RB2 _PTL_IG7_0|_TX|104 0  1.550338398468e-12
B_PTL_IG7_0|_RX|1 _PTL_IG7_0|_RX|1 _PTL_IG7_0|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IG7_0|_RX|2 _PTL_IG7_0|_RX|4 _PTL_IG7_0|_RX|5 JJMIT AREA=2.0
B_PTL_IG7_0|_RX|3 _PTL_IG7_0|_RX|7 _PTL_IG7_0|_RX|8 JJMIT AREA=2.5
I_PTL_IG7_0|_RX|B1 0 _PTL_IG7_0|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IG7_0|_RX|B1 _PTL_IG7_0|_RX|1 _PTL_IG7_0|_RX|3  2.777e-12
I_PTL_IG7_0|_RX|B2 0 _PTL_IG7_0|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IG7_0|_RX|B2 _PTL_IG7_0|_RX|4 _PTL_IG7_0|_RX|6  2.685e-12
I_PTL_IG7_0|_RX|B3 0 _PTL_IG7_0|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IG7_0|_RX|B3 _PTL_IG7_0|_RX|7 _PTL_IG7_0|_RX|9  2.764e-12
L_PTL_IG7_0|_RX|1 _PTL_IG7_0|A_PTL _PTL_IG7_0|_RX|1  1.346e-12
L_PTL_IG7_0|_RX|2 _PTL_IG7_0|_RX|1 _PTL_IG7_0|_RX|4  6.348e-12
L_PTL_IG7_0|_RX|3 _PTL_IG7_0|_RX|4 _PTL_IG7_0|_RX|7  5.197e-12
L_PTL_IG7_0|_RX|4 _PTL_IG7_0|_RX|7 IG7_0_TO7  2.058e-12
L_PTL_IG7_0|_RX|P1 _PTL_IG7_0|_RX|2 0  4.795e-13
L_PTL_IG7_0|_RX|P2 _PTL_IG7_0|_RX|5 0  5.431e-13
L_PTL_IG7_0|_RX|P3 _PTL_IG7_0|_RX|8 0  5.339e-13
R_PTL_IG7_0|_RX|B1 _PTL_IG7_0|_RX|1 _PTL_IG7_0|_RX|101  4.225701121488
R_PTL_IG7_0|_RX|B2 _PTL_IG7_0|_RX|4 _PTL_IG7_0|_RX|104  3.429952209
R_PTL_IG7_0|_RX|B3 _PTL_IG7_0|_RX|7 _PTL_IG7_0|_RX|107  2.7439617672
L_PTL_IG7_0|_RX|RB1 _PTL_IG7_0|_RX|101 0  2.38752113364072e-12
L_PTL_IG7_0|_RX|RB2 _PTL_IG7_0|_RX|104 0  1.937922998085e-12
L_PTL_IG7_0|_RX|RB3 _PTL_IG7_0|_RX|107 0  1.550338398468e-12
L_S0_01|I_1|B _S0_01|A1 _S0_01|I_1|MID  2e-12
I_S0_01|I_1|B 0 _S0_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0_01|I_3|B _S0_01|A3 _S0_01|I_3|MID  2e-12
I_S0_01|I_3|B 0 _S0_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0_01|I_T|B _S0_01|T1 _S0_01|I_T|MID  2e-12
I_S0_01|I_T|B 0 _S0_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0_01|I_6|B _S0_01|Q1 _S0_01|I_6|MID  2e-12
I_S0_01|I_6|B 0 _S0_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0_01|1|1 _S0_01|A1 _S0_01|1|MID_SERIES JJMIT AREA=2.5
L_S0_01|1|P _S0_01|1|MID_SERIES 0  2e-13
R_S0_01|1|B _S0_01|A1 _S0_01|1|MID_SHUNT  2.7439617672
L_S0_01|1|RB _S0_01|1|MID_SHUNT 0  1.550338398468e-12
B_S0_01|23|1 _S0_01|A2 _S0_01|A3 JJMIT AREA=1.7857142857142858
R_S0_01|23|B _S0_01|A2 _S0_01|23|MID_SHUNT  3.84154647408
L_S0_01|23|RB _S0_01|23|MID_SHUNT _S0_01|A3  2.1704737578552e-12
B_S0_01|3|1 _S0_01|A3 _S0_01|3|MID_SERIES JJMIT AREA=2.5
L_S0_01|3|P _S0_01|3|MID_SERIES 0  2e-13
R_S0_01|3|B _S0_01|A3 _S0_01|3|MID_SHUNT  2.7439617672
L_S0_01|3|RB _S0_01|3|MID_SHUNT 0  1.550338398468e-12
B_S0_01|4|1 _S0_01|A4 _S0_01|4|MID_SERIES JJMIT AREA=2.5
L_S0_01|4|P _S0_01|4|MID_SERIES 0  2e-13
R_S0_01|4|B _S0_01|A4 _S0_01|4|MID_SHUNT  2.7439617672
L_S0_01|4|RB _S0_01|4|MID_SHUNT 0  1.550338398468e-12
B_S0_01|T|1 _S0_01|T1 _S0_01|T|MID_SERIES JJMIT AREA=2.5
L_S0_01|T|P _S0_01|T|MID_SERIES 0  2e-13
R_S0_01|T|B _S0_01|T1 _S0_01|T|MID_SHUNT  2.7439617672
L_S0_01|T|RB _S0_01|T|MID_SHUNT 0  1.550338398468e-12
B_S0_01|45|1 _S0_01|T2 _S0_01|A4 JJMIT AREA=1.7857142857142858
R_S0_01|45|B _S0_01|T2 _S0_01|45|MID_SHUNT  3.84154647408
L_S0_01|45|RB _S0_01|45|MID_SHUNT _S0_01|A4  2.1704737578552e-12
B_S0_01|6|1 _S0_01|Q1 _S0_01|6|MID_SERIES JJMIT AREA=2.5
L_S0_01|6|P _S0_01|6|MID_SERIES 0  2e-13
R_S0_01|6|B _S0_01|Q1 _S0_01|6|MID_SHUNT  2.7439617672
L_S0_01|6|RB _S0_01|6|MID_SHUNT 0  1.550338398468e-12
L_S1_01|I_A1|B _S1_01|A1 _S1_01|I_A1|MID  2e-12
I_S1_01|I_A1|B 0 _S1_01|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S1_01|I_A3|B _S1_01|A3 _S1_01|I_A3|MID  2e-12
I_S1_01|I_A3|B 0 _S1_01|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S1_01|I_B1|B _S1_01|B1 _S1_01|I_B1|MID  2e-12
I_S1_01|I_B1|B 0 _S1_01|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S1_01|I_B3|B _S1_01|B3 _S1_01|I_B3|MID  2e-12
I_S1_01|I_B3|B 0 _S1_01|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S1_01|I_Q1|B _S1_01|Q1 _S1_01|I_Q1|MID  2e-12
I_S1_01|I_Q1|B 0 _S1_01|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S1_01|A1|1 _S1_01|A1 _S1_01|A1|MID_SERIES JJMIT AREA=2.5
L_S1_01|A1|P _S1_01|A1|MID_SERIES 0  5e-13
R_S1_01|A1|B _S1_01|A1 _S1_01|A1|MID_SHUNT  2.7439617672
L_S1_01|A1|RB _S1_01|A1|MID_SHUNT 0  2.050338398468e-12
B_S1_01|A2|1 _S1_01|A2 _S1_01|A2|MID_SERIES JJMIT AREA=2.5
L_S1_01|A2|P _S1_01|A2|MID_SERIES 0  5e-13
R_S1_01|A2|B _S1_01|A2 _S1_01|A2|MID_SHUNT  2.7439617672
L_S1_01|A2|RB _S1_01|A2|MID_SHUNT 0  2.050338398468e-12
B_S1_01|A3|1 _S1_01|A2 _S1_01|A3|MID_SERIES JJMIT AREA=2.5
L_S1_01|A3|P _S1_01|A3|MID_SERIES _S1_01|A3  1.2e-12
R_S1_01|A3|B _S1_01|A2 _S1_01|A3|MID_SHUNT  2.7439617672
L_S1_01|A3|RB _S1_01|A3|MID_SHUNT _S1_01|A3  2.050338398468e-12
B_S1_01|B1|1 _S1_01|B1 _S1_01|B1|MID_SERIES JJMIT AREA=2.5
L_S1_01|B1|P _S1_01|B1|MID_SERIES 0  5e-13
R_S1_01|B1|B _S1_01|B1 _S1_01|B1|MID_SHUNT  2.7439617672
L_S1_01|B1|RB _S1_01|B1|MID_SHUNT 0  2.050338398468e-12
B_S1_01|B2|1 _S1_01|B2 _S1_01|B2|MID_SERIES JJMIT AREA=2.5
L_S1_01|B2|P _S1_01|B2|MID_SERIES 0  5e-13
R_S1_01|B2|B _S1_01|B2 _S1_01|B2|MID_SHUNT  2.7439617672
L_S1_01|B2|RB _S1_01|B2|MID_SHUNT 0  2.050338398468e-12
B_S1_01|B3|1 _S1_01|B2 _S1_01|B3|MID_SERIES JJMIT AREA=2.5
L_S1_01|B3|P _S1_01|B3|MID_SERIES _S1_01|B3  1.2e-12
R_S1_01|B3|B _S1_01|B2 _S1_01|B3|MID_SHUNT  2.7439617672
L_S1_01|B3|RB _S1_01|B3|MID_SHUNT _S1_01|B3  2.050338398468e-12
B_S1_01|T1|1 _S1_01|T1 _S1_01|T1|MID_SERIES JJMIT AREA=2.5
L_S1_01|T1|P _S1_01|T1|MID_SERIES 0  5e-13
R_S1_01|T1|B _S1_01|T1 _S1_01|T1|MID_SHUNT  2.7439617672
L_S1_01|T1|RB _S1_01|T1|MID_SHUNT 0  2.050338398468e-12
B_S1_01|T2|1 _S1_01|T2 _S1_01|ABTQ JJMIT AREA=2.0
R_S1_01|T2|B _S1_01|T2 _S1_01|T2|MID_SHUNT  3.429952209
L_S1_01|T2|RB _S1_01|T2|MID_SHUNT _S1_01|ABTQ  2.437922998085e-12
B_S1_01|AB|1 _S1_01|AB _S1_01|AB|MID_SERIES JJMIT AREA=1.5
L_S1_01|AB|P _S1_01|AB|MID_SERIES _S1_01|ABTQ  1.2e-12
R_S1_01|AB|B _S1_01|AB _S1_01|AB|MID_SHUNT  4.573269612
L_S1_01|AB|RB _S1_01|AB|MID_SHUNT _S1_01|ABTQ  3.08389733078e-12
B_S1_01|ABTQ|1 _S1_01|ABTQ _S1_01|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S1_01|ABTQ|P _S1_01|ABTQ|MID_SERIES 0  5e-13
R_S1_01|ABTQ|B _S1_01|ABTQ _S1_01|ABTQ|MID_SHUNT  3.6586156896
L_S1_01|ABTQ|RB _S1_01|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S1_01|Q1|1 _S1_01|Q1 _S1_01|Q1|MID_SERIES JJMIT AREA=2.5
L_S1_01|Q1|P _S1_01|Q1|MID_SERIES 0  5e-13
R_S1_01|Q1|B _S1_01|Q1 _S1_01|Q1|MID_SHUNT  2.7439617672
L_S1_01|Q1|RB _S1_01|Q1|MID_SHUNT 0  2.050338398468e-12
L_PG1_01|_SPL_G1|1 IG1_0_TO1 _PG1_01|_SPL_G1|D1  2e-12
L_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|D2  4.135667696e-12
L_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG1_01|_SPL_G1|5 _PG1_01|_SPL_G1|QA1 _PG1_01|G1_COPY_1  2e-12
L_PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|QB1 _PG1_01|G1_COPY_2  2e-12
L_PG1_01|_SPL_P1|1 IP1_0_TO1 _PG1_01|_SPL_P1|D1  2e-12
L_PG1_01|_SPL_P1|2 _PG1_01|_SPL_P1|D1 _PG1_01|_SPL_P1|D2  4.135667696e-12
L_PG1_01|_SPL_P1|3 _PG1_01|_SPL_P1|D2 _PG1_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG1_01|_SPL_P1|4 _PG1_01|_SPL_P1|JCT _PG1_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG1_01|_SPL_P1|5 _PG1_01|_SPL_P1|QA1 _PG1_01|P1_COPY_1  2e-12
L_PG1_01|_SPL_P1|6 _PG1_01|_SPL_P1|JCT _PG1_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG1_01|_SPL_P1|7 _PG1_01|_SPL_P1|QB1 _PG1_01|P1_COPY_2  2e-12
L_PG1_01|_PG|A1 _PG1_01|P1_COPY_1 _PG1_01|_PG|A1  2.067833848e-12
L_PG1_01|_PG|A2 _PG1_01|_PG|A1 _PG1_01|_PG|A2  4.135667696e-12
L_PG1_01|_PG|A3 _PG1_01|_PG|A3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|B1 _PG1_01|G1_COPY_1 _PG1_01|_PG|B1  2.067833848e-12
L_PG1_01|_PG|B2 _PG1_01|_PG|B1 _PG1_01|_PG|B2  4.135667696e-12
L_PG1_01|_PG|B3 _PG1_01|_PG|B3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|Q3 _PG1_01|_PG|Q3 _PG1_01|_PG|Q2  4.135667696e-12
L_PG1_01|_PG|Q2 _PG1_01|_PG|Q2 _PG1_01|_PG|Q1  4.135667696e-12
L_PG1_01|_PG|Q1 _PG1_01|_PG|Q1 _PG1_01|PG  2.067833848e-12
L_PG1_01|_GG|A1 IG0_0_TO1 _PG1_01|_GG|A1  2.067833848e-12
L_PG1_01|_GG|A2 _PG1_01|_GG|A1 _PG1_01|_GG|A2  4.135667696e-12
L_PG1_01|_GG|A3 _PG1_01|_GG|A3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|B1 _PG1_01|G1_COPY_2 _PG1_01|_GG|B1  2.067833848e-12
L_PG1_01|_GG|B2 _PG1_01|_GG|B1 _PG1_01|_GG|B2  4.135667696e-12
L_PG1_01|_GG|B3 _PG1_01|_GG|B3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|Q3 _PG1_01|_GG|Q3 _PG1_01|_GG|Q2  4.135667696e-12
L_PG1_01|_GG|Q2 _PG1_01|_GG|Q2 _PG1_01|_GG|Q1  4.135667696e-12
L_PG1_01|_GG|Q1 _PG1_01|_GG|Q1 _PG1_01|GG  2.067833848e-12
L_PG1_01|_DFF_P0|1 IP0_0_TO1 _PG1_01|_DFF_P0|A1  2.067833848e-12
L_PG1_01|_DFF_P0|2 _PG1_01|_DFF_P0|A1 _PG1_01|_DFF_P0|A2  4.135667696e-12
L_PG1_01|_DFF_P0|3 _PG1_01|_DFF_P0|A3 _PG1_01|_DFF_P0|A4  8.271335392e-12
L_PG1_01|_DFF_P0|T T12 _PG1_01|_DFF_P0|T1  2.067833848e-12
L_PG1_01|_DFF_P0|4 _PG1_01|_DFF_P0|T1 _PG1_01|_DFF_P0|T2  4.135667696e-12
L_PG1_01|_DFF_P0|5 _PG1_01|_DFF_P0|A4 _PG1_01|_DFF_P0|Q1  4.135667696e-12
L_PG1_01|_DFF_P0|6 _PG1_01|_DFF_P0|Q1 _PG1_01|P0_SYNC  2.067833848e-12
L_PG1_01|_DFF_P1|1 _PG1_01|P1_COPY_2 _PG1_01|_DFF_P1|A1  2.067833848e-12
L_PG1_01|_DFF_P1|2 _PG1_01|_DFF_P1|A1 _PG1_01|_DFF_P1|A2  4.135667696e-12
L_PG1_01|_DFF_P1|3 _PG1_01|_DFF_P1|A3 _PG1_01|_DFF_P1|A4  8.271335392e-12
L_PG1_01|_DFF_P1|T T12 _PG1_01|_DFF_P1|T1  2.067833848e-12
L_PG1_01|_DFF_P1|4 _PG1_01|_DFF_P1|T1 _PG1_01|_DFF_P1|T2  4.135667696e-12
L_PG1_01|_DFF_P1|5 _PG1_01|_DFF_P1|A4 _PG1_01|_DFF_P1|Q1  4.135667696e-12
L_PG1_01|_DFF_P1|6 _PG1_01|_DFF_P1|Q1 _PG1_01|P1_SYNC  2.067833848e-12
L_PG1_01|_DFF_PG|1 _PG1_01|PG _PG1_01|_DFF_PG|A1  2.067833848e-12
L_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|A2  4.135667696e-12
L_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|A4  8.271335392e-12
L_PG1_01|_DFF_PG|T T12 _PG1_01|_DFF_PG|T1  2.067833848e-12
L_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T2  4.135667696e-12
L_PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|Q1  4.135667696e-12
L_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|Q1 _PG1_01|PG_SYNC  2.067833848e-12
L_PG1_01|_DFF_GG|1 _PG1_01|GG _PG1_01|_DFF_GG|A1  2.067833848e-12
L_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|A2  4.135667696e-12
L_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|A4  8.271335392e-12
L_PG1_01|_DFF_GG|T T12 _PG1_01|_DFF_GG|T1  2.067833848e-12
L_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T2  4.135667696e-12
L_PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|Q1  4.135667696e-12
L_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|Q1 _PG1_01|GG_SYNC  2.067833848e-12
L_PG1_01|_AND_G|A1 _PG1_01|PG_SYNC _PG1_01|_AND_G|A1  2.067833848e-12
L_PG1_01|_AND_G|A2 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A2  4.135667696e-12
L_PG1_01|_AND_G|A3 _PG1_01|_AND_G|A3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|B1 _PG1_01|GG_SYNC _PG1_01|_AND_G|B1  2.067833848e-12
L_PG1_01|_AND_G|B2 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B2  4.135667696e-12
L_PG1_01|_AND_G|B3 _PG1_01|_AND_G|B3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q2  4.135667696e-12
L_PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q1  4.135667696e-12
L_PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1 G1_1_TX  2.067833848e-12
L_PG1_01|_AND_P|A1 _PG1_01|P0_SYNC _PG1_01|_AND_P|A1  2.067833848e-12
L_PG1_01|_AND_P|A2 _PG1_01|_AND_P|A1 _PG1_01|_AND_P|A2  4.135667696e-12
L_PG1_01|_AND_P|A3 _PG1_01|_AND_P|A3 _PG1_01|_AND_P|Q3  1.2e-12
L_PG1_01|_AND_P|B1 _PG1_01|P1_SYNC _PG1_01|_AND_P|B1  2.067833848e-12
L_PG1_01|_AND_P|B2 _PG1_01|_AND_P|B1 _PG1_01|_AND_P|B2  4.135667696e-12
L_PG1_01|_AND_P|B3 _PG1_01|_AND_P|B3 _PG1_01|_AND_P|Q3  1.2e-12
L_PG1_01|_AND_P|Q3 _PG1_01|_AND_P|Q3 _PG1_01|_AND_P|Q2  4.135667696e-12
L_PG1_01|_AND_P|Q2 _PG1_01|_AND_P|Q2 _PG1_01|_AND_P|Q1  4.135667696e-12
L_PG1_01|_AND_P|Q1 _PG1_01|_AND_P|Q1 P1_1_TX  2.067833848e-12
L_PG2_01|P|1 IP2_0_TO2 _PG2_01|P|A1  2.067833848e-12
L_PG2_01|P|2 _PG2_01|P|A1 _PG2_01|P|A2  4.135667696e-12
L_PG2_01|P|3 _PG2_01|P|A3 _PG2_01|P|A4  8.271335392e-12
L_PG2_01|P|T T13 _PG2_01|P|T1  2.067833848e-12
L_PG2_01|P|4 _PG2_01|P|T1 _PG2_01|P|T2  4.135667696e-12
L_PG2_01|P|5 _PG2_01|P|A4 _PG2_01|P|Q1  4.135667696e-12
L_PG2_01|P|6 _PG2_01|P|Q1 P2_1_TX  2.067833848e-12
L_PG2_01|G|1 IG2_0_TO2 _PG2_01|G|A1  2.067833848e-12
L_PG2_01|G|2 _PG2_01|G|A1 _PG2_01|G|A2  4.135667696e-12
L_PG2_01|G|3 _PG2_01|G|A3 _PG2_01|G|A4  8.271335392e-12
L_PG2_01|G|T T13 _PG2_01|G|T1  2.067833848e-12
L_PG2_01|G|4 _PG2_01|G|T1 _PG2_01|G|T2  4.135667696e-12
L_PG2_01|G|5 _PG2_01|G|A4 _PG2_01|G|Q1  4.135667696e-12
L_PG2_01|G|6 _PG2_01|G|Q1 G2_1_TX  2.067833848e-12
L_PG3_01|_SPL_G1|1 IG3_0_TO3 _PG3_01|_SPL_G1|D1  2e-12
L_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|D2  4.135667696e-12
L_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_G1|5 _PG3_01|_SPL_G1|QA1 _PG3_01|G1_COPY_1  2e-12
L_PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|QB1 _PG3_01|G1_COPY_2  2e-12
L_PG3_01|_SPL_P1|1 IP3_0_TO3 _PG3_01|_SPL_P1|D1  2e-12
L_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|D2  4.135667696e-12
L_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_P1|5 _PG3_01|_SPL_P1|QA1 _PG3_01|P1_COPY_1  2e-12
L_PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|QB1 _PG3_01|P1_COPY_2  2e-12
L_PG3_01|_PG|A1 _PG3_01|P1_COPY_1 _PG3_01|_PG|A1  2.067833848e-12
L_PG3_01|_PG|A2 _PG3_01|_PG|A1 _PG3_01|_PG|A2  4.135667696e-12
L_PG3_01|_PG|A3 _PG3_01|_PG|A3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|B1 _PG3_01|G1_COPY_1 _PG3_01|_PG|B1  2.067833848e-12
L_PG3_01|_PG|B2 _PG3_01|_PG|B1 _PG3_01|_PG|B2  4.135667696e-12
L_PG3_01|_PG|B3 _PG3_01|_PG|B3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|Q3 _PG3_01|_PG|Q3 _PG3_01|_PG|Q2  4.135667696e-12
L_PG3_01|_PG|Q2 _PG3_01|_PG|Q2 _PG3_01|_PG|Q1  4.135667696e-12
L_PG3_01|_PG|Q1 _PG3_01|_PG|Q1 _PG3_01|PG  2.067833848e-12
L_PG3_01|_GG|A1 IG2_0_TO3 _PG3_01|_GG|A1  2.067833848e-12
L_PG3_01|_GG|A2 _PG3_01|_GG|A1 _PG3_01|_GG|A2  4.135667696e-12
L_PG3_01|_GG|A3 _PG3_01|_GG|A3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|B1 _PG3_01|G1_COPY_2 _PG3_01|_GG|B1  2.067833848e-12
L_PG3_01|_GG|B2 _PG3_01|_GG|B1 _PG3_01|_GG|B2  4.135667696e-12
L_PG3_01|_GG|B3 _PG3_01|_GG|B3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|Q3 _PG3_01|_GG|Q3 _PG3_01|_GG|Q2  4.135667696e-12
L_PG3_01|_GG|Q2 _PG3_01|_GG|Q2 _PG3_01|_GG|Q1  4.135667696e-12
L_PG3_01|_GG|Q1 _PG3_01|_GG|Q1 _PG3_01|GG  2.067833848e-12
L_PG3_01|_DFF_P0|1 IP2_0_TO3 _PG3_01|_DFF_P0|A1  2.067833848e-12
L_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|A2  4.135667696e-12
L_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|A4  8.271335392e-12
L_PG3_01|_DFF_P0|T T14 _PG3_01|_DFF_P0|T1  2.067833848e-12
L_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T2  4.135667696e-12
L_PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|Q1  4.135667696e-12
L_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|Q1 _PG3_01|P0_SYNC  2.067833848e-12
L_PG3_01|_DFF_P1|1 _PG3_01|P1_COPY_2 _PG3_01|_DFF_P1|A1  2.067833848e-12
L_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|A2  4.135667696e-12
L_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|A4  8.271335392e-12
L_PG3_01|_DFF_P1|T T14 _PG3_01|_DFF_P1|T1  2.067833848e-12
L_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T2  4.135667696e-12
L_PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|Q1  4.135667696e-12
L_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|Q1 _PG3_01|P1_SYNC  2.067833848e-12
L_PG3_01|_DFF_PG|1 _PG3_01|PG _PG3_01|_DFF_PG|A1  2.067833848e-12
L_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|A2  4.135667696e-12
L_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|A4  8.271335392e-12
L_PG3_01|_DFF_PG|T T14 _PG3_01|_DFF_PG|T1  2.067833848e-12
L_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T2  4.135667696e-12
L_PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|Q1  4.135667696e-12
L_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|Q1 _PG3_01|PG_SYNC  2.067833848e-12
L_PG3_01|_DFF_GG|1 _PG3_01|GG _PG3_01|_DFF_GG|A1  2.067833848e-12
L_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|A2  4.135667696e-12
L_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|A4  8.271335392e-12
L_PG3_01|_DFF_GG|T T14 _PG3_01|_DFF_GG|T1  2.067833848e-12
L_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T2  4.135667696e-12
L_PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|Q1  4.135667696e-12
L_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|Q1 _PG3_01|GG_SYNC  2.067833848e-12
L_PG3_01|_AND_G|A1 _PG3_01|PG_SYNC _PG3_01|_AND_G|A1  2.067833848e-12
L_PG3_01|_AND_G|A2 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A2  4.135667696e-12
L_PG3_01|_AND_G|A3 _PG3_01|_AND_G|A3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|B1 _PG3_01|GG_SYNC _PG3_01|_AND_G|B1  2.067833848e-12
L_PG3_01|_AND_G|B2 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B2  4.135667696e-12
L_PG3_01|_AND_G|B3 _PG3_01|_AND_G|B3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q2  4.135667696e-12
L_PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q1  4.135667696e-12
L_PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1 G3_1_TX  2.067833848e-12
L_PG3_01|_AND_P|A1 _PG3_01|P0_SYNC _PG3_01|_AND_P|A1  2.067833848e-12
L_PG3_01|_AND_P|A2 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A2  4.135667696e-12
L_PG3_01|_AND_P|A3 _PG3_01|_AND_P|A3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|B1 _PG3_01|P1_SYNC _PG3_01|_AND_P|B1  2.067833848e-12
L_PG3_01|_AND_P|B2 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B2  4.135667696e-12
L_PG3_01|_AND_P|B3 _PG3_01|_AND_P|B3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q2  4.135667696e-12
L_PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q1  4.135667696e-12
L_PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1 P3_1_TX  2.067833848e-12
L_IP3_OUT|I_1|B _IP3_OUT|A1 _IP3_OUT|I_1|MID  2e-12
I_IP3_OUT|I_1|B 0 _IP3_OUT|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP3_OUT|I_3|B _IP3_OUT|A3 _IP3_OUT|I_3|MID  2e-12
I_IP3_OUT|I_3|B 0 _IP3_OUT|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP3_OUT|I_T|B _IP3_OUT|T1 _IP3_OUT|I_T|MID  2e-12
I_IP3_OUT|I_T|B 0 _IP3_OUT|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP3_OUT|I_6|B _IP3_OUT|Q1 _IP3_OUT|I_6|MID  2e-12
I_IP3_OUT|I_6|B 0 _IP3_OUT|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP3_OUT|1|1 _IP3_OUT|A1 _IP3_OUT|1|MID_SERIES JJMIT AREA=2.5
L_IP3_OUT|1|P _IP3_OUT|1|MID_SERIES 0  2e-13
R_IP3_OUT|1|B _IP3_OUT|A1 _IP3_OUT|1|MID_SHUNT  2.7439617672
L_IP3_OUT|1|RB _IP3_OUT|1|MID_SHUNT 0  1.550338398468e-12
B_IP3_OUT|23|1 _IP3_OUT|A2 _IP3_OUT|A3 JJMIT AREA=1.7857142857142858
R_IP3_OUT|23|B _IP3_OUT|A2 _IP3_OUT|23|MID_SHUNT  3.84154647408
L_IP3_OUT|23|RB _IP3_OUT|23|MID_SHUNT _IP3_OUT|A3  2.1704737578552e-12
B_IP3_OUT|3|1 _IP3_OUT|A3 _IP3_OUT|3|MID_SERIES JJMIT AREA=2.5
L_IP3_OUT|3|P _IP3_OUT|3|MID_SERIES 0  2e-13
R_IP3_OUT|3|B _IP3_OUT|A3 _IP3_OUT|3|MID_SHUNT  2.7439617672
L_IP3_OUT|3|RB _IP3_OUT|3|MID_SHUNT 0  1.550338398468e-12
B_IP3_OUT|4|1 _IP3_OUT|A4 _IP3_OUT|4|MID_SERIES JJMIT AREA=2.5
L_IP3_OUT|4|P _IP3_OUT|4|MID_SERIES 0  2e-13
R_IP3_OUT|4|B _IP3_OUT|A4 _IP3_OUT|4|MID_SHUNT  2.7439617672
L_IP3_OUT|4|RB _IP3_OUT|4|MID_SHUNT 0  1.550338398468e-12
B_IP3_OUT|T|1 _IP3_OUT|T1 _IP3_OUT|T|MID_SERIES JJMIT AREA=2.5
L_IP3_OUT|T|P _IP3_OUT|T|MID_SERIES 0  2e-13
R_IP3_OUT|T|B _IP3_OUT|T1 _IP3_OUT|T|MID_SHUNT  2.7439617672
L_IP3_OUT|T|RB _IP3_OUT|T|MID_SHUNT 0  1.550338398468e-12
B_IP3_OUT|45|1 _IP3_OUT|T2 _IP3_OUT|A4 JJMIT AREA=1.7857142857142858
R_IP3_OUT|45|B _IP3_OUT|T2 _IP3_OUT|45|MID_SHUNT  3.84154647408
L_IP3_OUT|45|RB _IP3_OUT|45|MID_SHUNT _IP3_OUT|A4  2.1704737578552e-12
B_IP3_OUT|6|1 _IP3_OUT|Q1 _IP3_OUT|6|MID_SERIES JJMIT AREA=2.5
L_IP3_OUT|6|P _IP3_OUT|6|MID_SERIES 0  2e-13
R_IP3_OUT|6|B _IP3_OUT|Q1 _IP3_OUT|6|MID_SHUNT  2.7439617672
L_IP3_OUT|6|RB _IP3_OUT|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_01|P|1 IP4_0_TO4 _PG4_01|P|A1  2.067833848e-12
L_PG4_01|P|2 _PG4_01|P|A1 _PG4_01|P|A2  4.135667696e-12
L_PG4_01|P|3 _PG4_01|P|A3 _PG4_01|P|A4  8.271335392e-12
L_PG4_01|P|T T16 _PG4_01|P|T1  2.067833848e-12
L_PG4_01|P|4 _PG4_01|P|T1 _PG4_01|P|T2  4.135667696e-12
L_PG4_01|P|5 _PG4_01|P|A4 _PG4_01|P|Q1  4.135667696e-12
L_PG4_01|P|6 _PG4_01|P|Q1 P4_1_TX  2.067833848e-12
L_PG4_01|G|1 IG4_0_TO4 _PG4_01|G|A1  2.067833848e-12
L_PG4_01|G|2 _PG4_01|G|A1 _PG4_01|G|A2  4.135667696e-12
L_PG4_01|G|3 _PG4_01|G|A3 _PG4_01|G|A4  8.271335392e-12
L_PG4_01|G|T T16 _PG4_01|G|T1  2.067833848e-12
L_PG4_01|G|4 _PG4_01|G|T1 _PG4_01|G|T2  4.135667696e-12
L_PG4_01|G|5 _PG4_01|G|A4 _PG4_01|G|Q1  4.135667696e-12
L_PG4_01|G|6 _PG4_01|G|Q1 G4_1_TX  2.067833848e-12
L_PG5_01|_SPL_G1|1 IG5_0_TO5 _PG5_01|_SPL_G1|D1  2e-12
L_PG5_01|_SPL_G1|2 _PG5_01|_SPL_G1|D1 _PG5_01|_SPL_G1|D2  4.135667696e-12
L_PG5_01|_SPL_G1|3 _PG5_01|_SPL_G1|D2 _PG5_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG5_01|_SPL_G1|4 _PG5_01|_SPL_G1|JCT _PG5_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG5_01|_SPL_G1|5 _PG5_01|_SPL_G1|QA1 _PG5_01|G1_COPY_1  2e-12
L_PG5_01|_SPL_G1|6 _PG5_01|_SPL_G1|JCT _PG5_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG5_01|_SPL_G1|7 _PG5_01|_SPL_G1|QB1 _PG5_01|G1_COPY_2  2e-12
L_PG5_01|_SPL_P1|1 IP5_0_TO5 _PG5_01|_SPL_P1|D1  2e-12
L_PG5_01|_SPL_P1|2 _PG5_01|_SPL_P1|D1 _PG5_01|_SPL_P1|D2  4.135667696e-12
L_PG5_01|_SPL_P1|3 _PG5_01|_SPL_P1|D2 _PG5_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG5_01|_SPL_P1|4 _PG5_01|_SPL_P1|JCT _PG5_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG5_01|_SPL_P1|5 _PG5_01|_SPL_P1|QA1 _PG5_01|P1_COPY_1  2e-12
L_PG5_01|_SPL_P1|6 _PG5_01|_SPL_P1|JCT _PG5_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG5_01|_SPL_P1|7 _PG5_01|_SPL_P1|QB1 _PG5_01|P1_COPY_2  2e-12
L_PG5_01|_PG|A1 _PG5_01|P1_COPY_1 _PG5_01|_PG|A1  2.067833848e-12
L_PG5_01|_PG|A2 _PG5_01|_PG|A1 _PG5_01|_PG|A2  4.135667696e-12
L_PG5_01|_PG|A3 _PG5_01|_PG|A3 _PG5_01|_PG|Q3  1.2e-12
L_PG5_01|_PG|B1 _PG5_01|G1_COPY_1 _PG5_01|_PG|B1  2.067833848e-12
L_PG5_01|_PG|B2 _PG5_01|_PG|B1 _PG5_01|_PG|B2  4.135667696e-12
L_PG5_01|_PG|B3 _PG5_01|_PG|B3 _PG5_01|_PG|Q3  1.2e-12
L_PG5_01|_PG|Q3 _PG5_01|_PG|Q3 _PG5_01|_PG|Q2  4.135667696e-12
L_PG5_01|_PG|Q2 _PG5_01|_PG|Q2 _PG5_01|_PG|Q1  4.135667696e-12
L_PG5_01|_PG|Q1 _PG5_01|_PG|Q1 _PG5_01|PG  2.067833848e-12
L_PG5_01|_GG|A1 IG4_0_TO5 _PG5_01|_GG|A1  2.067833848e-12
L_PG5_01|_GG|A2 _PG5_01|_GG|A1 _PG5_01|_GG|A2  4.135667696e-12
L_PG5_01|_GG|A3 _PG5_01|_GG|A3 _PG5_01|_GG|Q3  1.2e-12
L_PG5_01|_GG|B1 _PG5_01|G1_COPY_2 _PG5_01|_GG|B1  2.067833848e-12
L_PG5_01|_GG|B2 _PG5_01|_GG|B1 _PG5_01|_GG|B2  4.135667696e-12
L_PG5_01|_GG|B3 _PG5_01|_GG|B3 _PG5_01|_GG|Q3  1.2e-12
L_PG5_01|_GG|Q3 _PG5_01|_GG|Q3 _PG5_01|_GG|Q2  4.135667696e-12
L_PG5_01|_GG|Q2 _PG5_01|_GG|Q2 _PG5_01|_GG|Q1  4.135667696e-12
L_PG5_01|_GG|Q1 _PG5_01|_GG|Q1 _PG5_01|GG  2.067833848e-12
L_PG5_01|_DFF_P0|1 IP4_0_TO5 _PG5_01|_DFF_P0|A1  2.067833848e-12
L_PG5_01|_DFF_P0|2 _PG5_01|_DFF_P0|A1 _PG5_01|_DFF_P0|A2  4.135667696e-12
L_PG5_01|_DFF_P0|3 _PG5_01|_DFF_P0|A3 _PG5_01|_DFF_P0|A4  8.271335392e-12
L_PG5_01|_DFF_P0|T T17 _PG5_01|_DFF_P0|T1  2.067833848e-12
L_PG5_01|_DFF_P0|4 _PG5_01|_DFF_P0|T1 _PG5_01|_DFF_P0|T2  4.135667696e-12
L_PG5_01|_DFF_P0|5 _PG5_01|_DFF_P0|A4 _PG5_01|_DFF_P0|Q1  4.135667696e-12
L_PG5_01|_DFF_P0|6 _PG5_01|_DFF_P0|Q1 _PG5_01|P0_SYNC  2.067833848e-12
L_PG5_01|_DFF_P1|1 _PG5_01|P1_COPY_2 _PG5_01|_DFF_P1|A1  2.067833848e-12
L_PG5_01|_DFF_P1|2 _PG5_01|_DFF_P1|A1 _PG5_01|_DFF_P1|A2  4.135667696e-12
L_PG5_01|_DFF_P1|3 _PG5_01|_DFF_P1|A3 _PG5_01|_DFF_P1|A4  8.271335392e-12
L_PG5_01|_DFF_P1|T T17 _PG5_01|_DFF_P1|T1  2.067833848e-12
L_PG5_01|_DFF_P1|4 _PG5_01|_DFF_P1|T1 _PG5_01|_DFF_P1|T2  4.135667696e-12
L_PG5_01|_DFF_P1|5 _PG5_01|_DFF_P1|A4 _PG5_01|_DFF_P1|Q1  4.135667696e-12
L_PG5_01|_DFF_P1|6 _PG5_01|_DFF_P1|Q1 _PG5_01|P1_SYNC  2.067833848e-12
L_PG5_01|_DFF_PG|1 _PG5_01|PG _PG5_01|_DFF_PG|A1  2.067833848e-12
L_PG5_01|_DFF_PG|2 _PG5_01|_DFF_PG|A1 _PG5_01|_DFF_PG|A2  4.135667696e-12
L_PG5_01|_DFF_PG|3 _PG5_01|_DFF_PG|A3 _PG5_01|_DFF_PG|A4  8.271335392e-12
L_PG5_01|_DFF_PG|T T17 _PG5_01|_DFF_PG|T1  2.067833848e-12
L_PG5_01|_DFF_PG|4 _PG5_01|_DFF_PG|T1 _PG5_01|_DFF_PG|T2  4.135667696e-12
L_PG5_01|_DFF_PG|5 _PG5_01|_DFF_PG|A4 _PG5_01|_DFF_PG|Q1  4.135667696e-12
L_PG5_01|_DFF_PG|6 _PG5_01|_DFF_PG|Q1 _PG5_01|PG_SYNC  2.067833848e-12
L_PG5_01|_DFF_GG|1 _PG5_01|GG _PG5_01|_DFF_GG|A1  2.067833848e-12
L_PG5_01|_DFF_GG|2 _PG5_01|_DFF_GG|A1 _PG5_01|_DFF_GG|A2  4.135667696e-12
L_PG5_01|_DFF_GG|3 _PG5_01|_DFF_GG|A3 _PG5_01|_DFF_GG|A4  8.271335392e-12
L_PG5_01|_DFF_GG|T T17 _PG5_01|_DFF_GG|T1  2.067833848e-12
L_PG5_01|_DFF_GG|4 _PG5_01|_DFF_GG|T1 _PG5_01|_DFF_GG|T2  4.135667696e-12
L_PG5_01|_DFF_GG|5 _PG5_01|_DFF_GG|A4 _PG5_01|_DFF_GG|Q1  4.135667696e-12
L_PG5_01|_DFF_GG|6 _PG5_01|_DFF_GG|Q1 _PG5_01|GG_SYNC  2.067833848e-12
L_PG5_01|_AND_G|A1 _PG5_01|PG_SYNC _PG5_01|_AND_G|A1  2.067833848e-12
L_PG5_01|_AND_G|A2 _PG5_01|_AND_G|A1 _PG5_01|_AND_G|A2  4.135667696e-12
L_PG5_01|_AND_G|A3 _PG5_01|_AND_G|A3 _PG5_01|_AND_G|Q3  1.2e-12
L_PG5_01|_AND_G|B1 _PG5_01|GG_SYNC _PG5_01|_AND_G|B1  2.067833848e-12
L_PG5_01|_AND_G|B2 _PG5_01|_AND_G|B1 _PG5_01|_AND_G|B2  4.135667696e-12
L_PG5_01|_AND_G|B3 _PG5_01|_AND_G|B3 _PG5_01|_AND_G|Q3  1.2e-12
L_PG5_01|_AND_G|Q3 _PG5_01|_AND_G|Q3 _PG5_01|_AND_G|Q2  4.135667696e-12
L_PG5_01|_AND_G|Q2 _PG5_01|_AND_G|Q2 _PG5_01|_AND_G|Q1  4.135667696e-12
L_PG5_01|_AND_G|Q1 _PG5_01|_AND_G|Q1 G5_1_TX  2.067833848e-12
L_PG5_01|_AND_P|A1 _PG5_01|P0_SYNC _PG5_01|_AND_P|A1  2.067833848e-12
L_PG5_01|_AND_P|A2 _PG5_01|_AND_P|A1 _PG5_01|_AND_P|A2  4.135667696e-12
L_PG5_01|_AND_P|A3 _PG5_01|_AND_P|A3 _PG5_01|_AND_P|Q3  1.2e-12
L_PG5_01|_AND_P|B1 _PG5_01|P1_SYNC _PG5_01|_AND_P|B1  2.067833848e-12
L_PG5_01|_AND_P|B2 _PG5_01|_AND_P|B1 _PG5_01|_AND_P|B2  4.135667696e-12
L_PG5_01|_AND_P|B3 _PG5_01|_AND_P|B3 _PG5_01|_AND_P|Q3  1.2e-12
L_PG5_01|_AND_P|Q3 _PG5_01|_AND_P|Q3 _PG5_01|_AND_P|Q2  4.135667696e-12
L_PG5_01|_AND_P|Q2 _PG5_01|_AND_P|Q2 _PG5_01|_AND_P|Q1  4.135667696e-12
L_PG5_01|_AND_P|Q1 _PG5_01|_AND_P|Q1 P5_1_TX  2.067833848e-12
L_IP5_OUT|I_1|B _IP5_OUT|A1 _IP5_OUT|I_1|MID  2e-12
I_IP5_OUT|I_1|B 0 _IP5_OUT|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP5_OUT|I_3|B _IP5_OUT|A3 _IP5_OUT|I_3|MID  2e-12
I_IP5_OUT|I_3|B 0 _IP5_OUT|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP5_OUT|I_T|B _IP5_OUT|T1 _IP5_OUT|I_T|MID  2e-12
I_IP5_OUT|I_T|B 0 _IP5_OUT|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP5_OUT|I_6|B _IP5_OUT|Q1 _IP5_OUT|I_6|MID  2e-12
I_IP5_OUT|I_6|B 0 _IP5_OUT|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP5_OUT|1|1 _IP5_OUT|A1 _IP5_OUT|1|MID_SERIES JJMIT AREA=2.5
L_IP5_OUT|1|P _IP5_OUT|1|MID_SERIES 0  2e-13
R_IP5_OUT|1|B _IP5_OUT|A1 _IP5_OUT|1|MID_SHUNT  2.7439617672
L_IP5_OUT|1|RB _IP5_OUT|1|MID_SHUNT 0  1.550338398468e-12
B_IP5_OUT|23|1 _IP5_OUT|A2 _IP5_OUT|A3 JJMIT AREA=1.7857142857142858
R_IP5_OUT|23|B _IP5_OUT|A2 _IP5_OUT|23|MID_SHUNT  3.84154647408
L_IP5_OUT|23|RB _IP5_OUT|23|MID_SHUNT _IP5_OUT|A3  2.1704737578552e-12
B_IP5_OUT|3|1 _IP5_OUT|A3 _IP5_OUT|3|MID_SERIES JJMIT AREA=2.5
L_IP5_OUT|3|P _IP5_OUT|3|MID_SERIES 0  2e-13
R_IP5_OUT|3|B _IP5_OUT|A3 _IP5_OUT|3|MID_SHUNT  2.7439617672
L_IP5_OUT|3|RB _IP5_OUT|3|MID_SHUNT 0  1.550338398468e-12
B_IP5_OUT|4|1 _IP5_OUT|A4 _IP5_OUT|4|MID_SERIES JJMIT AREA=2.5
L_IP5_OUT|4|P _IP5_OUT|4|MID_SERIES 0  2e-13
R_IP5_OUT|4|B _IP5_OUT|A4 _IP5_OUT|4|MID_SHUNT  2.7439617672
L_IP5_OUT|4|RB _IP5_OUT|4|MID_SHUNT 0  1.550338398468e-12
B_IP5_OUT|T|1 _IP5_OUT|T1 _IP5_OUT|T|MID_SERIES JJMIT AREA=2.5
L_IP5_OUT|T|P _IP5_OUT|T|MID_SERIES 0  2e-13
R_IP5_OUT|T|B _IP5_OUT|T1 _IP5_OUT|T|MID_SHUNT  2.7439617672
L_IP5_OUT|T|RB _IP5_OUT|T|MID_SHUNT 0  1.550338398468e-12
B_IP5_OUT|45|1 _IP5_OUT|T2 _IP5_OUT|A4 JJMIT AREA=1.7857142857142858
R_IP5_OUT|45|B _IP5_OUT|T2 _IP5_OUT|45|MID_SHUNT  3.84154647408
L_IP5_OUT|45|RB _IP5_OUT|45|MID_SHUNT _IP5_OUT|A4  2.1704737578552e-12
B_IP5_OUT|6|1 _IP5_OUT|Q1 _IP5_OUT|6|MID_SERIES JJMIT AREA=2.5
L_IP5_OUT|6|P _IP5_OUT|6|MID_SERIES 0  2e-13
R_IP5_OUT|6|B _IP5_OUT|Q1 _IP5_OUT|6|MID_SHUNT  2.7439617672
L_IP5_OUT|6|RB _IP5_OUT|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_01|P|1 IP6_0_TO6 _PG6_01|P|A1  2.067833848e-12
L_PG6_01|P|2 _PG6_01|P|A1 _PG6_01|P|A2  4.135667696e-12
L_PG6_01|P|3 _PG6_01|P|A3 _PG6_01|P|A4  8.271335392e-12
L_PG6_01|P|T T19 _PG6_01|P|T1  2.067833848e-12
L_PG6_01|P|4 _PG6_01|P|T1 _PG6_01|P|T2  4.135667696e-12
L_PG6_01|P|5 _PG6_01|P|A4 _PG6_01|P|Q1  4.135667696e-12
L_PG6_01|P|6 _PG6_01|P|Q1 P6_1_TX  2.067833848e-12
L_PG6_01|G|1 IG6_0_TO6 _PG6_01|G|A1  2.067833848e-12
L_PG6_01|G|2 _PG6_01|G|A1 _PG6_01|G|A2  4.135667696e-12
L_PG6_01|G|3 _PG6_01|G|A3 _PG6_01|G|A4  8.271335392e-12
L_PG6_01|G|T T19 _PG6_01|G|T1  2.067833848e-12
L_PG6_01|G|4 _PG6_01|G|T1 _PG6_01|G|T2  4.135667696e-12
L_PG6_01|G|5 _PG6_01|G|A4 _PG6_01|G|Q1  4.135667696e-12
L_PG6_01|G|6 _PG6_01|G|Q1 G6_1_TX  2.067833848e-12
L_PG7_01|_SPL_G1|1 IG7_0_TO7 _PG7_01|_SPL_G1|D1  2e-12
L_PG7_01|_SPL_G1|2 _PG7_01|_SPL_G1|D1 _PG7_01|_SPL_G1|D2  4.135667696e-12
L_PG7_01|_SPL_G1|3 _PG7_01|_SPL_G1|D2 _PG7_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG7_01|_SPL_G1|4 _PG7_01|_SPL_G1|JCT _PG7_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG7_01|_SPL_G1|5 _PG7_01|_SPL_G1|QA1 _PG7_01|G1_COPY_1  2e-12
L_PG7_01|_SPL_G1|6 _PG7_01|_SPL_G1|JCT _PG7_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG7_01|_SPL_G1|7 _PG7_01|_SPL_G1|QB1 _PG7_01|G1_COPY_2  2e-12
L_PG7_01|_SPL_P1|1 IP7_0_TO7 _PG7_01|_SPL_P1|D1  2e-12
L_PG7_01|_SPL_P1|2 _PG7_01|_SPL_P1|D1 _PG7_01|_SPL_P1|D2  4.135667696e-12
L_PG7_01|_SPL_P1|3 _PG7_01|_SPL_P1|D2 _PG7_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG7_01|_SPL_P1|4 _PG7_01|_SPL_P1|JCT _PG7_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG7_01|_SPL_P1|5 _PG7_01|_SPL_P1|QA1 _PG7_01|P1_COPY_1  2e-12
L_PG7_01|_SPL_P1|6 _PG7_01|_SPL_P1|JCT _PG7_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG7_01|_SPL_P1|7 _PG7_01|_SPL_P1|QB1 _PG7_01|P1_COPY_2  2e-12
L_PG7_01|_PG|A1 _PG7_01|P1_COPY_1 _PG7_01|_PG|A1  2.067833848e-12
L_PG7_01|_PG|A2 _PG7_01|_PG|A1 _PG7_01|_PG|A2  4.135667696e-12
L_PG7_01|_PG|A3 _PG7_01|_PG|A3 _PG7_01|_PG|Q3  1.2e-12
L_PG7_01|_PG|B1 _PG7_01|G1_COPY_1 _PG7_01|_PG|B1  2.067833848e-12
L_PG7_01|_PG|B2 _PG7_01|_PG|B1 _PG7_01|_PG|B2  4.135667696e-12
L_PG7_01|_PG|B3 _PG7_01|_PG|B3 _PG7_01|_PG|Q3  1.2e-12
L_PG7_01|_PG|Q3 _PG7_01|_PG|Q3 _PG7_01|_PG|Q2  4.135667696e-12
L_PG7_01|_PG|Q2 _PG7_01|_PG|Q2 _PG7_01|_PG|Q1  4.135667696e-12
L_PG7_01|_PG|Q1 _PG7_01|_PG|Q1 _PG7_01|PG  2.067833848e-12
L_PG7_01|_GG|A1 IG6_0_TO7 _PG7_01|_GG|A1  2.067833848e-12
L_PG7_01|_GG|A2 _PG7_01|_GG|A1 _PG7_01|_GG|A2  4.135667696e-12
L_PG7_01|_GG|A3 _PG7_01|_GG|A3 _PG7_01|_GG|Q3  1.2e-12
L_PG7_01|_GG|B1 _PG7_01|G1_COPY_2 _PG7_01|_GG|B1  2.067833848e-12
L_PG7_01|_GG|B2 _PG7_01|_GG|B1 _PG7_01|_GG|B2  4.135667696e-12
L_PG7_01|_GG|B3 _PG7_01|_GG|B3 _PG7_01|_GG|Q3  1.2e-12
L_PG7_01|_GG|Q3 _PG7_01|_GG|Q3 _PG7_01|_GG|Q2  4.135667696e-12
L_PG7_01|_GG|Q2 _PG7_01|_GG|Q2 _PG7_01|_GG|Q1  4.135667696e-12
L_PG7_01|_GG|Q1 _PG7_01|_GG|Q1 _PG7_01|GG  2.067833848e-12
L_PG7_01|_DFF_P0|1 IP6_0_TO7 _PG7_01|_DFF_P0|A1  2.067833848e-12
L_PG7_01|_DFF_P0|2 _PG7_01|_DFF_P0|A1 _PG7_01|_DFF_P0|A2  4.135667696e-12
L_PG7_01|_DFF_P0|3 _PG7_01|_DFF_P0|A3 _PG7_01|_DFF_P0|A4  8.271335392e-12
L_PG7_01|_DFF_P0|T T1A _PG7_01|_DFF_P0|T1  2.067833848e-12
L_PG7_01|_DFF_P0|4 _PG7_01|_DFF_P0|T1 _PG7_01|_DFF_P0|T2  4.135667696e-12
L_PG7_01|_DFF_P0|5 _PG7_01|_DFF_P0|A4 _PG7_01|_DFF_P0|Q1  4.135667696e-12
L_PG7_01|_DFF_P0|6 _PG7_01|_DFF_P0|Q1 _PG7_01|P0_SYNC  2.067833848e-12
L_PG7_01|_DFF_P1|1 _PG7_01|P1_COPY_2 _PG7_01|_DFF_P1|A1  2.067833848e-12
L_PG7_01|_DFF_P1|2 _PG7_01|_DFF_P1|A1 _PG7_01|_DFF_P1|A2  4.135667696e-12
L_PG7_01|_DFF_P1|3 _PG7_01|_DFF_P1|A3 _PG7_01|_DFF_P1|A4  8.271335392e-12
L_PG7_01|_DFF_P1|T T1A _PG7_01|_DFF_P1|T1  2.067833848e-12
L_PG7_01|_DFF_P1|4 _PG7_01|_DFF_P1|T1 _PG7_01|_DFF_P1|T2  4.135667696e-12
L_PG7_01|_DFF_P1|5 _PG7_01|_DFF_P1|A4 _PG7_01|_DFF_P1|Q1  4.135667696e-12
L_PG7_01|_DFF_P1|6 _PG7_01|_DFF_P1|Q1 _PG7_01|P1_SYNC  2.067833848e-12
L_PG7_01|_DFF_PG|1 _PG7_01|PG _PG7_01|_DFF_PG|A1  2.067833848e-12
L_PG7_01|_DFF_PG|2 _PG7_01|_DFF_PG|A1 _PG7_01|_DFF_PG|A2  4.135667696e-12
L_PG7_01|_DFF_PG|3 _PG7_01|_DFF_PG|A3 _PG7_01|_DFF_PG|A4  8.271335392e-12
L_PG7_01|_DFF_PG|T T1A _PG7_01|_DFF_PG|T1  2.067833848e-12
L_PG7_01|_DFF_PG|4 _PG7_01|_DFF_PG|T1 _PG7_01|_DFF_PG|T2  4.135667696e-12
L_PG7_01|_DFF_PG|5 _PG7_01|_DFF_PG|A4 _PG7_01|_DFF_PG|Q1  4.135667696e-12
L_PG7_01|_DFF_PG|6 _PG7_01|_DFF_PG|Q1 _PG7_01|PG_SYNC  2.067833848e-12
L_PG7_01|_DFF_GG|1 _PG7_01|GG _PG7_01|_DFF_GG|A1  2.067833848e-12
L_PG7_01|_DFF_GG|2 _PG7_01|_DFF_GG|A1 _PG7_01|_DFF_GG|A2  4.135667696e-12
L_PG7_01|_DFF_GG|3 _PG7_01|_DFF_GG|A3 _PG7_01|_DFF_GG|A4  8.271335392e-12
L_PG7_01|_DFF_GG|T T1A _PG7_01|_DFF_GG|T1  2.067833848e-12
L_PG7_01|_DFF_GG|4 _PG7_01|_DFF_GG|T1 _PG7_01|_DFF_GG|T2  4.135667696e-12
L_PG7_01|_DFF_GG|5 _PG7_01|_DFF_GG|A4 _PG7_01|_DFF_GG|Q1  4.135667696e-12
L_PG7_01|_DFF_GG|6 _PG7_01|_DFF_GG|Q1 _PG7_01|GG_SYNC  2.067833848e-12
L_PG7_01|_AND_G|A1 _PG7_01|PG_SYNC _PG7_01|_AND_G|A1  2.067833848e-12
L_PG7_01|_AND_G|A2 _PG7_01|_AND_G|A1 _PG7_01|_AND_G|A2  4.135667696e-12
L_PG7_01|_AND_G|A3 _PG7_01|_AND_G|A3 _PG7_01|_AND_G|Q3  1.2e-12
L_PG7_01|_AND_G|B1 _PG7_01|GG_SYNC _PG7_01|_AND_G|B1  2.067833848e-12
L_PG7_01|_AND_G|B2 _PG7_01|_AND_G|B1 _PG7_01|_AND_G|B2  4.135667696e-12
L_PG7_01|_AND_G|B3 _PG7_01|_AND_G|B3 _PG7_01|_AND_G|Q3  1.2e-12
L_PG7_01|_AND_G|Q3 _PG7_01|_AND_G|Q3 _PG7_01|_AND_G|Q2  4.135667696e-12
L_PG7_01|_AND_G|Q2 _PG7_01|_AND_G|Q2 _PG7_01|_AND_G|Q1  4.135667696e-12
L_PG7_01|_AND_G|Q1 _PG7_01|_AND_G|Q1 G7_1_TX  2.067833848e-12
L_PG7_01|_AND_P|A1 _PG7_01|P0_SYNC _PG7_01|_AND_P|A1  2.067833848e-12
L_PG7_01|_AND_P|A2 _PG7_01|_AND_P|A1 _PG7_01|_AND_P|A2  4.135667696e-12
L_PG7_01|_AND_P|A3 _PG7_01|_AND_P|A3 _PG7_01|_AND_P|Q3  1.2e-12
L_PG7_01|_AND_P|B1 _PG7_01|P1_SYNC _PG7_01|_AND_P|B1  2.067833848e-12
L_PG7_01|_AND_P|B2 _PG7_01|_AND_P|B1 _PG7_01|_AND_P|B2  4.135667696e-12
L_PG7_01|_AND_P|B3 _PG7_01|_AND_P|B3 _PG7_01|_AND_P|Q3  1.2e-12
L_PG7_01|_AND_P|Q3 _PG7_01|_AND_P|Q3 _PG7_01|_AND_P|Q2  4.135667696e-12
L_PG7_01|_AND_P|Q2 _PG7_01|_AND_P|Q2 _PG7_01|_AND_P|Q1  4.135667696e-12
L_PG7_01|_AND_P|Q1 _PG7_01|_AND_P|Q1 P7_1_TX  2.067833848e-12
L_IP7_OUT|I_1|B _IP7_OUT|A1 _IP7_OUT|I_1|MID  2e-12
I_IP7_OUT|I_1|B 0 _IP7_OUT|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP7_OUT|I_3|B _IP7_OUT|A3 _IP7_OUT|I_3|MID  2e-12
I_IP7_OUT|I_3|B 0 _IP7_OUT|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP7_OUT|I_T|B _IP7_OUT|T1 _IP7_OUT|I_T|MID  2e-12
I_IP7_OUT|I_T|B 0 _IP7_OUT|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP7_OUT|I_6|B _IP7_OUT|Q1 _IP7_OUT|I_6|MID  2e-12
I_IP7_OUT|I_6|B 0 _IP7_OUT|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP7_OUT|1|1 _IP7_OUT|A1 _IP7_OUT|1|MID_SERIES JJMIT AREA=2.5
L_IP7_OUT|1|P _IP7_OUT|1|MID_SERIES 0  2e-13
R_IP7_OUT|1|B _IP7_OUT|A1 _IP7_OUT|1|MID_SHUNT  2.7439617672
L_IP7_OUT|1|RB _IP7_OUT|1|MID_SHUNT 0  1.550338398468e-12
B_IP7_OUT|23|1 _IP7_OUT|A2 _IP7_OUT|A3 JJMIT AREA=1.7857142857142858
R_IP7_OUT|23|B _IP7_OUT|A2 _IP7_OUT|23|MID_SHUNT  3.84154647408
L_IP7_OUT|23|RB _IP7_OUT|23|MID_SHUNT _IP7_OUT|A3  2.1704737578552e-12
B_IP7_OUT|3|1 _IP7_OUT|A3 _IP7_OUT|3|MID_SERIES JJMIT AREA=2.5
L_IP7_OUT|3|P _IP7_OUT|3|MID_SERIES 0  2e-13
R_IP7_OUT|3|B _IP7_OUT|A3 _IP7_OUT|3|MID_SHUNT  2.7439617672
L_IP7_OUT|3|RB _IP7_OUT|3|MID_SHUNT 0  1.550338398468e-12
B_IP7_OUT|4|1 _IP7_OUT|A4 _IP7_OUT|4|MID_SERIES JJMIT AREA=2.5
L_IP7_OUT|4|P _IP7_OUT|4|MID_SERIES 0  2e-13
R_IP7_OUT|4|B _IP7_OUT|A4 _IP7_OUT|4|MID_SHUNT  2.7439617672
L_IP7_OUT|4|RB _IP7_OUT|4|MID_SHUNT 0  1.550338398468e-12
B_IP7_OUT|T|1 _IP7_OUT|T1 _IP7_OUT|T|MID_SERIES JJMIT AREA=2.5
L_IP7_OUT|T|P _IP7_OUT|T|MID_SERIES 0  2e-13
R_IP7_OUT|T|B _IP7_OUT|T1 _IP7_OUT|T|MID_SHUNT  2.7439617672
L_IP7_OUT|T|RB _IP7_OUT|T|MID_SHUNT 0  1.550338398468e-12
B_IP7_OUT|45|1 _IP7_OUT|T2 _IP7_OUT|A4 JJMIT AREA=1.7857142857142858
R_IP7_OUT|45|B _IP7_OUT|T2 _IP7_OUT|45|MID_SHUNT  3.84154647408
L_IP7_OUT|45|RB _IP7_OUT|45|MID_SHUNT _IP7_OUT|A4  2.1704737578552e-12
B_IP7_OUT|6|1 _IP7_OUT|Q1 _IP7_OUT|6|MID_SERIES JJMIT AREA=2.5
L_IP7_OUT|6|P _IP7_OUT|6|MID_SERIES 0  2e-13
R_IP7_OUT|6|B _IP7_OUT|Q1 _IP7_OUT|6|MID_SHUNT  2.7439617672
L_IP7_OUT|6|RB _IP7_OUT|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_S0_1|_TX|1 _PTL_S0_1|_TX|1 _PTL_S0_1|_TX|2 JJMIT AREA=2.5
B_PTL_S0_1|_TX|2 _PTL_S0_1|_TX|4 _PTL_S0_1|_TX|5 JJMIT AREA=2.5
I_PTL_S0_1|_TX|B1 0 _PTL_S0_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S0_1|_TX|B2 0 _PTL_S0_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S0_1|_TX|B1 _PTL_S0_1|_TX|1 _PTL_S0_1|_TX|3  1.684e-12
L_PTL_S0_1|_TX|B2 _PTL_S0_1|_TX|4 _PTL_S0_1|_TX|6  3.596e-12
L_PTL_S0_1|_TX|1 S0_1_TX _PTL_S0_1|_TX|1  2.063e-12
L_PTL_S0_1|_TX|2 _PTL_S0_1|_TX|1 _PTL_S0_1|_TX|4  4.123e-12
L_PTL_S0_1|_TX|3 _PTL_S0_1|_TX|4 _PTL_S0_1|_TX|7  2.193e-12
R_PTL_S0_1|_TX|D _PTL_S0_1|_TX|7 _PTL_S0_1|A_PTL  1.36
L_PTL_S0_1|_TX|P1 _PTL_S0_1|_TX|2 0  5.254e-13
L_PTL_S0_1|_TX|P2 _PTL_S0_1|_TX|5 0  5.141e-13
R_PTL_S0_1|_TX|B1 _PTL_S0_1|_TX|1 _PTL_S0_1|_TX|101  2.7439617672
R_PTL_S0_1|_TX|B2 _PTL_S0_1|_TX|4 _PTL_S0_1|_TX|104  2.7439617672
L_PTL_S0_1|_TX|RB1 _PTL_S0_1|_TX|101 0  1.550338398468e-12
L_PTL_S0_1|_TX|RB2 _PTL_S0_1|_TX|104 0  1.550338398468e-12
B_PTL_S0_1|_RX|1 _PTL_S0_1|_RX|1 _PTL_S0_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S0_1|_RX|2 _PTL_S0_1|_RX|4 _PTL_S0_1|_RX|5 JJMIT AREA=2.0
B_PTL_S0_1|_RX|3 _PTL_S0_1|_RX|7 _PTL_S0_1|_RX|8 JJMIT AREA=2.5
I_PTL_S0_1|_RX|B1 0 _PTL_S0_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S0_1|_RX|B1 _PTL_S0_1|_RX|1 _PTL_S0_1|_RX|3  2.777e-12
I_PTL_S0_1|_RX|B2 0 _PTL_S0_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S0_1|_RX|B2 _PTL_S0_1|_RX|4 _PTL_S0_1|_RX|6  2.685e-12
I_PTL_S0_1|_RX|B3 0 _PTL_S0_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S0_1|_RX|B3 _PTL_S0_1|_RX|7 _PTL_S0_1|_RX|9  2.764e-12
L_PTL_S0_1|_RX|1 _PTL_S0_1|A_PTL _PTL_S0_1|_RX|1  1.346e-12
L_PTL_S0_1|_RX|2 _PTL_S0_1|_RX|1 _PTL_S0_1|_RX|4  6.348e-12
L_PTL_S0_1|_RX|3 _PTL_S0_1|_RX|4 _PTL_S0_1|_RX|7  5.197e-12
L_PTL_S0_1|_RX|4 _PTL_S0_1|_RX|7 S0_1  2.058e-12
L_PTL_S0_1|_RX|P1 _PTL_S0_1|_RX|2 0  4.795e-13
L_PTL_S0_1|_RX|P2 _PTL_S0_1|_RX|5 0  5.431e-13
L_PTL_S0_1|_RX|P3 _PTL_S0_1|_RX|8 0  5.339e-13
R_PTL_S0_1|_RX|B1 _PTL_S0_1|_RX|1 _PTL_S0_1|_RX|101  4.225701121488
R_PTL_S0_1|_RX|B2 _PTL_S0_1|_RX|4 _PTL_S0_1|_RX|104  3.429952209
R_PTL_S0_1|_RX|B3 _PTL_S0_1|_RX|7 _PTL_S0_1|_RX|107  2.7439617672
L_PTL_S0_1|_RX|RB1 _PTL_S0_1|_RX|101 0  2.38752113364072e-12
L_PTL_S0_1|_RX|RB2 _PTL_S0_1|_RX|104 0  1.937922998085e-12
L_PTL_S0_1|_RX|RB3 _PTL_S0_1|_RX|107 0  1.550338398468e-12
B_PTL_S1_1|_TX|1 _PTL_S1_1|_TX|1 _PTL_S1_1|_TX|2 JJMIT AREA=2.5
B_PTL_S1_1|_TX|2 _PTL_S1_1|_TX|4 _PTL_S1_1|_TX|5 JJMIT AREA=2.5
I_PTL_S1_1|_TX|B1 0 _PTL_S1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S1_1|_TX|B2 0 _PTL_S1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S1_1|_TX|B1 _PTL_S1_1|_TX|1 _PTL_S1_1|_TX|3  1.684e-12
L_PTL_S1_1|_TX|B2 _PTL_S1_1|_TX|4 _PTL_S1_1|_TX|6  3.596e-12
L_PTL_S1_1|_TX|1 S1_1_TX _PTL_S1_1|_TX|1  2.063e-12
L_PTL_S1_1|_TX|2 _PTL_S1_1|_TX|1 _PTL_S1_1|_TX|4  4.123e-12
L_PTL_S1_1|_TX|3 _PTL_S1_1|_TX|4 _PTL_S1_1|_TX|7  2.193e-12
R_PTL_S1_1|_TX|D _PTL_S1_1|_TX|7 _PTL_S1_1|A_PTL  1.36
L_PTL_S1_1|_TX|P1 _PTL_S1_1|_TX|2 0  5.254e-13
L_PTL_S1_1|_TX|P2 _PTL_S1_1|_TX|5 0  5.141e-13
R_PTL_S1_1|_TX|B1 _PTL_S1_1|_TX|1 _PTL_S1_1|_TX|101  2.7439617672
R_PTL_S1_1|_TX|B2 _PTL_S1_1|_TX|4 _PTL_S1_1|_TX|104  2.7439617672
L_PTL_S1_1|_TX|RB1 _PTL_S1_1|_TX|101 0  1.550338398468e-12
L_PTL_S1_1|_TX|RB2 _PTL_S1_1|_TX|104 0  1.550338398468e-12
B_PTL_S1_1|_RX|1 _PTL_S1_1|_RX|1 _PTL_S1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S1_1|_RX|2 _PTL_S1_1|_RX|4 _PTL_S1_1|_RX|5 JJMIT AREA=2.0
B_PTL_S1_1|_RX|3 _PTL_S1_1|_RX|7 _PTL_S1_1|_RX|8 JJMIT AREA=2.5
I_PTL_S1_1|_RX|B1 0 _PTL_S1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S1_1|_RX|B1 _PTL_S1_1|_RX|1 _PTL_S1_1|_RX|3  2.777e-12
I_PTL_S1_1|_RX|B2 0 _PTL_S1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S1_1|_RX|B2 _PTL_S1_1|_RX|4 _PTL_S1_1|_RX|6  2.685e-12
I_PTL_S1_1|_RX|B3 0 _PTL_S1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S1_1|_RX|B3 _PTL_S1_1|_RX|7 _PTL_S1_1|_RX|9  2.764e-12
L_PTL_S1_1|_RX|1 _PTL_S1_1|A_PTL _PTL_S1_1|_RX|1  1.346e-12
L_PTL_S1_1|_RX|2 _PTL_S1_1|_RX|1 _PTL_S1_1|_RX|4  6.348e-12
L_PTL_S1_1|_RX|3 _PTL_S1_1|_RX|4 _PTL_S1_1|_RX|7  5.197e-12
L_PTL_S1_1|_RX|4 _PTL_S1_1|_RX|7 S1_1  2.058e-12
L_PTL_S1_1|_RX|P1 _PTL_S1_1|_RX|2 0  4.795e-13
L_PTL_S1_1|_RX|P2 _PTL_S1_1|_RX|5 0  5.431e-13
L_PTL_S1_1|_RX|P3 _PTL_S1_1|_RX|8 0  5.339e-13
R_PTL_S1_1|_RX|B1 _PTL_S1_1|_RX|1 _PTL_S1_1|_RX|101  4.225701121488
R_PTL_S1_1|_RX|B2 _PTL_S1_1|_RX|4 _PTL_S1_1|_RX|104  3.429952209
R_PTL_S1_1|_RX|B3 _PTL_S1_1|_RX|7 _PTL_S1_1|_RX|107  2.7439617672
L_PTL_S1_1|_RX|RB1 _PTL_S1_1|_RX|101 0  2.38752113364072e-12
L_PTL_S1_1|_RX|RB2 _PTL_S1_1|_RX|104 0  1.937922998085e-12
L_PTL_S1_1|_RX|RB3 _PTL_S1_1|_RX|107 0  1.550338398468e-12
B_PTL_P1_1|_TX|1 _PTL_P1_1|_TX|1 _PTL_P1_1|_TX|2 JJMIT AREA=2.5
B_PTL_P1_1|_TX|2 _PTL_P1_1|_TX|4 _PTL_P1_1|_TX|5 JJMIT AREA=2.5
I_PTL_P1_1|_TX|B1 0 _PTL_P1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P1_1|_TX|B2 0 _PTL_P1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P1_1|_TX|B1 _PTL_P1_1|_TX|1 _PTL_P1_1|_TX|3  1.684e-12
L_PTL_P1_1|_TX|B2 _PTL_P1_1|_TX|4 _PTL_P1_1|_TX|6  3.596e-12
L_PTL_P1_1|_TX|1 P1_1_TX _PTL_P1_1|_TX|1  2.063e-12
L_PTL_P1_1|_TX|2 _PTL_P1_1|_TX|1 _PTL_P1_1|_TX|4  4.123e-12
L_PTL_P1_1|_TX|3 _PTL_P1_1|_TX|4 _PTL_P1_1|_TX|7  2.193e-12
R_PTL_P1_1|_TX|D _PTL_P1_1|_TX|7 _PTL_P1_1|A_PTL  1.36
L_PTL_P1_1|_TX|P1 _PTL_P1_1|_TX|2 0  5.254e-13
L_PTL_P1_1|_TX|P2 _PTL_P1_1|_TX|5 0  5.141e-13
R_PTL_P1_1|_TX|B1 _PTL_P1_1|_TX|1 _PTL_P1_1|_TX|101  2.7439617672
R_PTL_P1_1|_TX|B2 _PTL_P1_1|_TX|4 _PTL_P1_1|_TX|104  2.7439617672
L_PTL_P1_1|_TX|RB1 _PTL_P1_1|_TX|101 0  1.550338398468e-12
L_PTL_P1_1|_TX|RB2 _PTL_P1_1|_TX|104 0  1.550338398468e-12
B_PTL_P1_1|_RX|1 _PTL_P1_1|_RX|1 _PTL_P1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P1_1|_RX|2 _PTL_P1_1|_RX|4 _PTL_P1_1|_RX|5 JJMIT AREA=2.0
B_PTL_P1_1|_RX|3 _PTL_P1_1|_RX|7 _PTL_P1_1|_RX|8 JJMIT AREA=2.5
I_PTL_P1_1|_RX|B1 0 _PTL_P1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P1_1|_RX|B1 _PTL_P1_1|_RX|1 _PTL_P1_1|_RX|3  2.777e-12
I_PTL_P1_1|_RX|B2 0 _PTL_P1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P1_1|_RX|B2 _PTL_P1_1|_RX|4 _PTL_P1_1|_RX|6  2.685e-12
I_PTL_P1_1|_RX|B3 0 _PTL_P1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P1_1|_RX|B3 _PTL_P1_1|_RX|7 _PTL_P1_1|_RX|9  2.764e-12
L_PTL_P1_1|_RX|1 _PTL_P1_1|A_PTL _PTL_P1_1|_RX|1  1.346e-12
L_PTL_P1_1|_RX|2 _PTL_P1_1|_RX|1 _PTL_P1_1|_RX|4  6.348e-12
L_PTL_P1_1|_RX|3 _PTL_P1_1|_RX|4 _PTL_P1_1|_RX|7  5.197e-12
L_PTL_P1_1|_RX|4 _PTL_P1_1|_RX|7 _PTL_P1_1|D  2.058e-12
L_PTL_P1_1|_RX|P1 _PTL_P1_1|_RX|2 0  4.795e-13
L_PTL_P1_1|_RX|P2 _PTL_P1_1|_RX|5 0  5.431e-13
L_PTL_P1_1|_RX|P3 _PTL_P1_1|_RX|8 0  5.339e-13
R_PTL_P1_1|_RX|B1 _PTL_P1_1|_RX|1 _PTL_P1_1|_RX|101  4.225701121488
R_PTL_P1_1|_RX|B2 _PTL_P1_1|_RX|4 _PTL_P1_1|_RX|104  3.429952209
R_PTL_P1_1|_RX|B3 _PTL_P1_1|_RX|7 _PTL_P1_1|_RX|107  2.7439617672
L_PTL_P1_1|_RX|RB1 _PTL_P1_1|_RX|101 0  2.38752113364072e-12
L_PTL_P1_1|_RX|RB2 _PTL_P1_1|_RX|104 0  1.937922998085e-12
L_PTL_P1_1|_RX|RB3 _PTL_P1_1|_RX|107 0  1.550338398468e-12
L_PTL_P1_1|_SPL|1 _PTL_P1_1|D _PTL_P1_1|_SPL|D1  2e-12
L_PTL_P1_1|_SPL|2 _PTL_P1_1|_SPL|D1 _PTL_P1_1|_SPL|D2  4.135667696e-12
L_PTL_P1_1|_SPL|3 _PTL_P1_1|_SPL|D2 _PTL_P1_1|_SPL|JCT  9.84682784761905e-13
L_PTL_P1_1|_SPL|4 _PTL_P1_1|_SPL|JCT _PTL_P1_1|_SPL|QA1  9.84682784761905e-13
L_PTL_P1_1|_SPL|5 _PTL_P1_1|_SPL|QA1 P1_1_TO2  2e-12
L_PTL_P1_1|_SPL|6 _PTL_P1_1|_SPL|JCT _PTL_P1_1|_SPL|QB1  9.84682784761905e-13
L_PTL_P1_1|_SPL|7 _PTL_P1_1|_SPL|QB1 P1_1_TO3  2e-12
B_PTL_G1_1|_TX|1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|2 JJMIT AREA=2.5
B_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|5 JJMIT AREA=2.5
I_PTL_G1_1|_TX|B1 0 _PTL_G1_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G1_1|_TX|B2 0 _PTL_G1_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|3  1.684e-12
L_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|6  3.596e-12
L_PTL_G1_1|_TX|1 G1_1_TX _PTL_G1_1|_TX|1  2.063e-12
L_PTL_G1_1|_TX|2 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|4  4.123e-12
L_PTL_G1_1|_TX|3 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|7  2.193e-12
R_PTL_G1_1|_TX|D _PTL_G1_1|_TX|7 _PTL_G1_1|A_PTL  1.36
L_PTL_G1_1|_TX|P1 _PTL_G1_1|_TX|2 0  5.254e-13
L_PTL_G1_1|_TX|P2 _PTL_G1_1|_TX|5 0  5.141e-13
R_PTL_G1_1|_TX|B1 _PTL_G1_1|_TX|1 _PTL_G1_1|_TX|101  2.7439617672
R_PTL_G1_1|_TX|B2 _PTL_G1_1|_TX|4 _PTL_G1_1|_TX|104  2.7439617672
L_PTL_G1_1|_TX|RB1 _PTL_G1_1|_TX|101 0  1.550338398468e-12
L_PTL_G1_1|_TX|RB2 _PTL_G1_1|_TX|104 0  1.550338398468e-12
B_PTL_G1_1|_RX|1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|5 JJMIT AREA=2.0
B_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|8 JJMIT AREA=2.5
I_PTL_G1_1|_RX|B1 0 _PTL_G1_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|3  2.777e-12
I_PTL_G1_1|_RX|B2 0 _PTL_G1_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|6  2.685e-12
I_PTL_G1_1|_RX|B3 0 _PTL_G1_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|9  2.764e-12
L_PTL_G1_1|_RX|1 _PTL_G1_1|A_PTL _PTL_G1_1|_RX|1  1.346e-12
L_PTL_G1_1|_RX|2 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|4  6.348e-12
L_PTL_G1_1|_RX|3 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7  5.197e-12
L_PTL_G1_1|_RX|4 _PTL_G1_1|_RX|7 _PTL_G1_1|D  2.058e-12
L_PTL_G1_1|_RX|P1 _PTL_G1_1|_RX|2 0  4.795e-13
L_PTL_G1_1|_RX|P2 _PTL_G1_1|_RX|5 0  5.431e-13
L_PTL_G1_1|_RX|P3 _PTL_G1_1|_RX|8 0  5.339e-13
R_PTL_G1_1|_RX|B1 _PTL_G1_1|_RX|1 _PTL_G1_1|_RX|101  4.225701121488
R_PTL_G1_1|_RX|B2 _PTL_G1_1|_RX|4 _PTL_G1_1|_RX|104  3.429952209
R_PTL_G1_1|_RX|B3 _PTL_G1_1|_RX|7 _PTL_G1_1|_RX|107  2.7439617672
L_PTL_G1_1|_RX|RB1 _PTL_G1_1|_RX|101 0  2.38752113364072e-12
L_PTL_G1_1|_RX|RB2 _PTL_G1_1|_RX|104 0  1.937922998085e-12
L_PTL_G1_1|_RX|RB3 _PTL_G1_1|_RX|107 0  1.550338398468e-12
B_PTL_P2_1|_TX|1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|2 JJMIT AREA=2.5
B_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|5 JJMIT AREA=2.5
I_PTL_P2_1|_TX|B1 0 _PTL_P2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P2_1|_TX|B2 0 _PTL_P2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|3  1.684e-12
L_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|6  3.596e-12
L_PTL_P2_1|_TX|1 P2_1_TX _PTL_P2_1|_TX|1  2.063e-12
L_PTL_P2_1|_TX|2 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|4  4.123e-12
L_PTL_P2_1|_TX|3 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|7  2.193e-12
R_PTL_P2_1|_TX|D _PTL_P2_1|_TX|7 _PTL_P2_1|A_PTL  1.36
L_PTL_P2_1|_TX|P1 _PTL_P2_1|_TX|2 0  5.254e-13
L_PTL_P2_1|_TX|P2 _PTL_P2_1|_TX|5 0  5.141e-13
R_PTL_P2_1|_TX|B1 _PTL_P2_1|_TX|1 _PTL_P2_1|_TX|101  2.7439617672
R_PTL_P2_1|_TX|B2 _PTL_P2_1|_TX|4 _PTL_P2_1|_TX|104  2.7439617672
L_PTL_P2_1|_TX|RB1 _PTL_P2_1|_TX|101 0  1.550338398468e-12
L_PTL_P2_1|_TX|RB2 _PTL_P2_1|_TX|104 0  1.550338398468e-12
B_PTL_P2_1|_RX|1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|5 JJMIT AREA=2.0
B_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|8 JJMIT AREA=2.5
I_PTL_P2_1|_RX|B1 0 _PTL_P2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|3  2.777e-12
I_PTL_P2_1|_RX|B2 0 _PTL_P2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|6  2.685e-12
I_PTL_P2_1|_RX|B3 0 _PTL_P2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|9  2.764e-12
L_PTL_P2_1|_RX|1 _PTL_P2_1|A_PTL _PTL_P2_1|_RX|1  1.346e-12
L_PTL_P2_1|_RX|2 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|4  6.348e-12
L_PTL_P2_1|_RX|3 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7  5.197e-12
L_PTL_P2_1|_RX|4 _PTL_P2_1|_RX|7 _PTL_P2_1|D  2.058e-12
L_PTL_P2_1|_RX|P1 _PTL_P2_1|_RX|2 0  4.795e-13
L_PTL_P2_1|_RX|P2 _PTL_P2_1|_RX|5 0  5.431e-13
L_PTL_P2_1|_RX|P3 _PTL_P2_1|_RX|8 0  5.339e-13
R_PTL_P2_1|_RX|B1 _PTL_P2_1|_RX|1 _PTL_P2_1|_RX|101  4.225701121488
R_PTL_P2_1|_RX|B2 _PTL_P2_1|_RX|4 _PTL_P2_1|_RX|104  3.429952209
R_PTL_P2_1|_RX|B3 _PTL_P2_1|_RX|7 _PTL_P2_1|_RX|107  2.7439617672
L_PTL_P2_1|_RX|RB1 _PTL_P2_1|_RX|101 0  2.38752113364072e-12
L_PTL_P2_1|_RX|RB2 _PTL_P2_1|_RX|104 0  1.937922998085e-12
L_PTL_P2_1|_RX|RB3 _PTL_P2_1|_RX|107 0  1.550338398468e-12
L_PTL_P2_1|_SPL|1 _PTL_P2_1|D _PTL_P2_1|_SPL|D1  2e-12
L_PTL_P2_1|_SPL|2 _PTL_P2_1|_SPL|D1 _PTL_P2_1|_SPL|D2  4.135667696e-12
L_PTL_P2_1|_SPL|3 _PTL_P2_1|_SPL|D2 _PTL_P2_1|_SPL|JCT  9.84682784761905e-13
L_PTL_P2_1|_SPL|4 _PTL_P2_1|_SPL|JCT _PTL_P2_1|_SPL|QA1  9.84682784761905e-13
L_PTL_P2_1|_SPL|5 _PTL_P2_1|_SPL|QA1 P2_1_TO2  2e-12
L_PTL_P2_1|_SPL|6 _PTL_P2_1|_SPL|JCT _PTL_P2_1|_SPL|QB1  9.84682784761905e-13
L_PTL_P2_1|_SPL|7 _PTL_P2_1|_SPL|QB1 P2_1_OUT  2e-12
B_PTL_G2_1|_TX|1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|2 JJMIT AREA=2.5
B_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|5 JJMIT AREA=2.5
I_PTL_G2_1|_TX|B1 0 _PTL_G2_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_1|_TX|B2 0 _PTL_G2_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|3  1.684e-12
L_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|6  3.596e-12
L_PTL_G2_1|_TX|1 G2_1_TX _PTL_G2_1|_TX|1  2.063e-12
L_PTL_G2_1|_TX|2 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|4  4.123e-12
L_PTL_G2_1|_TX|3 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|7  2.193e-12
R_PTL_G2_1|_TX|D _PTL_G2_1|_TX|7 _PTL_G2_1|A_PTL  1.36
L_PTL_G2_1|_TX|P1 _PTL_G2_1|_TX|2 0  5.254e-13
L_PTL_G2_1|_TX|P2 _PTL_G2_1|_TX|5 0  5.141e-13
R_PTL_G2_1|_TX|B1 _PTL_G2_1|_TX|1 _PTL_G2_1|_TX|101  2.7439617672
R_PTL_G2_1|_TX|B2 _PTL_G2_1|_TX|4 _PTL_G2_1|_TX|104  2.7439617672
L_PTL_G2_1|_TX|RB1 _PTL_G2_1|_TX|101 0  1.550338398468e-12
L_PTL_G2_1|_TX|RB2 _PTL_G2_1|_TX|104 0  1.550338398468e-12
B_PTL_G2_1|_RX|1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|5 JJMIT AREA=2.0
B_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|8 JJMIT AREA=2.5
I_PTL_G2_1|_RX|B1 0 _PTL_G2_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|3  2.777e-12
I_PTL_G2_1|_RX|B2 0 _PTL_G2_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|6  2.685e-12
I_PTL_G2_1|_RX|B3 0 _PTL_G2_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|9  2.764e-12
L_PTL_G2_1|_RX|1 _PTL_G2_1|A_PTL _PTL_G2_1|_RX|1  1.346e-12
L_PTL_G2_1|_RX|2 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|4  6.348e-12
L_PTL_G2_1|_RX|3 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7  5.197e-12
L_PTL_G2_1|_RX|4 _PTL_G2_1|_RX|7 G2_1_TO2  2.058e-12
L_PTL_G2_1|_RX|P1 _PTL_G2_1|_RX|2 0  4.795e-13
L_PTL_G2_1|_RX|P2 _PTL_G2_1|_RX|5 0  5.431e-13
L_PTL_G2_1|_RX|P3 _PTL_G2_1|_RX|8 0  5.339e-13
R_PTL_G2_1|_RX|B1 _PTL_G2_1|_RX|1 _PTL_G2_1|_RX|101  4.225701121488
R_PTL_G2_1|_RX|B2 _PTL_G2_1|_RX|4 _PTL_G2_1|_RX|104  3.429952209
R_PTL_G2_1|_RX|B3 _PTL_G2_1|_RX|7 _PTL_G2_1|_RX|107  2.7439617672
L_PTL_G2_1|_RX|RB1 _PTL_G2_1|_RX|101 0  2.38752113364072e-12
L_PTL_G2_1|_RX|RB2 _PTL_G2_1|_RX|104 0  1.937922998085e-12
L_PTL_G2_1|_RX|RB3 _PTL_G2_1|_RX|107 0  1.550338398468e-12
B_PTL_P3_1|_TX|1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|2 JJMIT AREA=2.5
B_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|5 JJMIT AREA=2.5
I_PTL_P3_1|_TX|B1 0 _PTL_P3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P3_1|_TX|B2 0 _PTL_P3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|3  1.684e-12
L_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|6  3.596e-12
L_PTL_P3_1|_TX|1 P3_1_TX _PTL_P3_1|_TX|1  2.063e-12
L_PTL_P3_1|_TX|2 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|4  4.123e-12
L_PTL_P3_1|_TX|3 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|7  2.193e-12
R_PTL_P3_1|_TX|D _PTL_P3_1|_TX|7 _PTL_P3_1|A_PTL  1.36
L_PTL_P3_1|_TX|P1 _PTL_P3_1|_TX|2 0  5.254e-13
L_PTL_P3_1|_TX|P2 _PTL_P3_1|_TX|5 0  5.141e-13
R_PTL_P3_1|_TX|B1 _PTL_P3_1|_TX|1 _PTL_P3_1|_TX|101  2.7439617672
R_PTL_P3_1|_TX|B2 _PTL_P3_1|_TX|4 _PTL_P3_1|_TX|104  2.7439617672
L_PTL_P3_1|_TX|RB1 _PTL_P3_1|_TX|101 0  1.550338398468e-12
L_PTL_P3_1|_TX|RB2 _PTL_P3_1|_TX|104 0  1.550338398468e-12
B_PTL_P3_1|_RX|1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|5 JJMIT AREA=2.0
B_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|8 JJMIT AREA=2.5
I_PTL_P3_1|_RX|B1 0 _PTL_P3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|3  2.777e-12
I_PTL_P3_1|_RX|B2 0 _PTL_P3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|6  2.685e-12
I_PTL_P3_1|_RX|B3 0 _PTL_P3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|9  2.764e-12
L_PTL_P3_1|_RX|1 _PTL_P3_1|A_PTL _PTL_P3_1|_RX|1  1.346e-12
L_PTL_P3_1|_RX|2 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|4  6.348e-12
L_PTL_P3_1|_RX|3 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7  5.197e-12
L_PTL_P3_1|_RX|4 _PTL_P3_1|_RX|7 P3_1_TO3  2.058e-12
L_PTL_P3_1|_RX|P1 _PTL_P3_1|_RX|2 0  4.795e-13
L_PTL_P3_1|_RX|P2 _PTL_P3_1|_RX|5 0  5.431e-13
L_PTL_P3_1|_RX|P3 _PTL_P3_1|_RX|8 0  5.339e-13
R_PTL_P3_1|_RX|B1 _PTL_P3_1|_RX|1 _PTL_P3_1|_RX|101  4.225701121488
R_PTL_P3_1|_RX|B2 _PTL_P3_1|_RX|4 _PTL_P3_1|_RX|104  3.429952209
R_PTL_P3_1|_RX|B3 _PTL_P3_1|_RX|7 _PTL_P3_1|_RX|107  2.7439617672
L_PTL_P3_1|_RX|RB1 _PTL_P3_1|_RX|101 0  2.38752113364072e-12
L_PTL_P3_1|_RX|RB2 _PTL_P3_1|_RX|104 0  1.937922998085e-12
L_PTL_P3_1|_RX|RB3 _PTL_P3_1|_RX|107 0  1.550338398468e-12
B_PTL_G3_1|_TX|1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|2 JJMIT AREA=2.5
B_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|5 JJMIT AREA=2.5
I_PTL_G3_1|_TX|B1 0 _PTL_G3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_1|_TX|B2 0 _PTL_G3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|3  1.684e-12
L_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|6  3.596e-12
L_PTL_G3_1|_TX|1 G3_1_TX _PTL_G3_1|_TX|1  2.063e-12
L_PTL_G3_1|_TX|2 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|4  4.123e-12
L_PTL_G3_1|_TX|3 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|7  2.193e-12
R_PTL_G3_1|_TX|D _PTL_G3_1|_TX|7 _PTL_G3_1|A_PTL  1.36
L_PTL_G3_1|_TX|P1 _PTL_G3_1|_TX|2 0  5.254e-13
L_PTL_G3_1|_TX|P2 _PTL_G3_1|_TX|5 0  5.141e-13
R_PTL_G3_1|_TX|B1 _PTL_G3_1|_TX|1 _PTL_G3_1|_TX|101  2.7439617672
R_PTL_G3_1|_TX|B2 _PTL_G3_1|_TX|4 _PTL_G3_1|_TX|104  2.7439617672
L_PTL_G3_1|_TX|RB1 _PTL_G3_1|_TX|101 0  1.550338398468e-12
L_PTL_G3_1|_TX|RB2 _PTL_G3_1|_TX|104 0  1.550338398468e-12
B_PTL_G3_1|_RX|1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|5 JJMIT AREA=2.0
B_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|8 JJMIT AREA=2.5
I_PTL_G3_1|_RX|B1 0 _PTL_G3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|3  2.777e-12
I_PTL_G3_1|_RX|B2 0 _PTL_G3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|6  2.685e-12
I_PTL_G3_1|_RX|B3 0 _PTL_G3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|9  2.764e-12
L_PTL_G3_1|_RX|1 _PTL_G3_1|A_PTL _PTL_G3_1|_RX|1  1.346e-12
L_PTL_G3_1|_RX|2 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|4  6.348e-12
L_PTL_G3_1|_RX|3 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7  5.197e-12
L_PTL_G3_1|_RX|4 _PTL_G3_1|_RX|7 G3_1_TO3  2.058e-12
L_PTL_G3_1|_RX|P1 _PTL_G3_1|_RX|2 0  4.795e-13
L_PTL_G3_1|_RX|P2 _PTL_G3_1|_RX|5 0  5.431e-13
L_PTL_G3_1|_RX|P3 _PTL_G3_1|_RX|8 0  5.339e-13
R_PTL_G3_1|_RX|B1 _PTL_G3_1|_RX|1 _PTL_G3_1|_RX|101  4.225701121488
R_PTL_G3_1|_RX|B2 _PTL_G3_1|_RX|4 _PTL_G3_1|_RX|104  3.429952209
R_PTL_G3_1|_RX|B3 _PTL_G3_1|_RX|7 _PTL_G3_1|_RX|107  2.7439617672
L_PTL_G3_1|_RX|RB1 _PTL_G3_1|_RX|101 0  2.38752113364072e-12
L_PTL_G3_1|_RX|RB2 _PTL_G3_1|_RX|104 0  1.937922998085e-12
L_PTL_G3_1|_RX|RB3 _PTL_G3_1|_RX|107 0  1.550338398468e-12
B_PTL_P4_1|_TX|1 _PTL_P4_1|_TX|1 _PTL_P4_1|_TX|2 JJMIT AREA=2.5
B_PTL_P4_1|_TX|2 _PTL_P4_1|_TX|4 _PTL_P4_1|_TX|5 JJMIT AREA=2.5
I_PTL_P4_1|_TX|B1 0 _PTL_P4_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P4_1|_TX|B2 0 _PTL_P4_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P4_1|_TX|B1 _PTL_P4_1|_TX|1 _PTL_P4_1|_TX|3  1.684e-12
L_PTL_P4_1|_TX|B2 _PTL_P4_1|_TX|4 _PTL_P4_1|_TX|6  3.596e-12
L_PTL_P4_1|_TX|1 P4_1_TX _PTL_P4_1|_TX|1  2.063e-12
L_PTL_P4_1|_TX|2 _PTL_P4_1|_TX|1 _PTL_P4_1|_TX|4  4.123e-12
L_PTL_P4_1|_TX|3 _PTL_P4_1|_TX|4 _PTL_P4_1|_TX|7  2.193e-12
R_PTL_P4_1|_TX|D _PTL_P4_1|_TX|7 _PTL_P4_1|A_PTL  1.36
L_PTL_P4_1|_TX|P1 _PTL_P4_1|_TX|2 0  5.254e-13
L_PTL_P4_1|_TX|P2 _PTL_P4_1|_TX|5 0  5.141e-13
R_PTL_P4_1|_TX|B1 _PTL_P4_1|_TX|1 _PTL_P4_1|_TX|101  2.7439617672
R_PTL_P4_1|_TX|B2 _PTL_P4_1|_TX|4 _PTL_P4_1|_TX|104  2.7439617672
L_PTL_P4_1|_TX|RB1 _PTL_P4_1|_TX|101 0  1.550338398468e-12
L_PTL_P4_1|_TX|RB2 _PTL_P4_1|_TX|104 0  1.550338398468e-12
B_PTL_P4_1|_RX|1 _PTL_P4_1|_RX|1 _PTL_P4_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P4_1|_RX|2 _PTL_P4_1|_RX|4 _PTL_P4_1|_RX|5 JJMIT AREA=2.0
B_PTL_P4_1|_RX|3 _PTL_P4_1|_RX|7 _PTL_P4_1|_RX|8 JJMIT AREA=2.5
I_PTL_P4_1|_RX|B1 0 _PTL_P4_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P4_1|_RX|B1 _PTL_P4_1|_RX|1 _PTL_P4_1|_RX|3  2.777e-12
I_PTL_P4_1|_RX|B2 0 _PTL_P4_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P4_1|_RX|B2 _PTL_P4_1|_RX|4 _PTL_P4_1|_RX|6  2.685e-12
I_PTL_P4_1|_RX|B3 0 _PTL_P4_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P4_1|_RX|B3 _PTL_P4_1|_RX|7 _PTL_P4_1|_RX|9  2.764e-12
L_PTL_P4_1|_RX|1 _PTL_P4_1|A_PTL _PTL_P4_1|_RX|1  1.346e-12
L_PTL_P4_1|_RX|2 _PTL_P4_1|_RX|1 _PTL_P4_1|_RX|4  6.348e-12
L_PTL_P4_1|_RX|3 _PTL_P4_1|_RX|4 _PTL_P4_1|_RX|7  5.197e-12
L_PTL_P4_1|_RX|4 _PTL_P4_1|_RX|7 P4_1_TO4  2.058e-12
L_PTL_P4_1|_RX|P1 _PTL_P4_1|_RX|2 0  4.795e-13
L_PTL_P4_1|_RX|P2 _PTL_P4_1|_RX|5 0  5.431e-13
L_PTL_P4_1|_RX|P3 _PTL_P4_1|_RX|8 0  5.339e-13
R_PTL_P4_1|_RX|B1 _PTL_P4_1|_RX|1 _PTL_P4_1|_RX|101  4.225701121488
R_PTL_P4_1|_RX|B2 _PTL_P4_1|_RX|4 _PTL_P4_1|_RX|104  3.429952209
R_PTL_P4_1|_RX|B3 _PTL_P4_1|_RX|7 _PTL_P4_1|_RX|107  2.7439617672
L_PTL_P4_1|_RX|RB1 _PTL_P4_1|_RX|101 0  2.38752113364072e-12
L_PTL_P4_1|_RX|RB2 _PTL_P4_1|_RX|104 0  1.937922998085e-12
L_PTL_P4_1|_RX|RB3 _PTL_P4_1|_RX|107 0  1.550338398468e-12
B_PTL_G4_1|_TX|1 _PTL_G4_1|_TX|1 _PTL_G4_1|_TX|2 JJMIT AREA=2.5
B_PTL_G4_1|_TX|2 _PTL_G4_1|_TX|4 _PTL_G4_1|_TX|5 JJMIT AREA=2.5
I_PTL_G4_1|_TX|B1 0 _PTL_G4_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G4_1|_TX|B2 0 _PTL_G4_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G4_1|_TX|B1 _PTL_G4_1|_TX|1 _PTL_G4_1|_TX|3  1.684e-12
L_PTL_G4_1|_TX|B2 _PTL_G4_1|_TX|4 _PTL_G4_1|_TX|6  3.596e-12
L_PTL_G4_1|_TX|1 G4_1_TX _PTL_G4_1|_TX|1  2.063e-12
L_PTL_G4_1|_TX|2 _PTL_G4_1|_TX|1 _PTL_G4_1|_TX|4  4.123e-12
L_PTL_G4_1|_TX|3 _PTL_G4_1|_TX|4 _PTL_G4_1|_TX|7  2.193e-12
R_PTL_G4_1|_TX|D _PTL_G4_1|_TX|7 _PTL_G4_1|A_PTL  1.36
L_PTL_G4_1|_TX|P1 _PTL_G4_1|_TX|2 0  5.254e-13
L_PTL_G4_1|_TX|P2 _PTL_G4_1|_TX|5 0  5.141e-13
R_PTL_G4_1|_TX|B1 _PTL_G4_1|_TX|1 _PTL_G4_1|_TX|101  2.7439617672
R_PTL_G4_1|_TX|B2 _PTL_G4_1|_TX|4 _PTL_G4_1|_TX|104  2.7439617672
L_PTL_G4_1|_TX|RB1 _PTL_G4_1|_TX|101 0  1.550338398468e-12
L_PTL_G4_1|_TX|RB2 _PTL_G4_1|_TX|104 0  1.550338398468e-12
B_PTL_G4_1|_RX|1 _PTL_G4_1|_RX|1 _PTL_G4_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G4_1|_RX|2 _PTL_G4_1|_RX|4 _PTL_G4_1|_RX|5 JJMIT AREA=2.0
B_PTL_G4_1|_RX|3 _PTL_G4_1|_RX|7 _PTL_G4_1|_RX|8 JJMIT AREA=2.5
I_PTL_G4_1|_RX|B1 0 _PTL_G4_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G4_1|_RX|B1 _PTL_G4_1|_RX|1 _PTL_G4_1|_RX|3  2.777e-12
I_PTL_G4_1|_RX|B2 0 _PTL_G4_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G4_1|_RX|B2 _PTL_G4_1|_RX|4 _PTL_G4_1|_RX|6  2.685e-12
I_PTL_G4_1|_RX|B3 0 _PTL_G4_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G4_1|_RX|B3 _PTL_G4_1|_RX|7 _PTL_G4_1|_RX|9  2.764e-12
L_PTL_G4_1|_RX|1 _PTL_G4_1|A_PTL _PTL_G4_1|_RX|1  1.346e-12
L_PTL_G4_1|_RX|2 _PTL_G4_1|_RX|1 _PTL_G4_1|_RX|4  6.348e-12
L_PTL_G4_1|_RX|3 _PTL_G4_1|_RX|4 _PTL_G4_1|_RX|7  5.197e-12
L_PTL_G4_1|_RX|4 _PTL_G4_1|_RX|7 G4_1_TO4  2.058e-12
L_PTL_G4_1|_RX|P1 _PTL_G4_1|_RX|2 0  4.795e-13
L_PTL_G4_1|_RX|P2 _PTL_G4_1|_RX|5 0  5.431e-13
L_PTL_G4_1|_RX|P3 _PTL_G4_1|_RX|8 0  5.339e-13
R_PTL_G4_1|_RX|B1 _PTL_G4_1|_RX|1 _PTL_G4_1|_RX|101  4.225701121488
R_PTL_G4_1|_RX|B2 _PTL_G4_1|_RX|4 _PTL_G4_1|_RX|104  3.429952209
R_PTL_G4_1|_RX|B3 _PTL_G4_1|_RX|7 _PTL_G4_1|_RX|107  2.7439617672
L_PTL_G4_1|_RX|RB1 _PTL_G4_1|_RX|101 0  2.38752113364072e-12
L_PTL_G4_1|_RX|RB2 _PTL_G4_1|_RX|104 0  1.937922998085e-12
L_PTL_G4_1|_RX|RB3 _PTL_G4_1|_RX|107 0  1.550338398468e-12
B_PTL_P5_1|_TX|1 _PTL_P5_1|_TX|1 _PTL_P5_1|_TX|2 JJMIT AREA=2.5
B_PTL_P5_1|_TX|2 _PTL_P5_1|_TX|4 _PTL_P5_1|_TX|5 JJMIT AREA=2.5
I_PTL_P5_1|_TX|B1 0 _PTL_P5_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P5_1|_TX|B2 0 _PTL_P5_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P5_1|_TX|B1 _PTL_P5_1|_TX|1 _PTL_P5_1|_TX|3  1.684e-12
L_PTL_P5_1|_TX|B2 _PTL_P5_1|_TX|4 _PTL_P5_1|_TX|6  3.596e-12
L_PTL_P5_1|_TX|1 P5_1_TX _PTL_P5_1|_TX|1  2.063e-12
L_PTL_P5_1|_TX|2 _PTL_P5_1|_TX|1 _PTL_P5_1|_TX|4  4.123e-12
L_PTL_P5_1|_TX|3 _PTL_P5_1|_TX|4 _PTL_P5_1|_TX|7  2.193e-12
R_PTL_P5_1|_TX|D _PTL_P5_1|_TX|7 _PTL_P5_1|A_PTL  1.36
L_PTL_P5_1|_TX|P1 _PTL_P5_1|_TX|2 0  5.254e-13
L_PTL_P5_1|_TX|P2 _PTL_P5_1|_TX|5 0  5.141e-13
R_PTL_P5_1|_TX|B1 _PTL_P5_1|_TX|1 _PTL_P5_1|_TX|101  2.7439617672
R_PTL_P5_1|_TX|B2 _PTL_P5_1|_TX|4 _PTL_P5_1|_TX|104  2.7439617672
L_PTL_P5_1|_TX|RB1 _PTL_P5_1|_TX|101 0  1.550338398468e-12
L_PTL_P5_1|_TX|RB2 _PTL_P5_1|_TX|104 0  1.550338398468e-12
B_PTL_P5_1|_RX|1 _PTL_P5_1|_RX|1 _PTL_P5_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P5_1|_RX|2 _PTL_P5_1|_RX|4 _PTL_P5_1|_RX|5 JJMIT AREA=2.0
B_PTL_P5_1|_RX|3 _PTL_P5_1|_RX|7 _PTL_P5_1|_RX|8 JJMIT AREA=2.5
I_PTL_P5_1|_RX|B1 0 _PTL_P5_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P5_1|_RX|B1 _PTL_P5_1|_RX|1 _PTL_P5_1|_RX|3  2.777e-12
I_PTL_P5_1|_RX|B2 0 _PTL_P5_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P5_1|_RX|B2 _PTL_P5_1|_RX|4 _PTL_P5_1|_RX|6  2.685e-12
I_PTL_P5_1|_RX|B3 0 _PTL_P5_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P5_1|_RX|B3 _PTL_P5_1|_RX|7 _PTL_P5_1|_RX|9  2.764e-12
L_PTL_P5_1|_RX|1 _PTL_P5_1|A_PTL _PTL_P5_1|_RX|1  1.346e-12
L_PTL_P5_1|_RX|2 _PTL_P5_1|_RX|1 _PTL_P5_1|_RX|4  6.348e-12
L_PTL_P5_1|_RX|3 _PTL_P5_1|_RX|4 _PTL_P5_1|_RX|7  5.197e-12
L_PTL_P5_1|_RX|4 _PTL_P5_1|_RX|7 _PTL_P5_1|D  2.058e-12
L_PTL_P5_1|_RX|P1 _PTL_P5_1|_RX|2 0  4.795e-13
L_PTL_P5_1|_RX|P2 _PTL_P5_1|_RX|5 0  5.431e-13
L_PTL_P5_1|_RX|P3 _PTL_P5_1|_RX|8 0  5.339e-13
R_PTL_P5_1|_RX|B1 _PTL_P5_1|_RX|1 _PTL_P5_1|_RX|101  4.225701121488
R_PTL_P5_1|_RX|B2 _PTL_P5_1|_RX|4 _PTL_P5_1|_RX|104  3.429952209
R_PTL_P5_1|_RX|B3 _PTL_P5_1|_RX|7 _PTL_P5_1|_RX|107  2.7439617672
L_PTL_P5_1|_RX|RB1 _PTL_P5_1|_RX|101 0  2.38752113364072e-12
L_PTL_P5_1|_RX|RB2 _PTL_P5_1|_RX|104 0  1.937922998085e-12
L_PTL_P5_1|_RX|RB3 _PTL_P5_1|_RX|107 0  1.550338398468e-12
L_PTL_P5_1|_SPL|1 _PTL_P5_1|D _PTL_P5_1|_SPL|D1  2e-12
L_PTL_P5_1|_SPL|2 _PTL_P5_1|_SPL|D1 _PTL_P5_1|_SPL|D2  4.135667696e-12
L_PTL_P5_1|_SPL|3 _PTL_P5_1|_SPL|D2 _PTL_P5_1|_SPL|JCT  9.84682784761905e-13
L_PTL_P5_1|_SPL|4 _PTL_P5_1|_SPL|JCT _PTL_P5_1|_SPL|QA1  9.84682784761905e-13
L_PTL_P5_1|_SPL|5 _PTL_P5_1|_SPL|QA1 P5_1_TO5  2e-12
L_PTL_P5_1|_SPL|6 _PTL_P5_1|_SPL|JCT _PTL_P5_1|_SPL|QB1  9.84682784761905e-13
L_PTL_P5_1|_SPL|7 _PTL_P5_1|_SPL|QB1 P5_1_TO7  2e-12
B_PTL_G5_1|_TX|1 _PTL_G5_1|_TX|1 _PTL_G5_1|_TX|2 JJMIT AREA=2.5
B_PTL_G5_1|_TX|2 _PTL_G5_1|_TX|4 _PTL_G5_1|_TX|5 JJMIT AREA=2.5
I_PTL_G5_1|_TX|B1 0 _PTL_G5_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G5_1|_TX|B2 0 _PTL_G5_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G5_1|_TX|B1 _PTL_G5_1|_TX|1 _PTL_G5_1|_TX|3  1.684e-12
L_PTL_G5_1|_TX|B2 _PTL_G5_1|_TX|4 _PTL_G5_1|_TX|6  3.596e-12
L_PTL_G5_1|_TX|1 G5_1_TX _PTL_G5_1|_TX|1  2.063e-12
L_PTL_G5_1|_TX|2 _PTL_G5_1|_TX|1 _PTL_G5_1|_TX|4  4.123e-12
L_PTL_G5_1|_TX|3 _PTL_G5_1|_TX|4 _PTL_G5_1|_TX|7  2.193e-12
R_PTL_G5_1|_TX|D _PTL_G5_1|_TX|7 _PTL_G5_1|A_PTL  1.36
L_PTL_G5_1|_TX|P1 _PTL_G5_1|_TX|2 0  5.254e-13
L_PTL_G5_1|_TX|P2 _PTL_G5_1|_TX|5 0  5.141e-13
R_PTL_G5_1|_TX|B1 _PTL_G5_1|_TX|1 _PTL_G5_1|_TX|101  2.7439617672
R_PTL_G5_1|_TX|B2 _PTL_G5_1|_TX|4 _PTL_G5_1|_TX|104  2.7439617672
L_PTL_G5_1|_TX|RB1 _PTL_G5_1|_TX|101 0  1.550338398468e-12
L_PTL_G5_1|_TX|RB2 _PTL_G5_1|_TX|104 0  1.550338398468e-12
B_PTL_G5_1|_RX|1 _PTL_G5_1|_RX|1 _PTL_G5_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G5_1|_RX|2 _PTL_G5_1|_RX|4 _PTL_G5_1|_RX|5 JJMIT AREA=2.0
B_PTL_G5_1|_RX|3 _PTL_G5_1|_RX|7 _PTL_G5_1|_RX|8 JJMIT AREA=2.5
I_PTL_G5_1|_RX|B1 0 _PTL_G5_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G5_1|_RX|B1 _PTL_G5_1|_RX|1 _PTL_G5_1|_RX|3  2.777e-12
I_PTL_G5_1|_RX|B2 0 _PTL_G5_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G5_1|_RX|B2 _PTL_G5_1|_RX|4 _PTL_G5_1|_RX|6  2.685e-12
I_PTL_G5_1|_RX|B3 0 _PTL_G5_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G5_1|_RX|B3 _PTL_G5_1|_RX|7 _PTL_G5_1|_RX|9  2.764e-12
L_PTL_G5_1|_RX|1 _PTL_G5_1|A_PTL _PTL_G5_1|_RX|1  1.346e-12
L_PTL_G5_1|_RX|2 _PTL_G5_1|_RX|1 _PTL_G5_1|_RX|4  6.348e-12
L_PTL_G5_1|_RX|3 _PTL_G5_1|_RX|4 _PTL_G5_1|_RX|7  5.197e-12
L_PTL_G5_1|_RX|4 _PTL_G5_1|_RX|7 _PTL_G5_1|D  2.058e-12
L_PTL_G5_1|_RX|P1 _PTL_G5_1|_RX|2 0  4.795e-13
L_PTL_G5_1|_RX|P2 _PTL_G5_1|_RX|5 0  5.431e-13
L_PTL_G5_1|_RX|P3 _PTL_G5_1|_RX|8 0  5.339e-13
R_PTL_G5_1|_RX|B1 _PTL_G5_1|_RX|1 _PTL_G5_1|_RX|101  4.225701121488
R_PTL_G5_1|_RX|B2 _PTL_G5_1|_RX|4 _PTL_G5_1|_RX|104  3.429952209
R_PTL_G5_1|_RX|B3 _PTL_G5_1|_RX|7 _PTL_G5_1|_RX|107  2.7439617672
L_PTL_G5_1|_RX|RB1 _PTL_G5_1|_RX|101 0  2.38752113364072e-12
L_PTL_G5_1|_RX|RB2 _PTL_G5_1|_RX|104 0  1.937922998085e-12
L_PTL_G5_1|_RX|RB3 _PTL_G5_1|_RX|107 0  1.550338398468e-12
L_PTL_G5_1|_SPL|1 _PTL_G5_1|D _PTL_G5_1|_SPL|D1  2e-12
L_PTL_G5_1|_SPL|2 _PTL_G5_1|_SPL|D1 _PTL_G5_1|_SPL|D2  4.135667696e-12
L_PTL_G5_1|_SPL|3 _PTL_G5_1|_SPL|D2 _PTL_G5_1|_SPL|JCT  9.84682784761905e-13
L_PTL_G5_1|_SPL|4 _PTL_G5_1|_SPL|JCT _PTL_G5_1|_SPL|QA1  9.84682784761905e-13
L_PTL_G5_1|_SPL|5 _PTL_G5_1|_SPL|QA1 G5_1_TO5  2e-12
L_PTL_G5_1|_SPL|6 _PTL_G5_1|_SPL|JCT _PTL_G5_1|_SPL|QB1  9.84682784761905e-13
L_PTL_G5_1|_SPL|7 _PTL_G5_1|_SPL|QB1 G5_1_TO7  2e-12
B_PTL_P6_1|_TX|1 _PTL_P6_1|_TX|1 _PTL_P6_1|_TX|2 JJMIT AREA=2.5
B_PTL_P6_1|_TX|2 _PTL_P6_1|_TX|4 _PTL_P6_1|_TX|5 JJMIT AREA=2.5
I_PTL_P6_1|_TX|B1 0 _PTL_P6_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P6_1|_TX|B2 0 _PTL_P6_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P6_1|_TX|B1 _PTL_P6_1|_TX|1 _PTL_P6_1|_TX|3  1.684e-12
L_PTL_P6_1|_TX|B2 _PTL_P6_1|_TX|4 _PTL_P6_1|_TX|6  3.596e-12
L_PTL_P6_1|_TX|1 P6_1_TX _PTL_P6_1|_TX|1  2.063e-12
L_PTL_P6_1|_TX|2 _PTL_P6_1|_TX|1 _PTL_P6_1|_TX|4  4.123e-12
L_PTL_P6_1|_TX|3 _PTL_P6_1|_TX|4 _PTL_P6_1|_TX|7  2.193e-12
R_PTL_P6_1|_TX|D _PTL_P6_1|_TX|7 _PTL_P6_1|A_PTL  1.36
L_PTL_P6_1|_TX|P1 _PTL_P6_1|_TX|2 0  5.254e-13
L_PTL_P6_1|_TX|P2 _PTL_P6_1|_TX|5 0  5.141e-13
R_PTL_P6_1|_TX|B1 _PTL_P6_1|_TX|1 _PTL_P6_1|_TX|101  2.7439617672
R_PTL_P6_1|_TX|B2 _PTL_P6_1|_TX|4 _PTL_P6_1|_TX|104  2.7439617672
L_PTL_P6_1|_TX|RB1 _PTL_P6_1|_TX|101 0  1.550338398468e-12
L_PTL_P6_1|_TX|RB2 _PTL_P6_1|_TX|104 0  1.550338398468e-12
B_PTL_P6_1|_RX|1 _PTL_P6_1|_RX|1 _PTL_P6_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P6_1|_RX|2 _PTL_P6_1|_RX|4 _PTL_P6_1|_RX|5 JJMIT AREA=2.0
B_PTL_P6_1|_RX|3 _PTL_P6_1|_RX|7 _PTL_P6_1|_RX|8 JJMIT AREA=2.5
I_PTL_P6_1|_RX|B1 0 _PTL_P6_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P6_1|_RX|B1 _PTL_P6_1|_RX|1 _PTL_P6_1|_RX|3  2.777e-12
I_PTL_P6_1|_RX|B2 0 _PTL_P6_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P6_1|_RX|B2 _PTL_P6_1|_RX|4 _PTL_P6_1|_RX|6  2.685e-12
I_PTL_P6_1|_RX|B3 0 _PTL_P6_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P6_1|_RX|B3 _PTL_P6_1|_RX|7 _PTL_P6_1|_RX|9  2.764e-12
L_PTL_P6_1|_RX|1 _PTL_P6_1|A_PTL _PTL_P6_1|_RX|1  1.346e-12
L_PTL_P6_1|_RX|2 _PTL_P6_1|_RX|1 _PTL_P6_1|_RX|4  6.348e-12
L_PTL_P6_1|_RX|3 _PTL_P6_1|_RX|4 _PTL_P6_1|_RX|7  5.197e-12
L_PTL_P6_1|_RX|4 _PTL_P6_1|_RX|7 P6_1_TO6  2.058e-12
L_PTL_P6_1|_RX|P1 _PTL_P6_1|_RX|2 0  4.795e-13
L_PTL_P6_1|_RX|P2 _PTL_P6_1|_RX|5 0  5.431e-13
L_PTL_P6_1|_RX|P3 _PTL_P6_1|_RX|8 0  5.339e-13
R_PTL_P6_1|_RX|B1 _PTL_P6_1|_RX|1 _PTL_P6_1|_RX|101  4.225701121488
R_PTL_P6_1|_RX|B2 _PTL_P6_1|_RX|4 _PTL_P6_1|_RX|104  3.429952209
R_PTL_P6_1|_RX|B3 _PTL_P6_1|_RX|7 _PTL_P6_1|_RX|107  2.7439617672
L_PTL_P6_1|_RX|RB1 _PTL_P6_1|_RX|101 0  2.38752113364072e-12
L_PTL_P6_1|_RX|RB2 _PTL_P6_1|_RX|104 0  1.937922998085e-12
L_PTL_P6_1|_RX|RB3 _PTL_P6_1|_RX|107 0  1.550338398468e-12
B_PTL_G6_1|_TX|1 _PTL_G6_1|_TX|1 _PTL_G6_1|_TX|2 JJMIT AREA=2.5
B_PTL_G6_1|_TX|2 _PTL_G6_1|_TX|4 _PTL_G6_1|_TX|5 JJMIT AREA=2.5
I_PTL_G6_1|_TX|B1 0 _PTL_G6_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G6_1|_TX|B2 0 _PTL_G6_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G6_1|_TX|B1 _PTL_G6_1|_TX|1 _PTL_G6_1|_TX|3  1.684e-12
L_PTL_G6_1|_TX|B2 _PTL_G6_1|_TX|4 _PTL_G6_1|_TX|6  3.596e-12
L_PTL_G6_1|_TX|1 G6_1_TX _PTL_G6_1|_TX|1  2.063e-12
L_PTL_G6_1|_TX|2 _PTL_G6_1|_TX|1 _PTL_G6_1|_TX|4  4.123e-12
L_PTL_G6_1|_TX|3 _PTL_G6_1|_TX|4 _PTL_G6_1|_TX|7  2.193e-12
R_PTL_G6_1|_TX|D _PTL_G6_1|_TX|7 _PTL_G6_1|A_PTL  1.36
L_PTL_G6_1|_TX|P1 _PTL_G6_1|_TX|2 0  5.254e-13
L_PTL_G6_1|_TX|P2 _PTL_G6_1|_TX|5 0  5.141e-13
R_PTL_G6_1|_TX|B1 _PTL_G6_1|_TX|1 _PTL_G6_1|_TX|101  2.7439617672
R_PTL_G6_1|_TX|B2 _PTL_G6_1|_TX|4 _PTL_G6_1|_TX|104  2.7439617672
L_PTL_G6_1|_TX|RB1 _PTL_G6_1|_TX|101 0  1.550338398468e-12
L_PTL_G6_1|_TX|RB2 _PTL_G6_1|_TX|104 0  1.550338398468e-12
B_PTL_G6_1|_RX|1 _PTL_G6_1|_RX|1 _PTL_G6_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G6_1|_RX|2 _PTL_G6_1|_RX|4 _PTL_G6_1|_RX|5 JJMIT AREA=2.0
B_PTL_G6_1|_RX|3 _PTL_G6_1|_RX|7 _PTL_G6_1|_RX|8 JJMIT AREA=2.5
I_PTL_G6_1|_RX|B1 0 _PTL_G6_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G6_1|_RX|B1 _PTL_G6_1|_RX|1 _PTL_G6_1|_RX|3  2.777e-12
I_PTL_G6_1|_RX|B2 0 _PTL_G6_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G6_1|_RX|B2 _PTL_G6_1|_RX|4 _PTL_G6_1|_RX|6  2.685e-12
I_PTL_G6_1|_RX|B3 0 _PTL_G6_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G6_1|_RX|B3 _PTL_G6_1|_RX|7 _PTL_G6_1|_RX|9  2.764e-12
L_PTL_G6_1|_RX|1 _PTL_G6_1|A_PTL _PTL_G6_1|_RX|1  1.346e-12
L_PTL_G6_1|_RX|2 _PTL_G6_1|_RX|1 _PTL_G6_1|_RX|4  6.348e-12
L_PTL_G6_1|_RX|3 _PTL_G6_1|_RX|4 _PTL_G6_1|_RX|7  5.197e-12
L_PTL_G6_1|_RX|4 _PTL_G6_1|_RX|7 G6_1_TO6  2.058e-12
L_PTL_G6_1|_RX|P1 _PTL_G6_1|_RX|2 0  4.795e-13
L_PTL_G6_1|_RX|P2 _PTL_G6_1|_RX|5 0  5.431e-13
L_PTL_G6_1|_RX|P3 _PTL_G6_1|_RX|8 0  5.339e-13
R_PTL_G6_1|_RX|B1 _PTL_G6_1|_RX|1 _PTL_G6_1|_RX|101  4.225701121488
R_PTL_G6_1|_RX|B2 _PTL_G6_1|_RX|4 _PTL_G6_1|_RX|104  3.429952209
R_PTL_G6_1|_RX|B3 _PTL_G6_1|_RX|7 _PTL_G6_1|_RX|107  2.7439617672
L_PTL_G6_1|_RX|RB1 _PTL_G6_1|_RX|101 0  2.38752113364072e-12
L_PTL_G6_1|_RX|RB2 _PTL_G6_1|_RX|104 0  1.937922998085e-12
L_PTL_G6_1|_RX|RB3 _PTL_G6_1|_RX|107 0  1.550338398468e-12
B_PTL_P7_1|_TX|1 _PTL_P7_1|_TX|1 _PTL_P7_1|_TX|2 JJMIT AREA=2.5
B_PTL_P7_1|_TX|2 _PTL_P7_1|_TX|4 _PTL_P7_1|_TX|5 JJMIT AREA=2.5
I_PTL_P7_1|_TX|B1 0 _PTL_P7_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P7_1|_TX|B2 0 _PTL_P7_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P7_1|_TX|B1 _PTL_P7_1|_TX|1 _PTL_P7_1|_TX|3  1.684e-12
L_PTL_P7_1|_TX|B2 _PTL_P7_1|_TX|4 _PTL_P7_1|_TX|6  3.596e-12
L_PTL_P7_1|_TX|1 P7_1_TX _PTL_P7_1|_TX|1  2.063e-12
L_PTL_P7_1|_TX|2 _PTL_P7_1|_TX|1 _PTL_P7_1|_TX|4  4.123e-12
L_PTL_P7_1|_TX|3 _PTL_P7_1|_TX|4 _PTL_P7_1|_TX|7  2.193e-12
R_PTL_P7_1|_TX|D _PTL_P7_1|_TX|7 _PTL_P7_1|A_PTL  1.36
L_PTL_P7_1|_TX|P1 _PTL_P7_1|_TX|2 0  5.254e-13
L_PTL_P7_1|_TX|P2 _PTL_P7_1|_TX|5 0  5.141e-13
R_PTL_P7_1|_TX|B1 _PTL_P7_1|_TX|1 _PTL_P7_1|_TX|101  2.7439617672
R_PTL_P7_1|_TX|B2 _PTL_P7_1|_TX|4 _PTL_P7_1|_TX|104  2.7439617672
L_PTL_P7_1|_TX|RB1 _PTL_P7_1|_TX|101 0  1.550338398468e-12
L_PTL_P7_1|_TX|RB2 _PTL_P7_1|_TX|104 0  1.550338398468e-12
B_PTL_P7_1|_RX|1 _PTL_P7_1|_RX|1 _PTL_P7_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P7_1|_RX|2 _PTL_P7_1|_RX|4 _PTL_P7_1|_RX|5 JJMIT AREA=2.0
B_PTL_P7_1|_RX|3 _PTL_P7_1|_RX|7 _PTL_P7_1|_RX|8 JJMIT AREA=2.5
I_PTL_P7_1|_RX|B1 0 _PTL_P7_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P7_1|_RX|B1 _PTL_P7_1|_RX|1 _PTL_P7_1|_RX|3  2.777e-12
I_PTL_P7_1|_RX|B2 0 _PTL_P7_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P7_1|_RX|B2 _PTL_P7_1|_RX|4 _PTL_P7_1|_RX|6  2.685e-12
I_PTL_P7_1|_RX|B3 0 _PTL_P7_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P7_1|_RX|B3 _PTL_P7_1|_RX|7 _PTL_P7_1|_RX|9  2.764e-12
L_PTL_P7_1|_RX|1 _PTL_P7_1|A_PTL _PTL_P7_1|_RX|1  1.346e-12
L_PTL_P7_1|_RX|2 _PTL_P7_1|_RX|1 _PTL_P7_1|_RX|4  6.348e-12
L_PTL_P7_1|_RX|3 _PTL_P7_1|_RX|4 _PTL_P7_1|_RX|7  5.197e-12
L_PTL_P7_1|_RX|4 _PTL_P7_1|_RX|7 P7_1_TO7  2.058e-12
L_PTL_P7_1|_RX|P1 _PTL_P7_1|_RX|2 0  4.795e-13
L_PTL_P7_1|_RX|P2 _PTL_P7_1|_RX|5 0  5.431e-13
L_PTL_P7_1|_RX|P3 _PTL_P7_1|_RX|8 0  5.339e-13
R_PTL_P7_1|_RX|B1 _PTL_P7_1|_RX|1 _PTL_P7_1|_RX|101  4.225701121488
R_PTL_P7_1|_RX|B2 _PTL_P7_1|_RX|4 _PTL_P7_1|_RX|104  3.429952209
R_PTL_P7_1|_RX|B3 _PTL_P7_1|_RX|7 _PTL_P7_1|_RX|107  2.7439617672
L_PTL_P7_1|_RX|RB1 _PTL_P7_1|_RX|101 0  2.38752113364072e-12
L_PTL_P7_1|_RX|RB2 _PTL_P7_1|_RX|104 0  1.937922998085e-12
L_PTL_P7_1|_RX|RB3 _PTL_P7_1|_RX|107 0  1.550338398468e-12
B_PTL_G7_1|_TX|1 _PTL_G7_1|_TX|1 _PTL_G7_1|_TX|2 JJMIT AREA=2.5
B_PTL_G7_1|_TX|2 _PTL_G7_1|_TX|4 _PTL_G7_1|_TX|5 JJMIT AREA=2.5
I_PTL_G7_1|_TX|B1 0 _PTL_G7_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G7_1|_TX|B2 0 _PTL_G7_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G7_1|_TX|B1 _PTL_G7_1|_TX|1 _PTL_G7_1|_TX|3  1.684e-12
L_PTL_G7_1|_TX|B2 _PTL_G7_1|_TX|4 _PTL_G7_1|_TX|6  3.596e-12
L_PTL_G7_1|_TX|1 G7_1_TX _PTL_G7_1|_TX|1  2.063e-12
L_PTL_G7_1|_TX|2 _PTL_G7_1|_TX|1 _PTL_G7_1|_TX|4  4.123e-12
L_PTL_G7_1|_TX|3 _PTL_G7_1|_TX|4 _PTL_G7_1|_TX|7  2.193e-12
R_PTL_G7_1|_TX|D _PTL_G7_1|_TX|7 _PTL_G7_1|A_PTL  1.36
L_PTL_G7_1|_TX|P1 _PTL_G7_1|_TX|2 0  5.254e-13
L_PTL_G7_1|_TX|P2 _PTL_G7_1|_TX|5 0  5.141e-13
R_PTL_G7_1|_TX|B1 _PTL_G7_1|_TX|1 _PTL_G7_1|_TX|101  2.7439617672
R_PTL_G7_1|_TX|B2 _PTL_G7_1|_TX|4 _PTL_G7_1|_TX|104  2.7439617672
L_PTL_G7_1|_TX|RB1 _PTL_G7_1|_TX|101 0  1.550338398468e-12
L_PTL_G7_1|_TX|RB2 _PTL_G7_1|_TX|104 0  1.550338398468e-12
B_PTL_G7_1|_RX|1 _PTL_G7_1|_RX|1 _PTL_G7_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G7_1|_RX|2 _PTL_G7_1|_RX|4 _PTL_G7_1|_RX|5 JJMIT AREA=2.0
B_PTL_G7_1|_RX|3 _PTL_G7_1|_RX|7 _PTL_G7_1|_RX|8 JJMIT AREA=2.5
I_PTL_G7_1|_RX|B1 0 _PTL_G7_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G7_1|_RX|B1 _PTL_G7_1|_RX|1 _PTL_G7_1|_RX|3  2.777e-12
I_PTL_G7_1|_RX|B2 0 _PTL_G7_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G7_1|_RX|B2 _PTL_G7_1|_RX|4 _PTL_G7_1|_RX|6  2.685e-12
I_PTL_G7_1|_RX|B3 0 _PTL_G7_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G7_1|_RX|B3 _PTL_G7_1|_RX|7 _PTL_G7_1|_RX|9  2.764e-12
L_PTL_G7_1|_RX|1 _PTL_G7_1|A_PTL _PTL_G7_1|_RX|1  1.346e-12
L_PTL_G7_1|_RX|2 _PTL_G7_1|_RX|1 _PTL_G7_1|_RX|4  6.348e-12
L_PTL_G7_1|_RX|3 _PTL_G7_1|_RX|4 _PTL_G7_1|_RX|7  5.197e-12
L_PTL_G7_1|_RX|4 _PTL_G7_1|_RX|7 G7_1_TO7  2.058e-12
L_PTL_G7_1|_RX|P1 _PTL_G7_1|_RX|2 0  4.795e-13
L_PTL_G7_1|_RX|P2 _PTL_G7_1|_RX|5 0  5.431e-13
L_PTL_G7_1|_RX|P3 _PTL_G7_1|_RX|8 0  5.339e-13
R_PTL_G7_1|_RX|B1 _PTL_G7_1|_RX|1 _PTL_G7_1|_RX|101  4.225701121488
R_PTL_G7_1|_RX|B2 _PTL_G7_1|_RX|4 _PTL_G7_1|_RX|104  3.429952209
R_PTL_G7_1|_RX|B3 _PTL_G7_1|_RX|7 _PTL_G7_1|_RX|107  2.7439617672
L_PTL_G7_1|_RX|RB1 _PTL_G7_1|_RX|101 0  2.38752113364072e-12
L_PTL_G7_1|_RX|RB2 _PTL_G7_1|_RX|104 0  1.937922998085e-12
L_PTL_G7_1|_RX|RB3 _PTL_G7_1|_RX|107 0  1.550338398468e-12
B_PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_1|_TX|B1 0 _PTL_IP3_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_1|_TX|B2 0 _PTL_IP3_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|3  1.684e-12
L_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|6  3.596e-12
L_PTL_IP3_1|_TX|1 IP3_1_OUT_TX _PTL_IP3_1|_TX|1  2.063e-12
L_PTL_IP3_1|_TX|2 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|4  4.123e-12
L_PTL_IP3_1|_TX|3 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|7  2.193e-12
R_PTL_IP3_1|_TX|D _PTL_IP3_1|_TX|7 _PTL_IP3_1|A_PTL  1.36
L_PTL_IP3_1|_TX|P1 _PTL_IP3_1|_TX|2 0  5.254e-13
L_PTL_IP3_1|_TX|P2 _PTL_IP3_1|_TX|5 0  5.141e-13
R_PTL_IP3_1|_TX|B1 _PTL_IP3_1|_TX|1 _PTL_IP3_1|_TX|101  2.7439617672
R_PTL_IP3_1|_TX|B2 _PTL_IP3_1|_TX|4 _PTL_IP3_1|_TX|104  2.7439617672
L_PTL_IP3_1|_TX|RB1 _PTL_IP3_1|_TX|101 0  1.550338398468e-12
L_PTL_IP3_1|_TX|RB2 _PTL_IP3_1|_TX|104 0  1.550338398468e-12
B_PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_1|_RX|B1 0 _PTL_IP3_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|3  2.777e-12
I_PTL_IP3_1|_RX|B2 0 _PTL_IP3_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|6  2.685e-12
I_PTL_IP3_1|_RX|B3 0 _PTL_IP3_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|9  2.764e-12
L_PTL_IP3_1|_RX|1 _PTL_IP3_1|A_PTL _PTL_IP3_1|_RX|1  1.346e-12
L_PTL_IP3_1|_RX|2 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|4  6.348e-12
L_PTL_IP3_1|_RX|3 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7  5.197e-12
L_PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|7 IP3_1_OUT  2.058e-12
L_PTL_IP3_1|_RX|P1 _PTL_IP3_1|_RX|2 0  4.795e-13
L_PTL_IP3_1|_RX|P2 _PTL_IP3_1|_RX|5 0  5.431e-13
L_PTL_IP3_1|_RX|P3 _PTL_IP3_1|_RX|8 0  5.339e-13
R_PTL_IP3_1|_RX|B1 _PTL_IP3_1|_RX|1 _PTL_IP3_1|_RX|101  4.225701121488
R_PTL_IP3_1|_RX|B2 _PTL_IP3_1|_RX|4 _PTL_IP3_1|_RX|104  3.429952209
R_PTL_IP3_1|_RX|B3 _PTL_IP3_1|_RX|7 _PTL_IP3_1|_RX|107  2.7439617672
L_PTL_IP3_1|_RX|RB1 _PTL_IP3_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_1|_RX|RB2 _PTL_IP3_1|_RX|104 0  1.937922998085e-12
L_PTL_IP3_1|_RX|RB3 _PTL_IP3_1|_RX|107 0  1.550338398468e-12
B_PTL_IP5_1|_TX|1 _PTL_IP5_1|_TX|1 _PTL_IP5_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP5_1|_TX|2 _PTL_IP5_1|_TX|4 _PTL_IP5_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP5_1|_TX|B1 0 _PTL_IP5_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP5_1|_TX|B2 0 _PTL_IP5_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_1|_TX|B1 _PTL_IP5_1|_TX|1 _PTL_IP5_1|_TX|3  1.684e-12
L_PTL_IP5_1|_TX|B2 _PTL_IP5_1|_TX|4 _PTL_IP5_1|_TX|6  3.596e-12
L_PTL_IP5_1|_TX|1 IP5_1_OUT_TX _PTL_IP5_1|_TX|1  2.063e-12
L_PTL_IP5_1|_TX|2 _PTL_IP5_1|_TX|1 _PTL_IP5_1|_TX|4  4.123e-12
L_PTL_IP5_1|_TX|3 _PTL_IP5_1|_TX|4 _PTL_IP5_1|_TX|7  2.193e-12
R_PTL_IP5_1|_TX|D _PTL_IP5_1|_TX|7 _PTL_IP5_1|A_PTL  1.36
L_PTL_IP5_1|_TX|P1 _PTL_IP5_1|_TX|2 0  5.254e-13
L_PTL_IP5_1|_TX|P2 _PTL_IP5_1|_TX|5 0  5.141e-13
R_PTL_IP5_1|_TX|B1 _PTL_IP5_1|_TX|1 _PTL_IP5_1|_TX|101  2.7439617672
R_PTL_IP5_1|_TX|B2 _PTL_IP5_1|_TX|4 _PTL_IP5_1|_TX|104  2.7439617672
L_PTL_IP5_1|_TX|RB1 _PTL_IP5_1|_TX|101 0  1.550338398468e-12
L_PTL_IP5_1|_TX|RB2 _PTL_IP5_1|_TX|104 0  1.550338398468e-12
B_PTL_IP5_1|_RX|1 _PTL_IP5_1|_RX|1 _PTL_IP5_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP5_1|_RX|2 _PTL_IP5_1|_RX|4 _PTL_IP5_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP5_1|_RX|3 _PTL_IP5_1|_RX|7 _PTL_IP5_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP5_1|_RX|B1 0 _PTL_IP5_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP5_1|_RX|B1 _PTL_IP5_1|_RX|1 _PTL_IP5_1|_RX|3  2.777e-12
I_PTL_IP5_1|_RX|B2 0 _PTL_IP5_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP5_1|_RX|B2 _PTL_IP5_1|_RX|4 _PTL_IP5_1|_RX|6  2.685e-12
I_PTL_IP5_1|_RX|B3 0 _PTL_IP5_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_1|_RX|B3 _PTL_IP5_1|_RX|7 _PTL_IP5_1|_RX|9  2.764e-12
L_PTL_IP5_1|_RX|1 _PTL_IP5_1|A_PTL _PTL_IP5_1|_RX|1  1.346e-12
L_PTL_IP5_1|_RX|2 _PTL_IP5_1|_RX|1 _PTL_IP5_1|_RX|4  6.348e-12
L_PTL_IP5_1|_RX|3 _PTL_IP5_1|_RX|4 _PTL_IP5_1|_RX|7  5.197e-12
L_PTL_IP5_1|_RX|4 _PTL_IP5_1|_RX|7 IP5_1_OUT  2.058e-12
L_PTL_IP5_1|_RX|P1 _PTL_IP5_1|_RX|2 0  4.795e-13
L_PTL_IP5_1|_RX|P2 _PTL_IP5_1|_RX|5 0  5.431e-13
L_PTL_IP5_1|_RX|P3 _PTL_IP5_1|_RX|8 0  5.339e-13
R_PTL_IP5_1|_RX|B1 _PTL_IP5_1|_RX|1 _PTL_IP5_1|_RX|101  4.225701121488
R_PTL_IP5_1|_RX|B2 _PTL_IP5_1|_RX|4 _PTL_IP5_1|_RX|104  3.429952209
R_PTL_IP5_1|_RX|B3 _PTL_IP5_1|_RX|7 _PTL_IP5_1|_RX|107  2.7439617672
L_PTL_IP5_1|_RX|RB1 _PTL_IP5_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP5_1|_RX|RB2 _PTL_IP5_1|_RX|104 0  1.937922998085e-12
L_PTL_IP5_1|_RX|RB3 _PTL_IP5_1|_RX|107 0  1.550338398468e-12
B_PTL_IP7_1|_TX|1 _PTL_IP7_1|_TX|1 _PTL_IP7_1|_TX|2 JJMIT AREA=2.5
B_PTL_IP7_1|_TX|2 _PTL_IP7_1|_TX|4 _PTL_IP7_1|_TX|5 JJMIT AREA=2.5
I_PTL_IP7_1|_TX|B1 0 _PTL_IP7_1|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP7_1|_TX|B2 0 _PTL_IP7_1|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_1|_TX|B1 _PTL_IP7_1|_TX|1 _PTL_IP7_1|_TX|3  1.684e-12
L_PTL_IP7_1|_TX|B2 _PTL_IP7_1|_TX|4 _PTL_IP7_1|_TX|6  3.596e-12
L_PTL_IP7_1|_TX|1 IP7_1_OUT_TX _PTL_IP7_1|_TX|1  2.063e-12
L_PTL_IP7_1|_TX|2 _PTL_IP7_1|_TX|1 _PTL_IP7_1|_TX|4  4.123e-12
L_PTL_IP7_1|_TX|3 _PTL_IP7_1|_TX|4 _PTL_IP7_1|_TX|7  2.193e-12
R_PTL_IP7_1|_TX|D _PTL_IP7_1|_TX|7 _PTL_IP7_1|A_PTL  1.36
L_PTL_IP7_1|_TX|P1 _PTL_IP7_1|_TX|2 0  5.254e-13
L_PTL_IP7_1|_TX|P2 _PTL_IP7_1|_TX|5 0  5.141e-13
R_PTL_IP7_1|_TX|B1 _PTL_IP7_1|_TX|1 _PTL_IP7_1|_TX|101  2.7439617672
R_PTL_IP7_1|_TX|B2 _PTL_IP7_1|_TX|4 _PTL_IP7_1|_TX|104  2.7439617672
L_PTL_IP7_1|_TX|RB1 _PTL_IP7_1|_TX|101 0  1.550338398468e-12
L_PTL_IP7_1|_TX|RB2 _PTL_IP7_1|_TX|104 0  1.550338398468e-12
B_PTL_IP7_1|_RX|1 _PTL_IP7_1|_RX|1 _PTL_IP7_1|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP7_1|_RX|2 _PTL_IP7_1|_RX|4 _PTL_IP7_1|_RX|5 JJMIT AREA=2.0
B_PTL_IP7_1|_RX|3 _PTL_IP7_1|_RX|7 _PTL_IP7_1|_RX|8 JJMIT AREA=2.5
I_PTL_IP7_1|_RX|B1 0 _PTL_IP7_1|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP7_1|_RX|B1 _PTL_IP7_1|_RX|1 _PTL_IP7_1|_RX|3  2.777e-12
I_PTL_IP7_1|_RX|B2 0 _PTL_IP7_1|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP7_1|_RX|B2 _PTL_IP7_1|_RX|4 _PTL_IP7_1|_RX|6  2.685e-12
I_PTL_IP7_1|_RX|B3 0 _PTL_IP7_1|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_1|_RX|B3 _PTL_IP7_1|_RX|7 _PTL_IP7_1|_RX|9  2.764e-12
L_PTL_IP7_1|_RX|1 _PTL_IP7_1|A_PTL _PTL_IP7_1|_RX|1  1.346e-12
L_PTL_IP7_1|_RX|2 _PTL_IP7_1|_RX|1 _PTL_IP7_1|_RX|4  6.348e-12
L_PTL_IP7_1|_RX|3 _PTL_IP7_1|_RX|4 _PTL_IP7_1|_RX|7  5.197e-12
L_PTL_IP7_1|_RX|4 _PTL_IP7_1|_RX|7 IP7_1_OUT  2.058e-12
L_PTL_IP7_1|_RX|P1 _PTL_IP7_1|_RX|2 0  4.795e-13
L_PTL_IP7_1|_RX|P2 _PTL_IP7_1|_RX|5 0  5.431e-13
L_PTL_IP7_1|_RX|P3 _PTL_IP7_1|_RX|8 0  5.339e-13
R_PTL_IP7_1|_RX|B1 _PTL_IP7_1|_RX|1 _PTL_IP7_1|_RX|101  4.225701121488
R_PTL_IP7_1|_RX|B2 _PTL_IP7_1|_RX|4 _PTL_IP7_1|_RX|104  3.429952209
R_PTL_IP7_1|_RX|B3 _PTL_IP7_1|_RX|7 _PTL_IP7_1|_RX|107  2.7439617672
L_PTL_IP7_1|_RX|RB1 _PTL_IP7_1|_RX|101 0  2.38752113364072e-12
L_PTL_IP7_1|_RX|RB2 _PTL_IP7_1|_RX|104 0  1.937922998085e-12
L_PTL_IP7_1|_RX|RB3 _PTL_IP7_1|_RX|107 0  1.550338398468e-12
L_S0_12|I_1|B _S0_12|A1 _S0_12|I_1|MID  2e-12
I_S0_12|I_1|B 0 _S0_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0_12|I_3|B _S0_12|A3 _S0_12|I_3|MID  2e-12
I_S0_12|I_3|B 0 _S0_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0_12|I_T|B _S0_12|T1 _S0_12|I_T|MID  2e-12
I_S0_12|I_T|B 0 _S0_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0_12|I_6|B _S0_12|Q1 _S0_12|I_6|MID  2e-12
I_S0_12|I_6|B 0 _S0_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0_12|1|1 _S0_12|A1 _S0_12|1|MID_SERIES JJMIT AREA=2.5
L_S0_12|1|P _S0_12|1|MID_SERIES 0  2e-13
R_S0_12|1|B _S0_12|A1 _S0_12|1|MID_SHUNT  2.7439617672
L_S0_12|1|RB _S0_12|1|MID_SHUNT 0  1.550338398468e-12
B_S0_12|23|1 _S0_12|A2 _S0_12|A3 JJMIT AREA=1.7857142857142858
R_S0_12|23|B _S0_12|A2 _S0_12|23|MID_SHUNT  3.84154647408
L_S0_12|23|RB _S0_12|23|MID_SHUNT _S0_12|A3  2.1704737578552e-12
B_S0_12|3|1 _S0_12|A3 _S0_12|3|MID_SERIES JJMIT AREA=2.5
L_S0_12|3|P _S0_12|3|MID_SERIES 0  2e-13
R_S0_12|3|B _S0_12|A3 _S0_12|3|MID_SHUNT  2.7439617672
L_S0_12|3|RB _S0_12|3|MID_SHUNT 0  1.550338398468e-12
B_S0_12|4|1 _S0_12|A4 _S0_12|4|MID_SERIES JJMIT AREA=2.5
L_S0_12|4|P _S0_12|4|MID_SERIES 0  2e-13
R_S0_12|4|B _S0_12|A4 _S0_12|4|MID_SHUNT  2.7439617672
L_S0_12|4|RB _S0_12|4|MID_SHUNT 0  1.550338398468e-12
B_S0_12|T|1 _S0_12|T1 _S0_12|T|MID_SERIES JJMIT AREA=2.5
L_S0_12|T|P _S0_12|T|MID_SERIES 0  2e-13
R_S0_12|T|B _S0_12|T1 _S0_12|T|MID_SHUNT  2.7439617672
L_S0_12|T|RB _S0_12|T|MID_SHUNT 0  1.550338398468e-12
B_S0_12|45|1 _S0_12|T2 _S0_12|A4 JJMIT AREA=1.7857142857142858
R_S0_12|45|B _S0_12|T2 _S0_12|45|MID_SHUNT  3.84154647408
L_S0_12|45|RB _S0_12|45|MID_SHUNT _S0_12|A4  2.1704737578552e-12
B_S0_12|6|1 _S0_12|Q1 _S0_12|6|MID_SERIES JJMIT AREA=2.5
L_S0_12|6|P _S0_12|6|MID_SERIES 0  2e-13
R_S0_12|6|B _S0_12|Q1 _S0_12|6|MID_SHUNT  2.7439617672
L_S0_12|6|RB _S0_12|6|MID_SHUNT 0  1.550338398468e-12
L_S1_12|I_1|B _S1_12|A1 _S1_12|I_1|MID  2e-12
I_S1_12|I_1|B 0 _S1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S1_12|I_3|B _S1_12|A3 _S1_12|I_3|MID  2e-12
I_S1_12|I_3|B 0 _S1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S1_12|I_T|B _S1_12|T1 _S1_12|I_T|MID  2e-12
I_S1_12|I_T|B 0 _S1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S1_12|I_6|B _S1_12|Q1 _S1_12|I_6|MID  2e-12
I_S1_12|I_6|B 0 _S1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S1_12|1|1 _S1_12|A1 _S1_12|1|MID_SERIES JJMIT AREA=2.5
L_S1_12|1|P _S1_12|1|MID_SERIES 0  2e-13
R_S1_12|1|B _S1_12|A1 _S1_12|1|MID_SHUNT  2.7439617672
L_S1_12|1|RB _S1_12|1|MID_SHUNT 0  1.550338398468e-12
B_S1_12|23|1 _S1_12|A2 _S1_12|A3 JJMIT AREA=1.7857142857142858
R_S1_12|23|B _S1_12|A2 _S1_12|23|MID_SHUNT  3.84154647408
L_S1_12|23|RB _S1_12|23|MID_SHUNT _S1_12|A3  2.1704737578552e-12
B_S1_12|3|1 _S1_12|A3 _S1_12|3|MID_SERIES JJMIT AREA=2.5
L_S1_12|3|P _S1_12|3|MID_SERIES 0  2e-13
R_S1_12|3|B _S1_12|A3 _S1_12|3|MID_SHUNT  2.7439617672
L_S1_12|3|RB _S1_12|3|MID_SHUNT 0  1.550338398468e-12
B_S1_12|4|1 _S1_12|A4 _S1_12|4|MID_SERIES JJMIT AREA=2.5
L_S1_12|4|P _S1_12|4|MID_SERIES 0  2e-13
R_S1_12|4|B _S1_12|A4 _S1_12|4|MID_SHUNT  2.7439617672
L_S1_12|4|RB _S1_12|4|MID_SHUNT 0  1.550338398468e-12
B_S1_12|T|1 _S1_12|T1 _S1_12|T|MID_SERIES JJMIT AREA=2.5
L_S1_12|T|P _S1_12|T|MID_SERIES 0  2e-13
R_S1_12|T|B _S1_12|T1 _S1_12|T|MID_SHUNT  2.7439617672
L_S1_12|T|RB _S1_12|T|MID_SHUNT 0  1.550338398468e-12
B_S1_12|45|1 _S1_12|T2 _S1_12|A4 JJMIT AREA=1.7857142857142858
R_S1_12|45|B _S1_12|T2 _S1_12|45|MID_SHUNT  3.84154647408
L_S1_12|45|RB _S1_12|45|MID_SHUNT _S1_12|A4  2.1704737578552e-12
B_S1_12|6|1 _S1_12|Q1 _S1_12|6|MID_SERIES JJMIT AREA=2.5
L_S1_12|6|P _S1_12|6|MID_SERIES 0  2e-13
R_S1_12|6|B _S1_12|Q1 _S1_12|6|MID_SHUNT  2.7439617672
L_S1_12|6|RB _S1_12|6|MID_SHUNT 0  1.550338398468e-12
L_S2_12|I_A1|B _S2_12|A1 _S2_12|I_A1|MID  2e-12
I_S2_12|I_A1|B 0 _S2_12|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S2_12|I_A3|B _S2_12|A3 _S2_12|I_A3|MID  2e-12
I_S2_12|I_A3|B 0 _S2_12|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S2_12|I_B1|B _S2_12|B1 _S2_12|I_B1|MID  2e-12
I_S2_12|I_B1|B 0 _S2_12|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S2_12|I_B3|B _S2_12|B3 _S2_12|I_B3|MID  2e-12
I_S2_12|I_B3|B 0 _S2_12|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S2_12|I_Q1|B _S2_12|Q1 _S2_12|I_Q1|MID  2e-12
I_S2_12|I_Q1|B 0 _S2_12|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S2_12|A1|1 _S2_12|A1 _S2_12|A1|MID_SERIES JJMIT AREA=2.5
L_S2_12|A1|P _S2_12|A1|MID_SERIES 0  5e-13
R_S2_12|A1|B _S2_12|A1 _S2_12|A1|MID_SHUNT  2.7439617672
L_S2_12|A1|RB _S2_12|A1|MID_SHUNT 0  2.050338398468e-12
B_S2_12|A2|1 _S2_12|A2 _S2_12|A2|MID_SERIES JJMIT AREA=2.5
L_S2_12|A2|P _S2_12|A2|MID_SERIES 0  5e-13
R_S2_12|A2|B _S2_12|A2 _S2_12|A2|MID_SHUNT  2.7439617672
L_S2_12|A2|RB _S2_12|A2|MID_SHUNT 0  2.050338398468e-12
B_S2_12|A3|1 _S2_12|A2 _S2_12|A3|MID_SERIES JJMIT AREA=2.5
L_S2_12|A3|P _S2_12|A3|MID_SERIES _S2_12|A3  1.2e-12
R_S2_12|A3|B _S2_12|A2 _S2_12|A3|MID_SHUNT  2.7439617672
L_S2_12|A3|RB _S2_12|A3|MID_SHUNT _S2_12|A3  2.050338398468e-12
B_S2_12|B1|1 _S2_12|B1 _S2_12|B1|MID_SERIES JJMIT AREA=2.5
L_S2_12|B1|P _S2_12|B1|MID_SERIES 0  5e-13
R_S2_12|B1|B _S2_12|B1 _S2_12|B1|MID_SHUNT  2.7439617672
L_S2_12|B1|RB _S2_12|B1|MID_SHUNT 0  2.050338398468e-12
B_S2_12|B2|1 _S2_12|B2 _S2_12|B2|MID_SERIES JJMIT AREA=2.5
L_S2_12|B2|P _S2_12|B2|MID_SERIES 0  5e-13
R_S2_12|B2|B _S2_12|B2 _S2_12|B2|MID_SHUNT  2.7439617672
L_S2_12|B2|RB _S2_12|B2|MID_SHUNT 0  2.050338398468e-12
B_S2_12|B3|1 _S2_12|B2 _S2_12|B3|MID_SERIES JJMIT AREA=2.5
L_S2_12|B3|P _S2_12|B3|MID_SERIES _S2_12|B3  1.2e-12
R_S2_12|B3|B _S2_12|B2 _S2_12|B3|MID_SHUNT  2.7439617672
L_S2_12|B3|RB _S2_12|B3|MID_SHUNT _S2_12|B3  2.050338398468e-12
B_S2_12|T1|1 _S2_12|T1 _S2_12|T1|MID_SERIES JJMIT AREA=2.5
L_S2_12|T1|P _S2_12|T1|MID_SERIES 0  5e-13
R_S2_12|T1|B _S2_12|T1 _S2_12|T1|MID_SHUNT  2.7439617672
L_S2_12|T1|RB _S2_12|T1|MID_SHUNT 0  2.050338398468e-12
B_S2_12|T2|1 _S2_12|T2 _S2_12|ABTQ JJMIT AREA=2.0
R_S2_12|T2|B _S2_12|T2 _S2_12|T2|MID_SHUNT  3.429952209
L_S2_12|T2|RB _S2_12|T2|MID_SHUNT _S2_12|ABTQ  2.437922998085e-12
B_S2_12|AB|1 _S2_12|AB _S2_12|AB|MID_SERIES JJMIT AREA=1.5
L_S2_12|AB|P _S2_12|AB|MID_SERIES _S2_12|ABTQ  1.2e-12
R_S2_12|AB|B _S2_12|AB _S2_12|AB|MID_SHUNT  4.573269612
L_S2_12|AB|RB _S2_12|AB|MID_SHUNT _S2_12|ABTQ  3.08389733078e-12
B_S2_12|ABTQ|1 _S2_12|ABTQ _S2_12|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S2_12|ABTQ|P _S2_12|ABTQ|MID_SERIES 0  5e-13
R_S2_12|ABTQ|B _S2_12|ABTQ _S2_12|ABTQ|MID_SHUNT  3.6586156896
L_S2_12|ABTQ|RB _S2_12|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S2_12|Q1|1 _S2_12|Q1 _S2_12|Q1|MID_SERIES JJMIT AREA=2.5
L_S2_12|Q1|P _S2_12|Q1|MID_SERIES 0  5e-13
R_S2_12|Q1|B _S2_12|Q1 _S2_12|Q1|MID_SHUNT  2.7439617672
L_S2_12|Q1|RB _S2_12|Q1|MID_SHUNT 0  2.050338398468e-12
L_PG2_12|_SPL_G1|1 G2_1_TO2 _PG2_12|_SPL_G1|D1  2e-12
L_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|D2  4.135667696e-12
L_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG2_12|_SPL_G1|5 _PG2_12|_SPL_G1|QA1 _PG2_12|G1_COPY_1  2e-12
L_PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|QB1 _PG2_12|G1_COPY_2  2e-12
L_PG2_12|_SPL_P1|1 P2_1_TO2 _PG2_12|_SPL_P1|D1  2e-12
L_PG2_12|_SPL_P1|2 _PG2_12|_SPL_P1|D1 _PG2_12|_SPL_P1|D2  4.135667696e-12
L_PG2_12|_SPL_P1|3 _PG2_12|_SPL_P1|D2 _PG2_12|_SPL_P1|JCT  9.84682784761905e-13
L_PG2_12|_SPL_P1|4 _PG2_12|_SPL_P1|JCT _PG2_12|_SPL_P1|QA1  9.84682784761905e-13
L_PG2_12|_SPL_P1|5 _PG2_12|_SPL_P1|QA1 _PG2_12|P1_COPY_1  2e-12
L_PG2_12|_SPL_P1|6 _PG2_12|_SPL_P1|JCT _PG2_12|_SPL_P1|QB1  9.84682784761905e-13
L_PG2_12|_SPL_P1|7 _PG2_12|_SPL_P1|QB1 _PG2_12|P1_COPY_2  2e-12
L_PG2_12|_PG|A1 _PG2_12|P1_COPY_1 _PG2_12|_PG|A1  2.067833848e-12
L_PG2_12|_PG|A2 _PG2_12|_PG|A1 _PG2_12|_PG|A2  4.135667696e-12
L_PG2_12|_PG|A3 _PG2_12|_PG|A3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|B1 _PG2_12|G1_COPY_1 _PG2_12|_PG|B1  2.067833848e-12
L_PG2_12|_PG|B2 _PG2_12|_PG|B1 _PG2_12|_PG|B2  4.135667696e-12
L_PG2_12|_PG|B3 _PG2_12|_PG|B3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|Q3 _PG2_12|_PG|Q3 _PG2_12|_PG|Q2  4.135667696e-12
L_PG2_12|_PG|Q2 _PG2_12|_PG|Q2 _PG2_12|_PG|Q1  4.135667696e-12
L_PG2_12|_PG|Q1 _PG2_12|_PG|Q1 _PG2_12|PG  2.067833848e-12
L_PG2_12|_GG|A1 G1_1_TO2 _PG2_12|_GG|A1  2.067833848e-12
L_PG2_12|_GG|A2 _PG2_12|_GG|A1 _PG2_12|_GG|A2  4.135667696e-12
L_PG2_12|_GG|A3 _PG2_12|_GG|A3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|B1 _PG2_12|G1_COPY_2 _PG2_12|_GG|B1  2.067833848e-12
L_PG2_12|_GG|B2 _PG2_12|_GG|B1 _PG2_12|_GG|B2  4.135667696e-12
L_PG2_12|_GG|B3 _PG2_12|_GG|B3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|Q3 _PG2_12|_GG|Q3 _PG2_12|_GG|Q2  4.135667696e-12
L_PG2_12|_GG|Q2 _PG2_12|_GG|Q2 _PG2_12|_GG|Q1  4.135667696e-12
L_PG2_12|_GG|Q1 _PG2_12|_GG|Q1 _PG2_12|GG  2.067833848e-12
L_PG2_12|_DFF_P0|1 P1_1_TO2 _PG2_12|_DFF_P0|A1  2.067833848e-12
L_PG2_12|_DFF_P0|2 _PG2_12|_DFF_P0|A1 _PG2_12|_DFF_P0|A2  4.135667696e-12
L_PG2_12|_DFF_P0|3 _PG2_12|_DFF_P0|A3 _PG2_12|_DFF_P0|A4  8.271335392e-12
L_PG2_12|_DFF_P0|T T23 _PG2_12|_DFF_P0|T1  2.067833848e-12
L_PG2_12|_DFF_P0|4 _PG2_12|_DFF_P0|T1 _PG2_12|_DFF_P0|T2  4.135667696e-12
L_PG2_12|_DFF_P0|5 _PG2_12|_DFF_P0|A4 _PG2_12|_DFF_P0|Q1  4.135667696e-12
L_PG2_12|_DFF_P0|6 _PG2_12|_DFF_P0|Q1 _PG2_12|P0_SYNC  2.067833848e-12
L_PG2_12|_DFF_P1|1 _PG2_12|P1_COPY_2 _PG2_12|_DFF_P1|A1  2.067833848e-12
L_PG2_12|_DFF_P1|2 _PG2_12|_DFF_P1|A1 _PG2_12|_DFF_P1|A2  4.135667696e-12
L_PG2_12|_DFF_P1|3 _PG2_12|_DFF_P1|A3 _PG2_12|_DFF_P1|A4  8.271335392e-12
L_PG2_12|_DFF_P1|T T23 _PG2_12|_DFF_P1|T1  2.067833848e-12
L_PG2_12|_DFF_P1|4 _PG2_12|_DFF_P1|T1 _PG2_12|_DFF_P1|T2  4.135667696e-12
L_PG2_12|_DFF_P1|5 _PG2_12|_DFF_P1|A4 _PG2_12|_DFF_P1|Q1  4.135667696e-12
L_PG2_12|_DFF_P1|6 _PG2_12|_DFF_P1|Q1 _PG2_12|P1_SYNC  2.067833848e-12
L_PG2_12|_DFF_PG|1 _PG2_12|PG _PG2_12|_DFF_PG|A1  2.067833848e-12
L_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|A2  4.135667696e-12
L_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|A4  8.271335392e-12
L_PG2_12|_DFF_PG|T T23 _PG2_12|_DFF_PG|T1  2.067833848e-12
L_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T2  4.135667696e-12
L_PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|Q1  4.135667696e-12
L_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|Q1 _PG2_12|PG_SYNC  2.067833848e-12
L_PG2_12|_DFF_GG|1 _PG2_12|GG _PG2_12|_DFF_GG|A1  2.067833848e-12
L_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|A2  4.135667696e-12
L_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|A4  8.271335392e-12
L_PG2_12|_DFF_GG|T T23 _PG2_12|_DFF_GG|T1  2.067833848e-12
L_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T2  4.135667696e-12
L_PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|Q1  4.135667696e-12
L_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|Q1 _PG2_12|GG_SYNC  2.067833848e-12
L_PG2_12|_AND_G|A1 _PG2_12|PG_SYNC _PG2_12|_AND_G|A1  2.067833848e-12
L_PG2_12|_AND_G|A2 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A2  4.135667696e-12
L_PG2_12|_AND_G|A3 _PG2_12|_AND_G|A3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|B1 _PG2_12|GG_SYNC _PG2_12|_AND_G|B1  2.067833848e-12
L_PG2_12|_AND_G|B2 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B2  4.135667696e-12
L_PG2_12|_AND_G|B3 _PG2_12|_AND_G|B3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q2  4.135667696e-12
L_PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q1  4.135667696e-12
L_PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1 G2_2_TX  2.067833848e-12
L_PG2_12|_AND_P|A1 _PG2_12|P0_SYNC _PG2_12|_AND_P|A1  2.067833848e-12
L_PG2_12|_AND_P|A2 _PG2_12|_AND_P|A1 _PG2_12|_AND_P|A2  4.135667696e-12
L_PG2_12|_AND_P|A3 _PG2_12|_AND_P|A3 _PG2_12|_AND_P|Q3  1.2e-12
L_PG2_12|_AND_P|B1 _PG2_12|P1_SYNC _PG2_12|_AND_P|B1  2.067833848e-12
L_PG2_12|_AND_P|B2 _PG2_12|_AND_P|B1 _PG2_12|_AND_P|B2  4.135667696e-12
L_PG2_12|_AND_P|B3 _PG2_12|_AND_P|B3 _PG2_12|_AND_P|Q3  1.2e-12
L_PG2_12|_AND_P|Q3 _PG2_12|_AND_P|Q3 _PG2_12|_AND_P|Q2  4.135667696e-12
L_PG2_12|_AND_P|Q2 _PG2_12|_AND_P|Q2 _PG2_12|_AND_P|Q1  4.135667696e-12
L_PG2_12|_AND_P|Q1 _PG2_12|_AND_P|Q1 P2_2_TX  2.067833848e-12
L_PG3_12|_SPL_G1|1 G3_1_TO3 _PG3_12|_SPL_G1|D1  2e-12
L_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|D2  4.135667696e-12
L_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_12|_SPL_G1|5 _PG3_12|_SPL_G1|QA1 _PG3_12|G1_COPY_1  2e-12
L_PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|QB1 _PG3_12|G1_COPY_2  2e-12
L_PG3_12|_SPL_P1|1 P3_1_TO3 _PG3_12|_SPL_P1|D1  2e-12
L_PG3_12|_SPL_P1|2 _PG3_12|_SPL_P1|D1 _PG3_12|_SPL_P1|D2  4.135667696e-12
L_PG3_12|_SPL_P1|3 _PG3_12|_SPL_P1|D2 _PG3_12|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_12|_SPL_P1|4 _PG3_12|_SPL_P1|JCT _PG3_12|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_12|_SPL_P1|5 _PG3_12|_SPL_P1|QA1 _PG3_12|P1_COPY_1  2e-12
L_PG3_12|_SPL_P1|6 _PG3_12|_SPL_P1|JCT _PG3_12|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_12|_SPL_P1|7 _PG3_12|_SPL_P1|QB1 _PG3_12|P1_COPY_2  2e-12
L_PG3_12|_PG|A1 _PG3_12|P1_COPY_1 _PG3_12|_PG|A1  2.067833848e-12
L_PG3_12|_PG|A2 _PG3_12|_PG|A1 _PG3_12|_PG|A2  4.135667696e-12
L_PG3_12|_PG|A3 _PG3_12|_PG|A3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|B1 _PG3_12|G1_COPY_1 _PG3_12|_PG|B1  2.067833848e-12
L_PG3_12|_PG|B2 _PG3_12|_PG|B1 _PG3_12|_PG|B2  4.135667696e-12
L_PG3_12|_PG|B3 _PG3_12|_PG|B3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|Q3 _PG3_12|_PG|Q3 _PG3_12|_PG|Q2  4.135667696e-12
L_PG3_12|_PG|Q2 _PG3_12|_PG|Q2 _PG3_12|_PG|Q1  4.135667696e-12
L_PG3_12|_PG|Q1 _PG3_12|_PG|Q1 _PG3_12|PG  2.067833848e-12
L_PG3_12|_GG|A1 G1_1_TO3 _PG3_12|_GG|A1  2.067833848e-12
L_PG3_12|_GG|A2 _PG3_12|_GG|A1 _PG3_12|_GG|A2  4.135667696e-12
L_PG3_12|_GG|A3 _PG3_12|_GG|A3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|B1 _PG3_12|G1_COPY_2 _PG3_12|_GG|B1  2.067833848e-12
L_PG3_12|_GG|B2 _PG3_12|_GG|B1 _PG3_12|_GG|B2  4.135667696e-12
L_PG3_12|_GG|B3 _PG3_12|_GG|B3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|Q3 _PG3_12|_GG|Q3 _PG3_12|_GG|Q2  4.135667696e-12
L_PG3_12|_GG|Q2 _PG3_12|_GG|Q2 _PG3_12|_GG|Q1  4.135667696e-12
L_PG3_12|_GG|Q1 _PG3_12|_GG|Q1 _PG3_12|GG  2.067833848e-12
L_PG3_12|_DFF_P0|1 P1_1_TO3 _PG3_12|_DFF_P0|A1  2.067833848e-12
L_PG3_12|_DFF_P0|2 _PG3_12|_DFF_P0|A1 _PG3_12|_DFF_P0|A2  4.135667696e-12
L_PG3_12|_DFF_P0|3 _PG3_12|_DFF_P0|A3 _PG3_12|_DFF_P0|A4  8.271335392e-12
L_PG3_12|_DFF_P0|T T24 _PG3_12|_DFF_P0|T1  2.067833848e-12
L_PG3_12|_DFF_P0|4 _PG3_12|_DFF_P0|T1 _PG3_12|_DFF_P0|T2  4.135667696e-12
L_PG3_12|_DFF_P0|5 _PG3_12|_DFF_P0|A4 _PG3_12|_DFF_P0|Q1  4.135667696e-12
L_PG3_12|_DFF_P0|6 _PG3_12|_DFF_P0|Q1 _PG3_12|P0_SYNC  2.067833848e-12
L_PG3_12|_DFF_P1|1 _PG3_12|P1_COPY_2 _PG3_12|_DFF_P1|A1  2.067833848e-12
L_PG3_12|_DFF_P1|2 _PG3_12|_DFF_P1|A1 _PG3_12|_DFF_P1|A2  4.135667696e-12
L_PG3_12|_DFF_P1|3 _PG3_12|_DFF_P1|A3 _PG3_12|_DFF_P1|A4  8.271335392e-12
L_PG3_12|_DFF_P1|T T24 _PG3_12|_DFF_P1|T1  2.067833848e-12
L_PG3_12|_DFF_P1|4 _PG3_12|_DFF_P1|T1 _PG3_12|_DFF_P1|T2  4.135667696e-12
L_PG3_12|_DFF_P1|5 _PG3_12|_DFF_P1|A4 _PG3_12|_DFF_P1|Q1  4.135667696e-12
L_PG3_12|_DFF_P1|6 _PG3_12|_DFF_P1|Q1 _PG3_12|P1_SYNC  2.067833848e-12
L_PG3_12|_DFF_PG|1 _PG3_12|PG _PG3_12|_DFF_PG|A1  2.067833848e-12
L_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|A2  4.135667696e-12
L_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|A4  8.271335392e-12
L_PG3_12|_DFF_PG|T T24 _PG3_12|_DFF_PG|T1  2.067833848e-12
L_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T2  4.135667696e-12
L_PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|Q1  4.135667696e-12
L_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|Q1 _PG3_12|PG_SYNC  2.067833848e-12
L_PG3_12|_DFF_GG|1 _PG3_12|GG _PG3_12|_DFF_GG|A1  2.067833848e-12
L_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|A2  4.135667696e-12
L_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|A4  8.271335392e-12
L_PG3_12|_DFF_GG|T T24 _PG3_12|_DFF_GG|T1  2.067833848e-12
L_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T2  4.135667696e-12
L_PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|Q1  4.135667696e-12
L_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|Q1 _PG3_12|GG_SYNC  2.067833848e-12
L_PG3_12|_AND_G|A1 _PG3_12|PG_SYNC _PG3_12|_AND_G|A1  2.067833848e-12
L_PG3_12|_AND_G|A2 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A2  4.135667696e-12
L_PG3_12|_AND_G|A3 _PG3_12|_AND_G|A3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|B1 _PG3_12|GG_SYNC _PG3_12|_AND_G|B1  2.067833848e-12
L_PG3_12|_AND_G|B2 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B2  4.135667696e-12
L_PG3_12|_AND_G|B3 _PG3_12|_AND_G|B3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q2  4.135667696e-12
L_PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q1  4.135667696e-12
L_PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1 G3_2_TX  2.067833848e-12
L_PG3_12|_AND_P|A1 _PG3_12|P0_SYNC _PG3_12|_AND_P|A1  2.067833848e-12
L_PG3_12|_AND_P|A2 _PG3_12|_AND_P|A1 _PG3_12|_AND_P|A2  4.135667696e-12
L_PG3_12|_AND_P|A3 _PG3_12|_AND_P|A3 _PG3_12|_AND_P|Q3  1.2e-12
L_PG3_12|_AND_P|B1 _PG3_12|P1_SYNC _PG3_12|_AND_P|B1  2.067833848e-12
L_PG3_12|_AND_P|B2 _PG3_12|_AND_P|B1 _PG3_12|_AND_P|B2  4.135667696e-12
L_PG3_12|_AND_P|B3 _PG3_12|_AND_P|B3 _PG3_12|_AND_P|Q3  1.2e-12
L_PG3_12|_AND_P|Q3 _PG3_12|_AND_P|Q3 _PG3_12|_AND_P|Q2  4.135667696e-12
L_PG3_12|_AND_P|Q2 _PG3_12|_AND_P|Q2 _PG3_12|_AND_P|Q1  4.135667696e-12
L_PG3_12|_AND_P|Q1 _PG3_12|_AND_P|Q1 P3_2_TX  2.067833848e-12
L_PG4_12|P|1 P4_1_TO4 _PG4_12|P|A1  2.067833848e-12
L_PG4_12|P|2 _PG4_12|P|A1 _PG4_12|P|A2  4.135667696e-12
L_PG4_12|P|3 _PG4_12|P|A3 _PG4_12|P|A4  8.271335392e-12
L_PG4_12|P|T T25 _PG4_12|P|T1  2.067833848e-12
L_PG4_12|P|4 _PG4_12|P|T1 _PG4_12|P|T2  4.135667696e-12
L_PG4_12|P|5 _PG4_12|P|A4 _PG4_12|P|Q1  4.135667696e-12
L_PG4_12|P|6 _PG4_12|P|Q1 P4_2_TX  2.067833848e-12
L_PG4_12|G|1 G4_1_TO4 _PG4_12|G|A1  2.067833848e-12
L_PG4_12|G|2 _PG4_12|G|A1 _PG4_12|G|A2  4.135667696e-12
L_PG4_12|G|3 _PG4_12|G|A3 _PG4_12|G|A4  8.271335392e-12
L_PG4_12|G|T T25 _PG4_12|G|T1  2.067833848e-12
L_PG4_12|G|4 _PG4_12|G|T1 _PG4_12|G|T2  4.135667696e-12
L_PG4_12|G|5 _PG4_12|G|A4 _PG4_12|G|Q1  4.135667696e-12
L_PG4_12|G|6 _PG4_12|G|Q1 G4_2_TX  2.067833848e-12
L_PG5_12|P|1 P5_1_TO5 _PG5_12|P|A1  2.067833848e-12
L_PG5_12|P|2 _PG5_12|P|A1 _PG5_12|P|A2  4.135667696e-12
L_PG5_12|P|3 _PG5_12|P|A3 _PG5_12|P|A4  8.271335392e-12
L_PG5_12|P|T T26 _PG5_12|P|T1  2.067833848e-12
L_PG5_12|P|4 _PG5_12|P|T1 _PG5_12|P|T2  4.135667696e-12
L_PG5_12|P|5 _PG5_12|P|A4 _PG5_12|P|Q1  4.135667696e-12
L_PG5_12|P|6 _PG5_12|P|Q1 P5_2_TX  2.067833848e-12
L_PG5_12|G|1 G5_1_TO5 _PG5_12|G|A1  2.067833848e-12
L_PG5_12|G|2 _PG5_12|G|A1 _PG5_12|G|A2  4.135667696e-12
L_PG5_12|G|3 _PG5_12|G|A3 _PG5_12|G|A4  8.271335392e-12
L_PG5_12|G|T T26 _PG5_12|G|T1  2.067833848e-12
L_PG5_12|G|4 _PG5_12|G|T1 _PG5_12|G|T2  4.135667696e-12
L_PG5_12|G|5 _PG5_12|G|A4 _PG5_12|G|Q1  4.135667696e-12
L_PG5_12|G|6 _PG5_12|G|Q1 G5_2_TX  2.067833848e-12
L_PG6_12|P|1 P6_1_TO6 _PG6_12|P|A1  2.067833848e-12
L_PG6_12|P|2 _PG6_12|P|A1 _PG6_12|P|A2  4.135667696e-12
L_PG6_12|P|3 _PG6_12|P|A3 _PG6_12|P|A4  8.271335392e-12
L_PG6_12|P|T T27 _PG6_12|P|T1  2.067833848e-12
L_PG6_12|P|4 _PG6_12|P|T1 _PG6_12|P|T2  4.135667696e-12
L_PG6_12|P|5 _PG6_12|P|A4 _PG6_12|P|Q1  4.135667696e-12
L_PG6_12|P|6 _PG6_12|P|Q1 P6_2_TX  2.067833848e-12
L_PG6_12|G|1 G6_1_TO6 _PG6_12|G|A1  2.067833848e-12
L_PG6_12|G|2 _PG6_12|G|A1 _PG6_12|G|A2  4.135667696e-12
L_PG6_12|G|3 _PG6_12|G|A3 _PG6_12|G|A4  8.271335392e-12
L_PG6_12|G|T T27 _PG6_12|G|T1  2.067833848e-12
L_PG6_12|G|4 _PG6_12|G|T1 _PG6_12|G|T2  4.135667696e-12
L_PG6_12|G|5 _PG6_12|G|A4 _PG6_12|G|Q1  4.135667696e-12
L_PG6_12|G|6 _PG6_12|G|Q1 G6_2_TX  2.067833848e-12
L_PG7_12|_SPL_G1|1 G7_1_TO7 _PG7_12|_SPL_G1|D1  2e-12
L_PG7_12|_SPL_G1|2 _PG7_12|_SPL_G1|D1 _PG7_12|_SPL_G1|D2  4.135667696e-12
L_PG7_12|_SPL_G1|3 _PG7_12|_SPL_G1|D2 _PG7_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG7_12|_SPL_G1|4 _PG7_12|_SPL_G1|JCT _PG7_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG7_12|_SPL_G1|5 _PG7_12|_SPL_G1|QA1 _PG7_12|G1_COPY_1  2e-12
L_PG7_12|_SPL_G1|6 _PG7_12|_SPL_G1|JCT _PG7_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG7_12|_SPL_G1|7 _PG7_12|_SPL_G1|QB1 _PG7_12|G1_COPY_2  2e-12
L_PG7_12|_SPL_P1|1 P7_1_TO7 _PG7_12|_SPL_P1|D1  2e-12
L_PG7_12|_SPL_P1|2 _PG7_12|_SPL_P1|D1 _PG7_12|_SPL_P1|D2  4.135667696e-12
L_PG7_12|_SPL_P1|3 _PG7_12|_SPL_P1|D2 _PG7_12|_SPL_P1|JCT  9.84682784761905e-13
L_PG7_12|_SPL_P1|4 _PG7_12|_SPL_P1|JCT _PG7_12|_SPL_P1|QA1  9.84682784761905e-13
L_PG7_12|_SPL_P1|5 _PG7_12|_SPL_P1|QA1 _PG7_12|P1_COPY_1  2e-12
L_PG7_12|_SPL_P1|6 _PG7_12|_SPL_P1|JCT _PG7_12|_SPL_P1|QB1  9.84682784761905e-13
L_PG7_12|_SPL_P1|7 _PG7_12|_SPL_P1|QB1 _PG7_12|P1_COPY_2  2e-12
L_PG7_12|_PG|A1 _PG7_12|P1_COPY_1 _PG7_12|_PG|A1  2.067833848e-12
L_PG7_12|_PG|A2 _PG7_12|_PG|A1 _PG7_12|_PG|A2  4.135667696e-12
L_PG7_12|_PG|A3 _PG7_12|_PG|A3 _PG7_12|_PG|Q3  1.2e-12
L_PG7_12|_PG|B1 _PG7_12|G1_COPY_1 _PG7_12|_PG|B1  2.067833848e-12
L_PG7_12|_PG|B2 _PG7_12|_PG|B1 _PG7_12|_PG|B2  4.135667696e-12
L_PG7_12|_PG|B3 _PG7_12|_PG|B3 _PG7_12|_PG|Q3  1.2e-12
L_PG7_12|_PG|Q3 _PG7_12|_PG|Q3 _PG7_12|_PG|Q2  4.135667696e-12
L_PG7_12|_PG|Q2 _PG7_12|_PG|Q2 _PG7_12|_PG|Q1  4.135667696e-12
L_PG7_12|_PG|Q1 _PG7_12|_PG|Q1 _PG7_12|PG  2.067833848e-12
L_PG7_12|_GG|A1 G5_1_TO7 _PG7_12|_GG|A1  2.067833848e-12
L_PG7_12|_GG|A2 _PG7_12|_GG|A1 _PG7_12|_GG|A2  4.135667696e-12
L_PG7_12|_GG|A3 _PG7_12|_GG|A3 _PG7_12|_GG|Q3  1.2e-12
L_PG7_12|_GG|B1 _PG7_12|G1_COPY_2 _PG7_12|_GG|B1  2.067833848e-12
L_PG7_12|_GG|B2 _PG7_12|_GG|B1 _PG7_12|_GG|B2  4.135667696e-12
L_PG7_12|_GG|B3 _PG7_12|_GG|B3 _PG7_12|_GG|Q3  1.2e-12
L_PG7_12|_GG|Q3 _PG7_12|_GG|Q3 _PG7_12|_GG|Q2  4.135667696e-12
L_PG7_12|_GG|Q2 _PG7_12|_GG|Q2 _PG7_12|_GG|Q1  4.135667696e-12
L_PG7_12|_GG|Q1 _PG7_12|_GG|Q1 _PG7_12|GG  2.067833848e-12
L_PG7_12|_DFF_P0|1 P5_1_TO7 _PG7_12|_DFF_P0|A1  2.067833848e-12
L_PG7_12|_DFF_P0|2 _PG7_12|_DFF_P0|A1 _PG7_12|_DFF_P0|A2  4.135667696e-12
L_PG7_12|_DFF_P0|3 _PG7_12|_DFF_P0|A3 _PG7_12|_DFF_P0|A4  8.271335392e-12
L_PG7_12|_DFF_P0|T T28 _PG7_12|_DFF_P0|T1  2.067833848e-12
L_PG7_12|_DFF_P0|4 _PG7_12|_DFF_P0|T1 _PG7_12|_DFF_P0|T2  4.135667696e-12
L_PG7_12|_DFF_P0|5 _PG7_12|_DFF_P0|A4 _PG7_12|_DFF_P0|Q1  4.135667696e-12
L_PG7_12|_DFF_P0|6 _PG7_12|_DFF_P0|Q1 _PG7_12|P0_SYNC  2.067833848e-12
L_PG7_12|_DFF_P1|1 _PG7_12|P1_COPY_2 _PG7_12|_DFF_P1|A1  2.067833848e-12
L_PG7_12|_DFF_P1|2 _PG7_12|_DFF_P1|A1 _PG7_12|_DFF_P1|A2  4.135667696e-12
L_PG7_12|_DFF_P1|3 _PG7_12|_DFF_P1|A3 _PG7_12|_DFF_P1|A4  8.271335392e-12
L_PG7_12|_DFF_P1|T T28 _PG7_12|_DFF_P1|T1  2.067833848e-12
L_PG7_12|_DFF_P1|4 _PG7_12|_DFF_P1|T1 _PG7_12|_DFF_P1|T2  4.135667696e-12
L_PG7_12|_DFF_P1|5 _PG7_12|_DFF_P1|A4 _PG7_12|_DFF_P1|Q1  4.135667696e-12
L_PG7_12|_DFF_P1|6 _PG7_12|_DFF_P1|Q1 _PG7_12|P1_SYNC  2.067833848e-12
L_PG7_12|_DFF_PG|1 _PG7_12|PG _PG7_12|_DFF_PG|A1  2.067833848e-12
L_PG7_12|_DFF_PG|2 _PG7_12|_DFF_PG|A1 _PG7_12|_DFF_PG|A2  4.135667696e-12
L_PG7_12|_DFF_PG|3 _PG7_12|_DFF_PG|A3 _PG7_12|_DFF_PG|A4  8.271335392e-12
L_PG7_12|_DFF_PG|T T28 _PG7_12|_DFF_PG|T1  2.067833848e-12
L_PG7_12|_DFF_PG|4 _PG7_12|_DFF_PG|T1 _PG7_12|_DFF_PG|T2  4.135667696e-12
L_PG7_12|_DFF_PG|5 _PG7_12|_DFF_PG|A4 _PG7_12|_DFF_PG|Q1  4.135667696e-12
L_PG7_12|_DFF_PG|6 _PG7_12|_DFF_PG|Q1 _PG7_12|PG_SYNC  2.067833848e-12
L_PG7_12|_DFF_GG|1 _PG7_12|GG _PG7_12|_DFF_GG|A1  2.067833848e-12
L_PG7_12|_DFF_GG|2 _PG7_12|_DFF_GG|A1 _PG7_12|_DFF_GG|A2  4.135667696e-12
L_PG7_12|_DFF_GG|3 _PG7_12|_DFF_GG|A3 _PG7_12|_DFF_GG|A4  8.271335392e-12
L_PG7_12|_DFF_GG|T T28 _PG7_12|_DFF_GG|T1  2.067833848e-12
L_PG7_12|_DFF_GG|4 _PG7_12|_DFF_GG|T1 _PG7_12|_DFF_GG|T2  4.135667696e-12
L_PG7_12|_DFF_GG|5 _PG7_12|_DFF_GG|A4 _PG7_12|_DFF_GG|Q1  4.135667696e-12
L_PG7_12|_DFF_GG|6 _PG7_12|_DFF_GG|Q1 _PG7_12|GG_SYNC  2.067833848e-12
L_PG7_12|_AND_G|A1 _PG7_12|PG_SYNC _PG7_12|_AND_G|A1  2.067833848e-12
L_PG7_12|_AND_G|A2 _PG7_12|_AND_G|A1 _PG7_12|_AND_G|A2  4.135667696e-12
L_PG7_12|_AND_G|A3 _PG7_12|_AND_G|A3 _PG7_12|_AND_G|Q3  1.2e-12
L_PG7_12|_AND_G|B1 _PG7_12|GG_SYNC _PG7_12|_AND_G|B1  2.067833848e-12
L_PG7_12|_AND_G|B2 _PG7_12|_AND_G|B1 _PG7_12|_AND_G|B2  4.135667696e-12
L_PG7_12|_AND_G|B3 _PG7_12|_AND_G|B3 _PG7_12|_AND_G|Q3  1.2e-12
L_PG7_12|_AND_G|Q3 _PG7_12|_AND_G|Q3 _PG7_12|_AND_G|Q2  4.135667696e-12
L_PG7_12|_AND_G|Q2 _PG7_12|_AND_G|Q2 _PG7_12|_AND_G|Q1  4.135667696e-12
L_PG7_12|_AND_G|Q1 _PG7_12|_AND_G|Q1 G7_2_TX  2.067833848e-12
L_PG7_12|_AND_P|A1 _PG7_12|P0_SYNC _PG7_12|_AND_P|A1  2.067833848e-12
L_PG7_12|_AND_P|A2 _PG7_12|_AND_P|A1 _PG7_12|_AND_P|A2  4.135667696e-12
L_PG7_12|_AND_P|A3 _PG7_12|_AND_P|A3 _PG7_12|_AND_P|Q3  1.2e-12
L_PG7_12|_AND_P|B1 _PG7_12|P1_SYNC _PG7_12|_AND_P|B1  2.067833848e-12
L_PG7_12|_AND_P|B2 _PG7_12|_AND_P|B1 _PG7_12|_AND_P|B2  4.135667696e-12
L_PG7_12|_AND_P|B3 _PG7_12|_AND_P|B3 _PG7_12|_AND_P|Q3  1.2e-12
L_PG7_12|_AND_P|Q3 _PG7_12|_AND_P|Q3 _PG7_12|_AND_P|Q2  4.135667696e-12
L_PG7_12|_AND_P|Q2 _PG7_12|_AND_P|Q2 _PG7_12|_AND_P|Q1  4.135667696e-12
L_PG7_12|_AND_P|Q1 _PG7_12|_AND_P|Q1 P7_2_TX  2.067833848e-12
L_IP3_12|I_1|B _IP3_12|A1 _IP3_12|I_1|MID  2e-12
I_IP3_12|I_1|B 0 _IP3_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP3_12|I_3|B _IP3_12|A3 _IP3_12|I_3|MID  2e-12
I_IP3_12|I_3|B 0 _IP3_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP3_12|I_T|B _IP3_12|T1 _IP3_12|I_T|MID  2e-12
I_IP3_12|I_T|B 0 _IP3_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP3_12|I_6|B _IP3_12|Q1 _IP3_12|I_6|MID  2e-12
I_IP3_12|I_6|B 0 _IP3_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP3_12|1|1 _IP3_12|A1 _IP3_12|1|MID_SERIES JJMIT AREA=2.5
L_IP3_12|1|P _IP3_12|1|MID_SERIES 0  2e-13
R_IP3_12|1|B _IP3_12|A1 _IP3_12|1|MID_SHUNT  2.7439617672
L_IP3_12|1|RB _IP3_12|1|MID_SHUNT 0  1.550338398468e-12
B_IP3_12|23|1 _IP3_12|A2 _IP3_12|A3 JJMIT AREA=1.7857142857142858
R_IP3_12|23|B _IP3_12|A2 _IP3_12|23|MID_SHUNT  3.84154647408
L_IP3_12|23|RB _IP3_12|23|MID_SHUNT _IP3_12|A3  2.1704737578552e-12
B_IP3_12|3|1 _IP3_12|A3 _IP3_12|3|MID_SERIES JJMIT AREA=2.5
L_IP3_12|3|P _IP3_12|3|MID_SERIES 0  2e-13
R_IP3_12|3|B _IP3_12|A3 _IP3_12|3|MID_SHUNT  2.7439617672
L_IP3_12|3|RB _IP3_12|3|MID_SHUNT 0  1.550338398468e-12
B_IP3_12|4|1 _IP3_12|A4 _IP3_12|4|MID_SERIES JJMIT AREA=2.5
L_IP3_12|4|P _IP3_12|4|MID_SERIES 0  2e-13
R_IP3_12|4|B _IP3_12|A4 _IP3_12|4|MID_SHUNT  2.7439617672
L_IP3_12|4|RB _IP3_12|4|MID_SHUNT 0  1.550338398468e-12
B_IP3_12|T|1 _IP3_12|T1 _IP3_12|T|MID_SERIES JJMIT AREA=2.5
L_IP3_12|T|P _IP3_12|T|MID_SERIES 0  2e-13
R_IP3_12|T|B _IP3_12|T1 _IP3_12|T|MID_SHUNT  2.7439617672
L_IP3_12|T|RB _IP3_12|T|MID_SHUNT 0  1.550338398468e-12
B_IP3_12|45|1 _IP3_12|T2 _IP3_12|A4 JJMIT AREA=1.7857142857142858
R_IP3_12|45|B _IP3_12|T2 _IP3_12|45|MID_SHUNT  3.84154647408
L_IP3_12|45|RB _IP3_12|45|MID_SHUNT _IP3_12|A4  2.1704737578552e-12
B_IP3_12|6|1 _IP3_12|Q1 _IP3_12|6|MID_SERIES JJMIT AREA=2.5
L_IP3_12|6|P _IP3_12|6|MID_SERIES 0  2e-13
R_IP3_12|6|B _IP3_12|Q1 _IP3_12|6|MID_SHUNT  2.7439617672
L_IP3_12|6|RB _IP3_12|6|MID_SHUNT 0  1.550338398468e-12
L_IP5_12|I_1|B _IP5_12|A1 _IP5_12|I_1|MID  2e-12
I_IP5_12|I_1|B 0 _IP5_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP5_12|I_3|B _IP5_12|A3 _IP5_12|I_3|MID  2e-12
I_IP5_12|I_3|B 0 _IP5_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP5_12|I_T|B _IP5_12|T1 _IP5_12|I_T|MID  2e-12
I_IP5_12|I_T|B 0 _IP5_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP5_12|I_6|B _IP5_12|Q1 _IP5_12|I_6|MID  2e-12
I_IP5_12|I_6|B 0 _IP5_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP5_12|1|1 _IP5_12|A1 _IP5_12|1|MID_SERIES JJMIT AREA=2.5
L_IP5_12|1|P _IP5_12|1|MID_SERIES 0  2e-13
R_IP5_12|1|B _IP5_12|A1 _IP5_12|1|MID_SHUNT  2.7439617672
L_IP5_12|1|RB _IP5_12|1|MID_SHUNT 0  1.550338398468e-12
B_IP5_12|23|1 _IP5_12|A2 _IP5_12|A3 JJMIT AREA=1.7857142857142858
R_IP5_12|23|B _IP5_12|A2 _IP5_12|23|MID_SHUNT  3.84154647408
L_IP5_12|23|RB _IP5_12|23|MID_SHUNT _IP5_12|A3  2.1704737578552e-12
B_IP5_12|3|1 _IP5_12|A3 _IP5_12|3|MID_SERIES JJMIT AREA=2.5
L_IP5_12|3|P _IP5_12|3|MID_SERIES 0  2e-13
R_IP5_12|3|B _IP5_12|A3 _IP5_12|3|MID_SHUNT  2.7439617672
L_IP5_12|3|RB _IP5_12|3|MID_SHUNT 0  1.550338398468e-12
B_IP5_12|4|1 _IP5_12|A4 _IP5_12|4|MID_SERIES JJMIT AREA=2.5
L_IP5_12|4|P _IP5_12|4|MID_SERIES 0  2e-13
R_IP5_12|4|B _IP5_12|A4 _IP5_12|4|MID_SHUNT  2.7439617672
L_IP5_12|4|RB _IP5_12|4|MID_SHUNT 0  1.550338398468e-12
B_IP5_12|T|1 _IP5_12|T1 _IP5_12|T|MID_SERIES JJMIT AREA=2.5
L_IP5_12|T|P _IP5_12|T|MID_SERIES 0  2e-13
R_IP5_12|T|B _IP5_12|T1 _IP5_12|T|MID_SHUNT  2.7439617672
L_IP5_12|T|RB _IP5_12|T|MID_SHUNT 0  1.550338398468e-12
B_IP5_12|45|1 _IP5_12|T2 _IP5_12|A4 JJMIT AREA=1.7857142857142858
R_IP5_12|45|B _IP5_12|T2 _IP5_12|45|MID_SHUNT  3.84154647408
L_IP5_12|45|RB _IP5_12|45|MID_SHUNT _IP5_12|A4  2.1704737578552e-12
B_IP5_12|6|1 _IP5_12|Q1 _IP5_12|6|MID_SERIES JJMIT AREA=2.5
L_IP5_12|6|P _IP5_12|6|MID_SERIES 0  2e-13
R_IP5_12|6|B _IP5_12|Q1 _IP5_12|6|MID_SHUNT  2.7439617672
L_IP5_12|6|RB _IP5_12|6|MID_SHUNT 0  1.550338398468e-12
L_IP7_12|I_1|B _IP7_12|A1 _IP7_12|I_1|MID  2e-12
I_IP7_12|I_1|B 0 _IP7_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP7_12|I_3|B _IP7_12|A3 _IP7_12|I_3|MID  2e-12
I_IP7_12|I_3|B 0 _IP7_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP7_12|I_T|B _IP7_12|T1 _IP7_12|I_T|MID  2e-12
I_IP7_12|I_T|B 0 _IP7_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP7_12|I_6|B _IP7_12|Q1 _IP7_12|I_6|MID  2e-12
I_IP7_12|I_6|B 0 _IP7_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP7_12|1|1 _IP7_12|A1 _IP7_12|1|MID_SERIES JJMIT AREA=2.5
L_IP7_12|1|P _IP7_12|1|MID_SERIES 0  2e-13
R_IP7_12|1|B _IP7_12|A1 _IP7_12|1|MID_SHUNT  2.7439617672
L_IP7_12|1|RB _IP7_12|1|MID_SHUNT 0  1.550338398468e-12
B_IP7_12|23|1 _IP7_12|A2 _IP7_12|A3 JJMIT AREA=1.7857142857142858
R_IP7_12|23|B _IP7_12|A2 _IP7_12|23|MID_SHUNT  3.84154647408
L_IP7_12|23|RB _IP7_12|23|MID_SHUNT _IP7_12|A3  2.1704737578552e-12
B_IP7_12|3|1 _IP7_12|A3 _IP7_12|3|MID_SERIES JJMIT AREA=2.5
L_IP7_12|3|P _IP7_12|3|MID_SERIES 0  2e-13
R_IP7_12|3|B _IP7_12|A3 _IP7_12|3|MID_SHUNT  2.7439617672
L_IP7_12|3|RB _IP7_12|3|MID_SHUNT 0  1.550338398468e-12
B_IP7_12|4|1 _IP7_12|A4 _IP7_12|4|MID_SERIES JJMIT AREA=2.5
L_IP7_12|4|P _IP7_12|4|MID_SERIES 0  2e-13
R_IP7_12|4|B _IP7_12|A4 _IP7_12|4|MID_SHUNT  2.7439617672
L_IP7_12|4|RB _IP7_12|4|MID_SHUNT 0  1.550338398468e-12
B_IP7_12|T|1 _IP7_12|T1 _IP7_12|T|MID_SERIES JJMIT AREA=2.5
L_IP7_12|T|P _IP7_12|T|MID_SERIES 0  2e-13
R_IP7_12|T|B _IP7_12|T1 _IP7_12|T|MID_SHUNT  2.7439617672
L_IP7_12|T|RB _IP7_12|T|MID_SHUNT 0  1.550338398468e-12
B_IP7_12|45|1 _IP7_12|T2 _IP7_12|A4 JJMIT AREA=1.7857142857142858
R_IP7_12|45|B _IP7_12|T2 _IP7_12|45|MID_SHUNT  3.84154647408
L_IP7_12|45|RB _IP7_12|45|MID_SHUNT _IP7_12|A4  2.1704737578552e-12
B_IP7_12|6|1 _IP7_12|Q1 _IP7_12|6|MID_SERIES JJMIT AREA=2.5
L_IP7_12|6|P _IP7_12|6|MID_SERIES 0  2e-13
R_IP7_12|6|B _IP7_12|Q1 _IP7_12|6|MID_SHUNT  2.7439617672
L_IP7_12|6|RB _IP7_12|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_S0_2|_TX|1 _PTL_S0_2|_TX|1 _PTL_S0_2|_TX|2 JJMIT AREA=2.5
B_PTL_S0_2|_TX|2 _PTL_S0_2|_TX|4 _PTL_S0_2|_TX|5 JJMIT AREA=2.5
I_PTL_S0_2|_TX|B1 0 _PTL_S0_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S0_2|_TX|B2 0 _PTL_S0_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S0_2|_TX|B1 _PTL_S0_2|_TX|1 _PTL_S0_2|_TX|3  1.684e-12
L_PTL_S0_2|_TX|B2 _PTL_S0_2|_TX|4 _PTL_S0_2|_TX|6  3.596e-12
L_PTL_S0_2|_TX|1 S0_2_TX _PTL_S0_2|_TX|1  2.063e-12
L_PTL_S0_2|_TX|2 _PTL_S0_2|_TX|1 _PTL_S0_2|_TX|4  4.123e-12
L_PTL_S0_2|_TX|3 _PTL_S0_2|_TX|4 _PTL_S0_2|_TX|7  2.193e-12
R_PTL_S0_2|_TX|D _PTL_S0_2|_TX|7 _PTL_S0_2|A_PTL  1.36
L_PTL_S0_2|_TX|P1 _PTL_S0_2|_TX|2 0  5.254e-13
L_PTL_S0_2|_TX|P2 _PTL_S0_2|_TX|5 0  5.141e-13
R_PTL_S0_2|_TX|B1 _PTL_S0_2|_TX|1 _PTL_S0_2|_TX|101  2.7439617672
R_PTL_S0_2|_TX|B2 _PTL_S0_2|_TX|4 _PTL_S0_2|_TX|104  2.7439617672
L_PTL_S0_2|_TX|RB1 _PTL_S0_2|_TX|101 0  1.550338398468e-12
L_PTL_S0_2|_TX|RB2 _PTL_S0_2|_TX|104 0  1.550338398468e-12
B_PTL_S0_2|_RX|1 _PTL_S0_2|_RX|1 _PTL_S0_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S0_2|_RX|2 _PTL_S0_2|_RX|4 _PTL_S0_2|_RX|5 JJMIT AREA=2.0
B_PTL_S0_2|_RX|3 _PTL_S0_2|_RX|7 _PTL_S0_2|_RX|8 JJMIT AREA=2.5
I_PTL_S0_2|_RX|B1 0 _PTL_S0_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S0_2|_RX|B1 _PTL_S0_2|_RX|1 _PTL_S0_2|_RX|3  2.777e-12
I_PTL_S0_2|_RX|B2 0 _PTL_S0_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S0_2|_RX|B2 _PTL_S0_2|_RX|4 _PTL_S0_2|_RX|6  2.685e-12
I_PTL_S0_2|_RX|B3 0 _PTL_S0_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S0_2|_RX|B3 _PTL_S0_2|_RX|7 _PTL_S0_2|_RX|9  2.764e-12
L_PTL_S0_2|_RX|1 _PTL_S0_2|A_PTL _PTL_S0_2|_RX|1  1.346e-12
L_PTL_S0_2|_RX|2 _PTL_S0_2|_RX|1 _PTL_S0_2|_RX|4  6.348e-12
L_PTL_S0_2|_RX|3 _PTL_S0_2|_RX|4 _PTL_S0_2|_RX|7  5.197e-12
L_PTL_S0_2|_RX|4 _PTL_S0_2|_RX|7 S0_2  2.058e-12
L_PTL_S0_2|_RX|P1 _PTL_S0_2|_RX|2 0  4.795e-13
L_PTL_S0_2|_RX|P2 _PTL_S0_2|_RX|5 0  5.431e-13
L_PTL_S0_2|_RX|P3 _PTL_S0_2|_RX|8 0  5.339e-13
R_PTL_S0_2|_RX|B1 _PTL_S0_2|_RX|1 _PTL_S0_2|_RX|101  4.225701121488
R_PTL_S0_2|_RX|B2 _PTL_S0_2|_RX|4 _PTL_S0_2|_RX|104  3.429952209
R_PTL_S0_2|_RX|B3 _PTL_S0_2|_RX|7 _PTL_S0_2|_RX|107  2.7439617672
L_PTL_S0_2|_RX|RB1 _PTL_S0_2|_RX|101 0  2.38752113364072e-12
L_PTL_S0_2|_RX|RB2 _PTL_S0_2|_RX|104 0  1.937922998085e-12
L_PTL_S0_2|_RX|RB3 _PTL_S0_2|_RX|107 0  1.550338398468e-12
B_PTL_S1_2|_TX|1 _PTL_S1_2|_TX|1 _PTL_S1_2|_TX|2 JJMIT AREA=2.5
B_PTL_S1_2|_TX|2 _PTL_S1_2|_TX|4 _PTL_S1_2|_TX|5 JJMIT AREA=2.5
I_PTL_S1_2|_TX|B1 0 _PTL_S1_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S1_2|_TX|B2 0 _PTL_S1_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S1_2|_TX|B1 _PTL_S1_2|_TX|1 _PTL_S1_2|_TX|3  1.684e-12
L_PTL_S1_2|_TX|B2 _PTL_S1_2|_TX|4 _PTL_S1_2|_TX|6  3.596e-12
L_PTL_S1_2|_TX|1 S1_2_TX _PTL_S1_2|_TX|1  2.063e-12
L_PTL_S1_2|_TX|2 _PTL_S1_2|_TX|1 _PTL_S1_2|_TX|4  4.123e-12
L_PTL_S1_2|_TX|3 _PTL_S1_2|_TX|4 _PTL_S1_2|_TX|7  2.193e-12
R_PTL_S1_2|_TX|D _PTL_S1_2|_TX|7 _PTL_S1_2|A_PTL  1.36
L_PTL_S1_2|_TX|P1 _PTL_S1_2|_TX|2 0  5.254e-13
L_PTL_S1_2|_TX|P2 _PTL_S1_2|_TX|5 0  5.141e-13
R_PTL_S1_2|_TX|B1 _PTL_S1_2|_TX|1 _PTL_S1_2|_TX|101  2.7439617672
R_PTL_S1_2|_TX|B2 _PTL_S1_2|_TX|4 _PTL_S1_2|_TX|104  2.7439617672
L_PTL_S1_2|_TX|RB1 _PTL_S1_2|_TX|101 0  1.550338398468e-12
L_PTL_S1_2|_TX|RB2 _PTL_S1_2|_TX|104 0  1.550338398468e-12
B_PTL_S1_2|_RX|1 _PTL_S1_2|_RX|1 _PTL_S1_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S1_2|_RX|2 _PTL_S1_2|_RX|4 _PTL_S1_2|_RX|5 JJMIT AREA=2.0
B_PTL_S1_2|_RX|3 _PTL_S1_2|_RX|7 _PTL_S1_2|_RX|8 JJMIT AREA=2.5
I_PTL_S1_2|_RX|B1 0 _PTL_S1_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S1_2|_RX|B1 _PTL_S1_2|_RX|1 _PTL_S1_2|_RX|3  2.777e-12
I_PTL_S1_2|_RX|B2 0 _PTL_S1_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S1_2|_RX|B2 _PTL_S1_2|_RX|4 _PTL_S1_2|_RX|6  2.685e-12
I_PTL_S1_2|_RX|B3 0 _PTL_S1_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S1_2|_RX|B3 _PTL_S1_2|_RX|7 _PTL_S1_2|_RX|9  2.764e-12
L_PTL_S1_2|_RX|1 _PTL_S1_2|A_PTL _PTL_S1_2|_RX|1  1.346e-12
L_PTL_S1_2|_RX|2 _PTL_S1_2|_RX|1 _PTL_S1_2|_RX|4  6.348e-12
L_PTL_S1_2|_RX|3 _PTL_S1_2|_RX|4 _PTL_S1_2|_RX|7  5.197e-12
L_PTL_S1_2|_RX|4 _PTL_S1_2|_RX|7 S1_2  2.058e-12
L_PTL_S1_2|_RX|P1 _PTL_S1_2|_RX|2 0  4.795e-13
L_PTL_S1_2|_RX|P2 _PTL_S1_2|_RX|5 0  5.431e-13
L_PTL_S1_2|_RX|P3 _PTL_S1_2|_RX|8 0  5.339e-13
R_PTL_S1_2|_RX|B1 _PTL_S1_2|_RX|1 _PTL_S1_2|_RX|101  4.225701121488
R_PTL_S1_2|_RX|B2 _PTL_S1_2|_RX|4 _PTL_S1_2|_RX|104  3.429952209
R_PTL_S1_2|_RX|B3 _PTL_S1_2|_RX|7 _PTL_S1_2|_RX|107  2.7439617672
L_PTL_S1_2|_RX|RB1 _PTL_S1_2|_RX|101 0  2.38752113364072e-12
L_PTL_S1_2|_RX|RB2 _PTL_S1_2|_RX|104 0  1.937922998085e-12
L_PTL_S1_2|_RX|RB3 _PTL_S1_2|_RX|107 0  1.550338398468e-12
B_PTL_S2_2|_TX|1 _PTL_S2_2|_TX|1 _PTL_S2_2|_TX|2 JJMIT AREA=2.5
B_PTL_S2_2|_TX|2 _PTL_S2_2|_TX|4 _PTL_S2_2|_TX|5 JJMIT AREA=2.5
I_PTL_S2_2|_TX|B1 0 _PTL_S2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S2_2|_TX|B2 0 _PTL_S2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S2_2|_TX|B1 _PTL_S2_2|_TX|1 _PTL_S2_2|_TX|3  1.684e-12
L_PTL_S2_2|_TX|B2 _PTL_S2_2|_TX|4 _PTL_S2_2|_TX|6  3.596e-12
L_PTL_S2_2|_TX|1 S2_2_TX _PTL_S2_2|_TX|1  2.063e-12
L_PTL_S2_2|_TX|2 _PTL_S2_2|_TX|1 _PTL_S2_2|_TX|4  4.123e-12
L_PTL_S2_2|_TX|3 _PTL_S2_2|_TX|4 _PTL_S2_2|_TX|7  2.193e-12
R_PTL_S2_2|_TX|D _PTL_S2_2|_TX|7 _PTL_S2_2|A_PTL  1.36
L_PTL_S2_2|_TX|P1 _PTL_S2_2|_TX|2 0  5.254e-13
L_PTL_S2_2|_TX|P2 _PTL_S2_2|_TX|5 0  5.141e-13
R_PTL_S2_2|_TX|B1 _PTL_S2_2|_TX|1 _PTL_S2_2|_TX|101  2.7439617672
R_PTL_S2_2|_TX|B2 _PTL_S2_2|_TX|4 _PTL_S2_2|_TX|104  2.7439617672
L_PTL_S2_2|_TX|RB1 _PTL_S2_2|_TX|101 0  1.550338398468e-12
L_PTL_S2_2|_TX|RB2 _PTL_S2_2|_TX|104 0  1.550338398468e-12
B_PTL_S2_2|_RX|1 _PTL_S2_2|_RX|1 _PTL_S2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S2_2|_RX|2 _PTL_S2_2|_RX|4 _PTL_S2_2|_RX|5 JJMIT AREA=2.0
B_PTL_S2_2|_RX|3 _PTL_S2_2|_RX|7 _PTL_S2_2|_RX|8 JJMIT AREA=2.5
I_PTL_S2_2|_RX|B1 0 _PTL_S2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S2_2|_RX|B1 _PTL_S2_2|_RX|1 _PTL_S2_2|_RX|3  2.777e-12
I_PTL_S2_2|_RX|B2 0 _PTL_S2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S2_2|_RX|B2 _PTL_S2_2|_RX|4 _PTL_S2_2|_RX|6  2.685e-12
I_PTL_S2_2|_RX|B3 0 _PTL_S2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S2_2|_RX|B3 _PTL_S2_2|_RX|7 _PTL_S2_2|_RX|9  2.764e-12
L_PTL_S2_2|_RX|1 _PTL_S2_2|A_PTL _PTL_S2_2|_RX|1  1.346e-12
L_PTL_S2_2|_RX|2 _PTL_S2_2|_RX|1 _PTL_S2_2|_RX|4  6.348e-12
L_PTL_S2_2|_RX|3 _PTL_S2_2|_RX|4 _PTL_S2_2|_RX|7  5.197e-12
L_PTL_S2_2|_RX|4 _PTL_S2_2|_RX|7 S2_2  2.058e-12
L_PTL_S2_2|_RX|P1 _PTL_S2_2|_RX|2 0  4.795e-13
L_PTL_S2_2|_RX|P2 _PTL_S2_2|_RX|5 0  5.431e-13
L_PTL_S2_2|_RX|P3 _PTL_S2_2|_RX|8 0  5.339e-13
R_PTL_S2_2|_RX|B1 _PTL_S2_2|_RX|1 _PTL_S2_2|_RX|101  4.225701121488
R_PTL_S2_2|_RX|B2 _PTL_S2_2|_RX|4 _PTL_S2_2|_RX|104  3.429952209
R_PTL_S2_2|_RX|B3 _PTL_S2_2|_RX|7 _PTL_S2_2|_RX|107  2.7439617672
L_PTL_S2_2|_RX|RB1 _PTL_S2_2|_RX|101 0  2.38752113364072e-12
L_PTL_S2_2|_RX|RB2 _PTL_S2_2|_RX|104 0  1.937922998085e-12
L_PTL_S2_2|_RX|RB3 _PTL_S2_2|_RX|107 0  1.550338398468e-12
B_PTL_G2_2|_TX|1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|2 JJMIT AREA=2.5
B_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|5 JJMIT AREA=2.5
I_PTL_G2_2|_TX|B1 0 _PTL_G2_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G2_2|_TX|B2 0 _PTL_G2_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|3  1.684e-12
L_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|6  3.596e-12
L_PTL_G2_2|_TX|1 G2_2_TX _PTL_G2_2|_TX|1  2.063e-12
L_PTL_G2_2|_TX|2 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|4  4.123e-12
L_PTL_G2_2|_TX|3 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|7  2.193e-12
R_PTL_G2_2|_TX|D _PTL_G2_2|_TX|7 _PTL_G2_2|A_PTL  1.36
L_PTL_G2_2|_TX|P1 _PTL_G2_2|_TX|2 0  5.254e-13
L_PTL_G2_2|_TX|P2 _PTL_G2_2|_TX|5 0  5.141e-13
R_PTL_G2_2|_TX|B1 _PTL_G2_2|_TX|1 _PTL_G2_2|_TX|101  2.7439617672
R_PTL_G2_2|_TX|B2 _PTL_G2_2|_TX|4 _PTL_G2_2|_TX|104  2.7439617672
L_PTL_G2_2|_TX|RB1 _PTL_G2_2|_TX|101 0  1.550338398468e-12
L_PTL_G2_2|_TX|RB2 _PTL_G2_2|_TX|104 0  1.550338398468e-12
B_PTL_G2_2|_RX|1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|5 JJMIT AREA=2.0
B_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|8 JJMIT AREA=2.5
I_PTL_G2_2|_RX|B1 0 _PTL_G2_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|3  2.777e-12
I_PTL_G2_2|_RX|B2 0 _PTL_G2_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|6  2.685e-12
I_PTL_G2_2|_RX|B3 0 _PTL_G2_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|9  2.764e-12
L_PTL_G2_2|_RX|1 _PTL_G2_2|A_PTL _PTL_G2_2|_RX|1  1.346e-12
L_PTL_G2_2|_RX|2 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|4  6.348e-12
L_PTL_G2_2|_RX|3 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7  5.197e-12
L_PTL_G2_2|_RX|4 _PTL_G2_2|_RX|7 G2_2_OUT  2.058e-12
L_PTL_G2_2|_RX|P1 _PTL_G2_2|_RX|2 0  4.795e-13
L_PTL_G2_2|_RX|P2 _PTL_G2_2|_RX|5 0  5.431e-13
L_PTL_G2_2|_RX|P3 _PTL_G2_2|_RX|8 0  5.339e-13
R_PTL_G2_2|_RX|B1 _PTL_G2_2|_RX|1 _PTL_G2_2|_RX|101  4.225701121488
R_PTL_G2_2|_RX|B2 _PTL_G2_2|_RX|4 _PTL_G2_2|_RX|104  3.429952209
R_PTL_G2_2|_RX|B3 _PTL_G2_2|_RX|7 _PTL_G2_2|_RX|107  2.7439617672
L_PTL_G2_2|_RX|RB1 _PTL_G2_2|_RX|101 0  2.38752113364072e-12
L_PTL_G2_2|_RX|RB2 _PTL_G2_2|_RX|104 0  1.937922998085e-12
L_PTL_G2_2|_RX|RB3 _PTL_G2_2|_RX|107 0  1.550338398468e-12
B_PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP3_2|_TX|B1 0 _PTL_IP3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP3_2|_TX|B2 0 _PTL_IP3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|3  1.684e-12
L_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|6  3.596e-12
L_PTL_IP3_2|_TX|1 IP3_2_OUT_TX _PTL_IP3_2|_TX|1  2.063e-12
L_PTL_IP3_2|_TX|2 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|4  4.123e-12
L_PTL_IP3_2|_TX|3 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|7  2.193e-12
R_PTL_IP3_2|_TX|D _PTL_IP3_2|_TX|7 _PTL_IP3_2|A_PTL  1.36
L_PTL_IP3_2|_TX|P1 _PTL_IP3_2|_TX|2 0  5.254e-13
L_PTL_IP3_2|_TX|P2 _PTL_IP3_2|_TX|5 0  5.141e-13
R_PTL_IP3_2|_TX|B1 _PTL_IP3_2|_TX|1 _PTL_IP3_2|_TX|101  2.7439617672
R_PTL_IP3_2|_TX|B2 _PTL_IP3_2|_TX|4 _PTL_IP3_2|_TX|104  2.7439617672
L_PTL_IP3_2|_TX|RB1 _PTL_IP3_2|_TX|101 0  1.550338398468e-12
L_PTL_IP3_2|_TX|RB2 _PTL_IP3_2|_TX|104 0  1.550338398468e-12
B_PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP3_2|_RX|B1 0 _PTL_IP3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|3  2.777e-12
I_PTL_IP3_2|_RX|B2 0 _PTL_IP3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|6  2.685e-12
I_PTL_IP3_2|_RX|B3 0 _PTL_IP3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|9  2.764e-12
L_PTL_IP3_2|_RX|1 _PTL_IP3_2|A_PTL _PTL_IP3_2|_RX|1  1.346e-12
L_PTL_IP3_2|_RX|2 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|4  6.348e-12
L_PTL_IP3_2|_RX|3 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7  5.197e-12
L_PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|7 IP3_2_OUT  2.058e-12
L_PTL_IP3_2|_RX|P1 _PTL_IP3_2|_RX|2 0  4.795e-13
L_PTL_IP3_2|_RX|P2 _PTL_IP3_2|_RX|5 0  5.431e-13
L_PTL_IP3_2|_RX|P3 _PTL_IP3_2|_RX|8 0  5.339e-13
R_PTL_IP3_2|_RX|B1 _PTL_IP3_2|_RX|1 _PTL_IP3_2|_RX|101  4.225701121488
R_PTL_IP3_2|_RX|B2 _PTL_IP3_2|_RX|4 _PTL_IP3_2|_RX|104  3.429952209
R_PTL_IP3_2|_RX|B3 _PTL_IP3_2|_RX|7 _PTL_IP3_2|_RX|107  2.7439617672
L_PTL_IP3_2|_RX|RB1 _PTL_IP3_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP3_2|_RX|RB2 _PTL_IP3_2|_RX|104 0  1.937922998085e-12
L_PTL_IP3_2|_RX|RB3 _PTL_IP3_2|_RX|107 0  1.550338398468e-12
B_PTL_P3_2|_TX|1 _PTL_P3_2|_TX|1 _PTL_P3_2|_TX|2 JJMIT AREA=2.5
B_PTL_P3_2|_TX|2 _PTL_P3_2|_TX|4 _PTL_P3_2|_TX|5 JJMIT AREA=2.5
I_PTL_P3_2|_TX|B1 0 _PTL_P3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P3_2|_TX|B2 0 _PTL_P3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P3_2|_TX|B1 _PTL_P3_2|_TX|1 _PTL_P3_2|_TX|3  1.684e-12
L_PTL_P3_2|_TX|B2 _PTL_P3_2|_TX|4 _PTL_P3_2|_TX|6  3.596e-12
L_PTL_P3_2|_TX|1 P3_2_TX _PTL_P3_2|_TX|1  2.063e-12
L_PTL_P3_2|_TX|2 _PTL_P3_2|_TX|1 _PTL_P3_2|_TX|4  4.123e-12
L_PTL_P3_2|_TX|3 _PTL_P3_2|_TX|4 _PTL_P3_2|_TX|7  2.193e-12
R_PTL_P3_2|_TX|D _PTL_P3_2|_TX|7 _PTL_P3_2|A_PTL  1.36
L_PTL_P3_2|_TX|P1 _PTL_P3_2|_TX|2 0  5.254e-13
L_PTL_P3_2|_TX|P2 _PTL_P3_2|_TX|5 0  5.141e-13
R_PTL_P3_2|_TX|B1 _PTL_P3_2|_TX|1 _PTL_P3_2|_TX|101  2.7439617672
R_PTL_P3_2|_TX|B2 _PTL_P3_2|_TX|4 _PTL_P3_2|_TX|104  2.7439617672
L_PTL_P3_2|_TX|RB1 _PTL_P3_2|_TX|101 0  1.550338398468e-12
L_PTL_P3_2|_TX|RB2 _PTL_P3_2|_TX|104 0  1.550338398468e-12
B_PTL_P3_2|_RX|1 _PTL_P3_2|_RX|1 _PTL_P3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P3_2|_RX|2 _PTL_P3_2|_RX|4 _PTL_P3_2|_RX|5 JJMIT AREA=2.0
B_PTL_P3_2|_RX|3 _PTL_P3_2|_RX|7 _PTL_P3_2|_RX|8 JJMIT AREA=2.5
I_PTL_P3_2|_RX|B1 0 _PTL_P3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P3_2|_RX|B1 _PTL_P3_2|_RX|1 _PTL_P3_2|_RX|3  2.777e-12
I_PTL_P3_2|_RX|B2 0 _PTL_P3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P3_2|_RX|B2 _PTL_P3_2|_RX|4 _PTL_P3_2|_RX|6  2.685e-12
I_PTL_P3_2|_RX|B3 0 _PTL_P3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P3_2|_RX|B3 _PTL_P3_2|_RX|7 _PTL_P3_2|_RX|9  2.764e-12
L_PTL_P3_2|_RX|1 _PTL_P3_2|A_PTL _PTL_P3_2|_RX|1  1.346e-12
L_PTL_P3_2|_RX|2 _PTL_P3_2|_RX|1 _PTL_P3_2|_RX|4  6.348e-12
L_PTL_P3_2|_RX|3 _PTL_P3_2|_RX|4 _PTL_P3_2|_RX|7  5.197e-12
L_PTL_P3_2|_RX|4 _PTL_P3_2|_RX|7 _PTL_P3_2|D  2.058e-12
L_PTL_P3_2|_RX|P1 _PTL_P3_2|_RX|2 0  4.795e-13
L_PTL_P3_2|_RX|P2 _PTL_P3_2|_RX|5 0  5.431e-13
L_PTL_P3_2|_RX|P3 _PTL_P3_2|_RX|8 0  5.339e-13
R_PTL_P3_2|_RX|B1 _PTL_P3_2|_RX|1 _PTL_P3_2|_RX|101  4.225701121488
R_PTL_P3_2|_RX|B2 _PTL_P3_2|_RX|4 _PTL_P3_2|_RX|104  3.429952209
R_PTL_P3_2|_RX|B3 _PTL_P3_2|_RX|7 _PTL_P3_2|_RX|107  2.7439617672
L_PTL_P3_2|_RX|RB1 _PTL_P3_2|_RX|101 0  2.38752113364072e-12
L_PTL_P3_2|_RX|RB2 _PTL_P3_2|_RX|104 0  1.937922998085e-12
L_PTL_P3_2|_RX|RB3 _PTL_P3_2|_RX|107 0  1.550338398468e-12
B_PTL_G3_2|_TX|1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|2 JJMIT AREA=2.5
B_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|5 JJMIT AREA=2.5
I_PTL_G3_2|_TX|B1 0 _PTL_G3_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G3_2|_TX|B2 0 _PTL_G3_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|3  1.684e-12
L_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|6  3.596e-12
L_PTL_G3_2|_TX|1 G3_2_TX _PTL_G3_2|_TX|1  2.063e-12
L_PTL_G3_2|_TX|2 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|4  4.123e-12
L_PTL_G3_2|_TX|3 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|7  2.193e-12
R_PTL_G3_2|_TX|D _PTL_G3_2|_TX|7 _PTL_G3_2|A_PTL  1.36
L_PTL_G3_2|_TX|P1 _PTL_G3_2|_TX|2 0  5.254e-13
L_PTL_G3_2|_TX|P2 _PTL_G3_2|_TX|5 0  5.141e-13
R_PTL_G3_2|_TX|B1 _PTL_G3_2|_TX|1 _PTL_G3_2|_TX|101  2.7439617672
R_PTL_G3_2|_TX|B2 _PTL_G3_2|_TX|4 _PTL_G3_2|_TX|104  2.7439617672
L_PTL_G3_2|_TX|RB1 _PTL_G3_2|_TX|101 0  1.550338398468e-12
L_PTL_G3_2|_TX|RB2 _PTL_G3_2|_TX|104 0  1.550338398468e-12
B_PTL_G3_2|_RX|1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|5 JJMIT AREA=2.0
B_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|8 JJMIT AREA=2.5
I_PTL_G3_2|_RX|B1 0 _PTL_G3_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|3  2.777e-12
I_PTL_G3_2|_RX|B2 0 _PTL_G3_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|6  2.685e-12
I_PTL_G3_2|_RX|B3 0 _PTL_G3_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|9  2.764e-12
L_PTL_G3_2|_RX|1 _PTL_G3_2|A_PTL _PTL_G3_2|_RX|1  1.346e-12
L_PTL_G3_2|_RX|2 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|4  6.348e-12
L_PTL_G3_2|_RX|3 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7  5.197e-12
L_PTL_G3_2|_RX|4 _PTL_G3_2|_RX|7 _PTL_G3_2|D  2.058e-12
L_PTL_G3_2|_RX|P1 _PTL_G3_2|_RX|2 0  4.795e-13
L_PTL_G3_2|_RX|P2 _PTL_G3_2|_RX|5 0  5.431e-13
L_PTL_G3_2|_RX|P3 _PTL_G3_2|_RX|8 0  5.339e-13
R_PTL_G3_2|_RX|B1 _PTL_G3_2|_RX|1 _PTL_G3_2|_RX|101  4.225701121488
R_PTL_G3_2|_RX|B2 _PTL_G3_2|_RX|4 _PTL_G3_2|_RX|104  3.429952209
R_PTL_G3_2|_RX|B3 _PTL_G3_2|_RX|7 _PTL_G3_2|_RX|107  2.7439617672
L_PTL_G3_2|_RX|RB1 _PTL_G3_2|_RX|101 0  2.38752113364072e-12
L_PTL_G3_2|_RX|RB2 _PTL_G3_2|_RX|104 0  1.937922998085e-12
L_PTL_G3_2|_RX|RB3 _PTL_G3_2|_RX|107 0  1.550338398468e-12
L_PTL_G3_2|_SPL_1|1 _PTL_G3_2|D _PTL_G3_2|_SPL_1|D1  2e-12
L_PTL_G3_2|_SPL_1|2 _PTL_G3_2|_SPL_1|D1 _PTL_G3_2|_SPL_1|D2  4.135667696e-12
L_PTL_G3_2|_SPL_1|3 _PTL_G3_2|_SPL_1|D2 _PTL_G3_2|_SPL_1|JCT  9.84682784761905e-13
L_PTL_G3_2|_SPL_1|4 _PTL_G3_2|_SPL_1|JCT _PTL_G3_2|_SPL_1|QA1  9.84682784761905e-13
L_PTL_G3_2|_SPL_1|5 _PTL_G3_2|_SPL_1|QA1 _PTL_G3_2|Q1  2e-12
L_PTL_G3_2|_SPL_1|6 _PTL_G3_2|_SPL_1|JCT _PTL_G3_2|_SPL_1|QB1  9.84682784761905e-13
L_PTL_G3_2|_SPL_1|7 _PTL_G3_2|_SPL_1|QB1 _PTL_G3_2|Q2  2e-12
L_PTL_G3_2|_SPL_2|1 _PTL_G3_2|Q1 _PTL_G3_2|_SPL_2|D1  2e-12
L_PTL_G3_2|_SPL_2|2 _PTL_G3_2|_SPL_2|D1 _PTL_G3_2|_SPL_2|D2  4.135667696e-12
L_PTL_G3_2|_SPL_2|3 _PTL_G3_2|_SPL_2|D2 _PTL_G3_2|_SPL_2|JCT  9.84682784761905e-13
L_PTL_G3_2|_SPL_2|4 _PTL_G3_2|_SPL_2|JCT _PTL_G3_2|_SPL_2|QA1  9.84682784761905e-13
L_PTL_G3_2|_SPL_2|5 _PTL_G3_2|_SPL_2|QA1 G3_2_TO4  2e-12
L_PTL_G3_2|_SPL_2|6 _PTL_G3_2|_SPL_2|JCT _PTL_G3_2|_SPL_2|QB1  9.84682784761905e-13
L_PTL_G3_2|_SPL_2|7 _PTL_G3_2|_SPL_2|QB1 G3_2_TO5  2e-12
L_PTL_G3_2|_SPL_3|1 _PTL_G3_2|Q2 _PTL_G3_2|_SPL_3|D1  2e-12
L_PTL_G3_2|_SPL_3|2 _PTL_G3_2|_SPL_3|D1 _PTL_G3_2|_SPL_3|D2  4.135667696e-12
L_PTL_G3_2|_SPL_3|3 _PTL_G3_2|_SPL_3|D2 _PTL_G3_2|_SPL_3|JCT  9.84682784761905e-13
L_PTL_G3_2|_SPL_3|4 _PTL_G3_2|_SPL_3|JCT _PTL_G3_2|_SPL_3|QA1  9.84682784761905e-13
L_PTL_G3_2|_SPL_3|5 _PTL_G3_2|_SPL_3|QA1 G3_2_TO7  2e-12
L_PTL_G3_2|_SPL_3|6 _PTL_G3_2|_SPL_3|JCT _PTL_G3_2|_SPL_3|QB1  9.84682784761905e-13
L_PTL_G3_2|_SPL_3|7 _PTL_G3_2|_SPL_3|QB1 G3_2_OUT  2e-12
B_PTL_P4_2|_TX|1 _PTL_P4_2|_TX|1 _PTL_P4_2|_TX|2 JJMIT AREA=2.5
B_PTL_P4_2|_TX|2 _PTL_P4_2|_TX|4 _PTL_P4_2|_TX|5 JJMIT AREA=2.5
I_PTL_P4_2|_TX|B1 0 _PTL_P4_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P4_2|_TX|B2 0 _PTL_P4_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P4_2|_TX|B1 _PTL_P4_2|_TX|1 _PTL_P4_2|_TX|3  1.684e-12
L_PTL_P4_2|_TX|B2 _PTL_P4_2|_TX|4 _PTL_P4_2|_TX|6  3.596e-12
L_PTL_P4_2|_TX|1 P4_2_TX _PTL_P4_2|_TX|1  2.063e-12
L_PTL_P4_2|_TX|2 _PTL_P4_2|_TX|1 _PTL_P4_2|_TX|4  4.123e-12
L_PTL_P4_2|_TX|3 _PTL_P4_2|_TX|4 _PTL_P4_2|_TX|7  2.193e-12
R_PTL_P4_2|_TX|D _PTL_P4_2|_TX|7 _PTL_P4_2|A_PTL  1.36
L_PTL_P4_2|_TX|P1 _PTL_P4_2|_TX|2 0  5.254e-13
L_PTL_P4_2|_TX|P2 _PTL_P4_2|_TX|5 0  5.141e-13
R_PTL_P4_2|_TX|B1 _PTL_P4_2|_TX|1 _PTL_P4_2|_TX|101  2.7439617672
R_PTL_P4_2|_TX|B2 _PTL_P4_2|_TX|4 _PTL_P4_2|_TX|104  2.7439617672
L_PTL_P4_2|_TX|RB1 _PTL_P4_2|_TX|101 0  1.550338398468e-12
L_PTL_P4_2|_TX|RB2 _PTL_P4_2|_TX|104 0  1.550338398468e-12
B_PTL_P4_2|_RX|1 _PTL_P4_2|_RX|1 _PTL_P4_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P4_2|_RX|2 _PTL_P4_2|_RX|4 _PTL_P4_2|_RX|5 JJMIT AREA=2.0
B_PTL_P4_2|_RX|3 _PTL_P4_2|_RX|7 _PTL_P4_2|_RX|8 JJMIT AREA=2.5
I_PTL_P4_2|_RX|B1 0 _PTL_P4_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P4_2|_RX|B1 _PTL_P4_2|_RX|1 _PTL_P4_2|_RX|3  2.777e-12
I_PTL_P4_2|_RX|B2 0 _PTL_P4_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P4_2|_RX|B2 _PTL_P4_2|_RX|4 _PTL_P4_2|_RX|6  2.685e-12
I_PTL_P4_2|_RX|B3 0 _PTL_P4_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P4_2|_RX|B3 _PTL_P4_2|_RX|7 _PTL_P4_2|_RX|9  2.764e-12
L_PTL_P4_2|_RX|1 _PTL_P4_2|A_PTL _PTL_P4_2|_RX|1  1.346e-12
L_PTL_P4_2|_RX|2 _PTL_P4_2|_RX|1 _PTL_P4_2|_RX|4  6.348e-12
L_PTL_P4_2|_RX|3 _PTL_P4_2|_RX|4 _PTL_P4_2|_RX|7  5.197e-12
L_PTL_P4_2|_RX|4 _PTL_P4_2|_RX|7 _PTL_P4_2|D  2.058e-12
L_PTL_P4_2|_RX|P1 _PTL_P4_2|_RX|2 0  4.795e-13
L_PTL_P4_2|_RX|P2 _PTL_P4_2|_RX|5 0  5.431e-13
L_PTL_P4_2|_RX|P3 _PTL_P4_2|_RX|8 0  5.339e-13
R_PTL_P4_2|_RX|B1 _PTL_P4_2|_RX|1 _PTL_P4_2|_RX|101  4.225701121488
R_PTL_P4_2|_RX|B2 _PTL_P4_2|_RX|4 _PTL_P4_2|_RX|104  3.429952209
R_PTL_P4_2|_RX|B3 _PTL_P4_2|_RX|7 _PTL_P4_2|_RX|107  2.7439617672
L_PTL_P4_2|_RX|RB1 _PTL_P4_2|_RX|101 0  2.38752113364072e-12
L_PTL_P4_2|_RX|RB2 _PTL_P4_2|_RX|104 0  1.937922998085e-12
L_PTL_P4_2|_RX|RB3 _PTL_P4_2|_RX|107 0  1.550338398468e-12
L_PTL_P4_2|_SPL|1 _PTL_P4_2|D _PTL_P4_2|_SPL|D1  2e-12
L_PTL_P4_2|_SPL|2 _PTL_P4_2|_SPL|D1 _PTL_P4_2|_SPL|D2  4.135667696e-12
L_PTL_P4_2|_SPL|3 _PTL_P4_2|_SPL|D2 _PTL_P4_2|_SPL|JCT  9.84682784761905e-13
L_PTL_P4_2|_SPL|4 _PTL_P4_2|_SPL|JCT _PTL_P4_2|_SPL|QA1  9.84682784761905e-13
L_PTL_P4_2|_SPL|5 _PTL_P4_2|_SPL|QA1 P4_2_TO4  2e-12
L_PTL_P4_2|_SPL|6 _PTL_P4_2|_SPL|JCT _PTL_P4_2|_SPL|QB1  9.84682784761905e-13
L_PTL_P4_2|_SPL|7 _PTL_P4_2|_SPL|QB1 P4_2_OUT  2e-12
B_PTL_G4_2|_TX|1 _PTL_G4_2|_TX|1 _PTL_G4_2|_TX|2 JJMIT AREA=2.5
B_PTL_G4_2|_TX|2 _PTL_G4_2|_TX|4 _PTL_G4_2|_TX|5 JJMIT AREA=2.5
I_PTL_G4_2|_TX|B1 0 _PTL_G4_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G4_2|_TX|B2 0 _PTL_G4_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G4_2|_TX|B1 _PTL_G4_2|_TX|1 _PTL_G4_2|_TX|3  1.684e-12
L_PTL_G4_2|_TX|B2 _PTL_G4_2|_TX|4 _PTL_G4_2|_TX|6  3.596e-12
L_PTL_G4_2|_TX|1 G4_2_TX _PTL_G4_2|_TX|1  2.063e-12
L_PTL_G4_2|_TX|2 _PTL_G4_2|_TX|1 _PTL_G4_2|_TX|4  4.123e-12
L_PTL_G4_2|_TX|3 _PTL_G4_2|_TX|4 _PTL_G4_2|_TX|7  2.193e-12
R_PTL_G4_2|_TX|D _PTL_G4_2|_TX|7 _PTL_G4_2|A_PTL  1.36
L_PTL_G4_2|_TX|P1 _PTL_G4_2|_TX|2 0  5.254e-13
L_PTL_G4_2|_TX|P2 _PTL_G4_2|_TX|5 0  5.141e-13
R_PTL_G4_2|_TX|B1 _PTL_G4_2|_TX|1 _PTL_G4_2|_TX|101  2.7439617672
R_PTL_G4_2|_TX|B2 _PTL_G4_2|_TX|4 _PTL_G4_2|_TX|104  2.7439617672
L_PTL_G4_2|_TX|RB1 _PTL_G4_2|_TX|101 0  1.550338398468e-12
L_PTL_G4_2|_TX|RB2 _PTL_G4_2|_TX|104 0  1.550338398468e-12
B_PTL_G4_2|_RX|1 _PTL_G4_2|_RX|1 _PTL_G4_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G4_2|_RX|2 _PTL_G4_2|_RX|4 _PTL_G4_2|_RX|5 JJMIT AREA=2.0
B_PTL_G4_2|_RX|3 _PTL_G4_2|_RX|7 _PTL_G4_2|_RX|8 JJMIT AREA=2.5
I_PTL_G4_2|_RX|B1 0 _PTL_G4_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G4_2|_RX|B1 _PTL_G4_2|_RX|1 _PTL_G4_2|_RX|3  2.777e-12
I_PTL_G4_2|_RX|B2 0 _PTL_G4_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G4_2|_RX|B2 _PTL_G4_2|_RX|4 _PTL_G4_2|_RX|6  2.685e-12
I_PTL_G4_2|_RX|B3 0 _PTL_G4_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G4_2|_RX|B3 _PTL_G4_2|_RX|7 _PTL_G4_2|_RX|9  2.764e-12
L_PTL_G4_2|_RX|1 _PTL_G4_2|A_PTL _PTL_G4_2|_RX|1  1.346e-12
L_PTL_G4_2|_RX|2 _PTL_G4_2|_RX|1 _PTL_G4_2|_RX|4  6.348e-12
L_PTL_G4_2|_RX|3 _PTL_G4_2|_RX|4 _PTL_G4_2|_RX|7  5.197e-12
L_PTL_G4_2|_RX|4 _PTL_G4_2|_RX|7 G4_2_TO4  2.058e-12
L_PTL_G4_2|_RX|P1 _PTL_G4_2|_RX|2 0  4.795e-13
L_PTL_G4_2|_RX|P2 _PTL_G4_2|_RX|5 0  5.431e-13
L_PTL_G4_2|_RX|P3 _PTL_G4_2|_RX|8 0  5.339e-13
R_PTL_G4_2|_RX|B1 _PTL_G4_2|_RX|1 _PTL_G4_2|_RX|101  4.225701121488
R_PTL_G4_2|_RX|B2 _PTL_G4_2|_RX|4 _PTL_G4_2|_RX|104  3.429952209
R_PTL_G4_2|_RX|B3 _PTL_G4_2|_RX|7 _PTL_G4_2|_RX|107  2.7439617672
L_PTL_G4_2|_RX|RB1 _PTL_G4_2|_RX|101 0  2.38752113364072e-12
L_PTL_G4_2|_RX|RB2 _PTL_G4_2|_RX|104 0  1.937922998085e-12
L_PTL_G4_2|_RX|RB3 _PTL_G4_2|_RX|107 0  1.550338398468e-12
B_PTL_IP5_2|_TX|1 _PTL_IP5_2|_TX|1 _PTL_IP5_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP5_2|_TX|2 _PTL_IP5_2|_TX|4 _PTL_IP5_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP5_2|_TX|B1 0 _PTL_IP5_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP5_2|_TX|B2 0 _PTL_IP5_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_2|_TX|B1 _PTL_IP5_2|_TX|1 _PTL_IP5_2|_TX|3  1.684e-12
L_PTL_IP5_2|_TX|B2 _PTL_IP5_2|_TX|4 _PTL_IP5_2|_TX|6  3.596e-12
L_PTL_IP5_2|_TX|1 IP5_2_OUT_TX _PTL_IP5_2|_TX|1  2.063e-12
L_PTL_IP5_2|_TX|2 _PTL_IP5_2|_TX|1 _PTL_IP5_2|_TX|4  4.123e-12
L_PTL_IP5_2|_TX|3 _PTL_IP5_2|_TX|4 _PTL_IP5_2|_TX|7  2.193e-12
R_PTL_IP5_2|_TX|D _PTL_IP5_2|_TX|7 _PTL_IP5_2|A_PTL  1.36
L_PTL_IP5_2|_TX|P1 _PTL_IP5_2|_TX|2 0  5.254e-13
L_PTL_IP5_2|_TX|P2 _PTL_IP5_2|_TX|5 0  5.141e-13
R_PTL_IP5_2|_TX|B1 _PTL_IP5_2|_TX|1 _PTL_IP5_2|_TX|101  2.7439617672
R_PTL_IP5_2|_TX|B2 _PTL_IP5_2|_TX|4 _PTL_IP5_2|_TX|104  2.7439617672
L_PTL_IP5_2|_TX|RB1 _PTL_IP5_2|_TX|101 0  1.550338398468e-12
L_PTL_IP5_2|_TX|RB2 _PTL_IP5_2|_TX|104 0  1.550338398468e-12
B_PTL_IP5_2|_RX|1 _PTL_IP5_2|_RX|1 _PTL_IP5_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP5_2|_RX|2 _PTL_IP5_2|_RX|4 _PTL_IP5_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP5_2|_RX|3 _PTL_IP5_2|_RX|7 _PTL_IP5_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP5_2|_RX|B1 0 _PTL_IP5_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP5_2|_RX|B1 _PTL_IP5_2|_RX|1 _PTL_IP5_2|_RX|3  2.777e-12
I_PTL_IP5_2|_RX|B2 0 _PTL_IP5_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP5_2|_RX|B2 _PTL_IP5_2|_RX|4 _PTL_IP5_2|_RX|6  2.685e-12
I_PTL_IP5_2|_RX|B3 0 _PTL_IP5_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_2|_RX|B3 _PTL_IP5_2|_RX|7 _PTL_IP5_2|_RX|9  2.764e-12
L_PTL_IP5_2|_RX|1 _PTL_IP5_2|A_PTL _PTL_IP5_2|_RX|1  1.346e-12
L_PTL_IP5_2|_RX|2 _PTL_IP5_2|_RX|1 _PTL_IP5_2|_RX|4  6.348e-12
L_PTL_IP5_2|_RX|3 _PTL_IP5_2|_RX|4 _PTL_IP5_2|_RX|7  5.197e-12
L_PTL_IP5_2|_RX|4 _PTL_IP5_2|_RX|7 IP5_2_OUT  2.058e-12
L_PTL_IP5_2|_RX|P1 _PTL_IP5_2|_RX|2 0  4.795e-13
L_PTL_IP5_2|_RX|P2 _PTL_IP5_2|_RX|5 0  5.431e-13
L_PTL_IP5_2|_RX|P3 _PTL_IP5_2|_RX|8 0  5.339e-13
R_PTL_IP5_2|_RX|B1 _PTL_IP5_2|_RX|1 _PTL_IP5_2|_RX|101  4.225701121488
R_PTL_IP5_2|_RX|B2 _PTL_IP5_2|_RX|4 _PTL_IP5_2|_RX|104  3.429952209
R_PTL_IP5_2|_RX|B3 _PTL_IP5_2|_RX|7 _PTL_IP5_2|_RX|107  2.7439617672
L_PTL_IP5_2|_RX|RB1 _PTL_IP5_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP5_2|_RX|RB2 _PTL_IP5_2|_RX|104 0  1.937922998085e-12
L_PTL_IP5_2|_RX|RB3 _PTL_IP5_2|_RX|107 0  1.550338398468e-12
B_PTL_P5_2|_TX|1 _PTL_P5_2|_TX|1 _PTL_P5_2|_TX|2 JJMIT AREA=2.5
B_PTL_P5_2|_TX|2 _PTL_P5_2|_TX|4 _PTL_P5_2|_TX|5 JJMIT AREA=2.5
I_PTL_P5_2|_TX|B1 0 _PTL_P5_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P5_2|_TX|B2 0 _PTL_P5_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P5_2|_TX|B1 _PTL_P5_2|_TX|1 _PTL_P5_2|_TX|3  1.684e-12
L_PTL_P5_2|_TX|B2 _PTL_P5_2|_TX|4 _PTL_P5_2|_TX|6  3.596e-12
L_PTL_P5_2|_TX|1 P5_2_TX _PTL_P5_2|_TX|1  2.063e-12
L_PTL_P5_2|_TX|2 _PTL_P5_2|_TX|1 _PTL_P5_2|_TX|4  4.123e-12
L_PTL_P5_2|_TX|3 _PTL_P5_2|_TX|4 _PTL_P5_2|_TX|7  2.193e-12
R_PTL_P5_2|_TX|D _PTL_P5_2|_TX|7 _PTL_P5_2|A_PTL  1.36
L_PTL_P5_2|_TX|P1 _PTL_P5_2|_TX|2 0  5.254e-13
L_PTL_P5_2|_TX|P2 _PTL_P5_2|_TX|5 0  5.141e-13
R_PTL_P5_2|_TX|B1 _PTL_P5_2|_TX|1 _PTL_P5_2|_TX|101  2.7439617672
R_PTL_P5_2|_TX|B2 _PTL_P5_2|_TX|4 _PTL_P5_2|_TX|104  2.7439617672
L_PTL_P5_2|_TX|RB1 _PTL_P5_2|_TX|101 0  1.550338398468e-12
L_PTL_P5_2|_TX|RB2 _PTL_P5_2|_TX|104 0  1.550338398468e-12
B_PTL_P5_2|_RX|1 _PTL_P5_2|_RX|1 _PTL_P5_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P5_2|_RX|2 _PTL_P5_2|_RX|4 _PTL_P5_2|_RX|5 JJMIT AREA=2.0
B_PTL_P5_2|_RX|3 _PTL_P5_2|_RX|7 _PTL_P5_2|_RX|8 JJMIT AREA=2.5
I_PTL_P5_2|_RX|B1 0 _PTL_P5_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P5_2|_RX|B1 _PTL_P5_2|_RX|1 _PTL_P5_2|_RX|3  2.777e-12
I_PTL_P5_2|_RX|B2 0 _PTL_P5_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P5_2|_RX|B2 _PTL_P5_2|_RX|4 _PTL_P5_2|_RX|6  2.685e-12
I_PTL_P5_2|_RX|B3 0 _PTL_P5_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P5_2|_RX|B3 _PTL_P5_2|_RX|7 _PTL_P5_2|_RX|9  2.764e-12
L_PTL_P5_2|_RX|1 _PTL_P5_2|A_PTL _PTL_P5_2|_RX|1  1.346e-12
L_PTL_P5_2|_RX|2 _PTL_P5_2|_RX|1 _PTL_P5_2|_RX|4  6.348e-12
L_PTL_P5_2|_RX|3 _PTL_P5_2|_RX|4 _PTL_P5_2|_RX|7  5.197e-12
L_PTL_P5_2|_RX|4 _PTL_P5_2|_RX|7 P5_2_TO5  2.058e-12
L_PTL_P5_2|_RX|P1 _PTL_P5_2|_RX|2 0  4.795e-13
L_PTL_P5_2|_RX|P2 _PTL_P5_2|_RX|5 0  5.431e-13
L_PTL_P5_2|_RX|P3 _PTL_P5_2|_RX|8 0  5.339e-13
R_PTL_P5_2|_RX|B1 _PTL_P5_2|_RX|1 _PTL_P5_2|_RX|101  4.225701121488
R_PTL_P5_2|_RX|B2 _PTL_P5_2|_RX|4 _PTL_P5_2|_RX|104  3.429952209
R_PTL_P5_2|_RX|B3 _PTL_P5_2|_RX|7 _PTL_P5_2|_RX|107  2.7439617672
L_PTL_P5_2|_RX|RB1 _PTL_P5_2|_RX|101 0  2.38752113364072e-12
L_PTL_P5_2|_RX|RB2 _PTL_P5_2|_RX|104 0  1.937922998085e-12
L_PTL_P5_2|_RX|RB3 _PTL_P5_2|_RX|107 0  1.550338398468e-12
B_PTL_G5_2|_TX|1 _PTL_G5_2|_TX|1 _PTL_G5_2|_TX|2 JJMIT AREA=2.5
B_PTL_G5_2|_TX|2 _PTL_G5_2|_TX|4 _PTL_G5_2|_TX|5 JJMIT AREA=2.5
I_PTL_G5_2|_TX|B1 0 _PTL_G5_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G5_2|_TX|B2 0 _PTL_G5_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G5_2|_TX|B1 _PTL_G5_2|_TX|1 _PTL_G5_2|_TX|3  1.684e-12
L_PTL_G5_2|_TX|B2 _PTL_G5_2|_TX|4 _PTL_G5_2|_TX|6  3.596e-12
L_PTL_G5_2|_TX|1 G5_2_TX _PTL_G5_2|_TX|1  2.063e-12
L_PTL_G5_2|_TX|2 _PTL_G5_2|_TX|1 _PTL_G5_2|_TX|4  4.123e-12
L_PTL_G5_2|_TX|3 _PTL_G5_2|_TX|4 _PTL_G5_2|_TX|7  2.193e-12
R_PTL_G5_2|_TX|D _PTL_G5_2|_TX|7 _PTL_G5_2|A_PTL  1.36
L_PTL_G5_2|_TX|P1 _PTL_G5_2|_TX|2 0  5.254e-13
L_PTL_G5_2|_TX|P2 _PTL_G5_2|_TX|5 0  5.141e-13
R_PTL_G5_2|_TX|B1 _PTL_G5_2|_TX|1 _PTL_G5_2|_TX|101  2.7439617672
R_PTL_G5_2|_TX|B2 _PTL_G5_2|_TX|4 _PTL_G5_2|_TX|104  2.7439617672
L_PTL_G5_2|_TX|RB1 _PTL_G5_2|_TX|101 0  1.550338398468e-12
L_PTL_G5_2|_TX|RB2 _PTL_G5_2|_TX|104 0  1.550338398468e-12
B_PTL_G5_2|_RX|1 _PTL_G5_2|_RX|1 _PTL_G5_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G5_2|_RX|2 _PTL_G5_2|_RX|4 _PTL_G5_2|_RX|5 JJMIT AREA=2.0
B_PTL_G5_2|_RX|3 _PTL_G5_2|_RX|7 _PTL_G5_2|_RX|8 JJMIT AREA=2.5
I_PTL_G5_2|_RX|B1 0 _PTL_G5_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G5_2|_RX|B1 _PTL_G5_2|_RX|1 _PTL_G5_2|_RX|3  2.777e-12
I_PTL_G5_2|_RX|B2 0 _PTL_G5_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G5_2|_RX|B2 _PTL_G5_2|_RX|4 _PTL_G5_2|_RX|6  2.685e-12
I_PTL_G5_2|_RX|B3 0 _PTL_G5_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G5_2|_RX|B3 _PTL_G5_2|_RX|7 _PTL_G5_2|_RX|9  2.764e-12
L_PTL_G5_2|_RX|1 _PTL_G5_2|A_PTL _PTL_G5_2|_RX|1  1.346e-12
L_PTL_G5_2|_RX|2 _PTL_G5_2|_RX|1 _PTL_G5_2|_RX|4  6.348e-12
L_PTL_G5_2|_RX|3 _PTL_G5_2|_RX|4 _PTL_G5_2|_RX|7  5.197e-12
L_PTL_G5_2|_RX|4 _PTL_G5_2|_RX|7 G5_2_TO5  2.058e-12
L_PTL_G5_2|_RX|P1 _PTL_G5_2|_RX|2 0  4.795e-13
L_PTL_G5_2|_RX|P2 _PTL_G5_2|_RX|5 0  5.431e-13
L_PTL_G5_2|_RX|P3 _PTL_G5_2|_RX|8 0  5.339e-13
R_PTL_G5_2|_RX|B1 _PTL_G5_2|_RX|1 _PTL_G5_2|_RX|101  4.225701121488
R_PTL_G5_2|_RX|B2 _PTL_G5_2|_RX|4 _PTL_G5_2|_RX|104  3.429952209
R_PTL_G5_2|_RX|B3 _PTL_G5_2|_RX|7 _PTL_G5_2|_RX|107  2.7439617672
L_PTL_G5_2|_RX|RB1 _PTL_G5_2|_RX|101 0  2.38752113364072e-12
L_PTL_G5_2|_RX|RB2 _PTL_G5_2|_RX|104 0  1.937922998085e-12
L_PTL_G5_2|_RX|RB3 _PTL_G5_2|_RX|107 0  1.550338398468e-12
B_PTL_P6_2|_TX|1 _PTL_P6_2|_TX|1 _PTL_P6_2|_TX|2 JJMIT AREA=2.5
B_PTL_P6_2|_TX|2 _PTL_P6_2|_TX|4 _PTL_P6_2|_TX|5 JJMIT AREA=2.5
I_PTL_P6_2|_TX|B1 0 _PTL_P6_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P6_2|_TX|B2 0 _PTL_P6_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P6_2|_TX|B1 _PTL_P6_2|_TX|1 _PTL_P6_2|_TX|3  1.684e-12
L_PTL_P6_2|_TX|B2 _PTL_P6_2|_TX|4 _PTL_P6_2|_TX|6  3.596e-12
L_PTL_P6_2|_TX|1 P6_2_TX _PTL_P6_2|_TX|1  2.063e-12
L_PTL_P6_2|_TX|2 _PTL_P6_2|_TX|1 _PTL_P6_2|_TX|4  4.123e-12
L_PTL_P6_2|_TX|3 _PTL_P6_2|_TX|4 _PTL_P6_2|_TX|7  2.193e-12
R_PTL_P6_2|_TX|D _PTL_P6_2|_TX|7 _PTL_P6_2|A_PTL  1.36
L_PTL_P6_2|_TX|P1 _PTL_P6_2|_TX|2 0  5.254e-13
L_PTL_P6_2|_TX|P2 _PTL_P6_2|_TX|5 0  5.141e-13
R_PTL_P6_2|_TX|B1 _PTL_P6_2|_TX|1 _PTL_P6_2|_TX|101  2.7439617672
R_PTL_P6_2|_TX|B2 _PTL_P6_2|_TX|4 _PTL_P6_2|_TX|104  2.7439617672
L_PTL_P6_2|_TX|RB1 _PTL_P6_2|_TX|101 0  1.550338398468e-12
L_PTL_P6_2|_TX|RB2 _PTL_P6_2|_TX|104 0  1.550338398468e-12
B_PTL_P6_2|_RX|1 _PTL_P6_2|_RX|1 _PTL_P6_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P6_2|_RX|2 _PTL_P6_2|_RX|4 _PTL_P6_2|_RX|5 JJMIT AREA=2.0
B_PTL_P6_2|_RX|3 _PTL_P6_2|_RX|7 _PTL_P6_2|_RX|8 JJMIT AREA=2.5
I_PTL_P6_2|_RX|B1 0 _PTL_P6_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P6_2|_RX|B1 _PTL_P6_2|_RX|1 _PTL_P6_2|_RX|3  2.777e-12
I_PTL_P6_2|_RX|B2 0 _PTL_P6_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P6_2|_RX|B2 _PTL_P6_2|_RX|4 _PTL_P6_2|_RX|6  2.685e-12
I_PTL_P6_2|_RX|B3 0 _PTL_P6_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P6_2|_RX|B3 _PTL_P6_2|_RX|7 _PTL_P6_2|_RX|9  2.764e-12
L_PTL_P6_2|_RX|1 _PTL_P6_2|A_PTL _PTL_P6_2|_RX|1  1.346e-12
L_PTL_P6_2|_RX|2 _PTL_P6_2|_RX|1 _PTL_P6_2|_RX|4  6.348e-12
L_PTL_P6_2|_RX|3 _PTL_P6_2|_RX|4 _PTL_P6_2|_RX|7  5.197e-12
L_PTL_P6_2|_RX|4 _PTL_P6_2|_RX|7 P6_2_TO6  2.058e-12
L_PTL_P6_2|_RX|P1 _PTL_P6_2|_RX|2 0  4.795e-13
L_PTL_P6_2|_RX|P2 _PTL_P6_2|_RX|5 0  5.431e-13
L_PTL_P6_2|_RX|P3 _PTL_P6_2|_RX|8 0  5.339e-13
R_PTL_P6_2|_RX|B1 _PTL_P6_2|_RX|1 _PTL_P6_2|_RX|101  4.225701121488
R_PTL_P6_2|_RX|B2 _PTL_P6_2|_RX|4 _PTL_P6_2|_RX|104  3.429952209
R_PTL_P6_2|_RX|B3 _PTL_P6_2|_RX|7 _PTL_P6_2|_RX|107  2.7439617672
L_PTL_P6_2|_RX|RB1 _PTL_P6_2|_RX|101 0  2.38752113364072e-12
L_PTL_P6_2|_RX|RB2 _PTL_P6_2|_RX|104 0  1.937922998085e-12
L_PTL_P6_2|_RX|RB3 _PTL_P6_2|_RX|107 0  1.550338398468e-12
B_PTL_G6_2|_TX|1 _PTL_G6_2|_TX|1 _PTL_G6_2|_TX|2 JJMIT AREA=2.5
B_PTL_G6_2|_TX|2 _PTL_G6_2|_TX|4 _PTL_G6_2|_TX|5 JJMIT AREA=2.5
I_PTL_G6_2|_TX|B1 0 _PTL_G6_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G6_2|_TX|B2 0 _PTL_G6_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G6_2|_TX|B1 _PTL_G6_2|_TX|1 _PTL_G6_2|_TX|3  1.684e-12
L_PTL_G6_2|_TX|B2 _PTL_G6_2|_TX|4 _PTL_G6_2|_TX|6  3.596e-12
L_PTL_G6_2|_TX|1 G6_2_TX _PTL_G6_2|_TX|1  2.063e-12
L_PTL_G6_2|_TX|2 _PTL_G6_2|_TX|1 _PTL_G6_2|_TX|4  4.123e-12
L_PTL_G6_2|_TX|3 _PTL_G6_2|_TX|4 _PTL_G6_2|_TX|7  2.193e-12
R_PTL_G6_2|_TX|D _PTL_G6_2|_TX|7 _PTL_G6_2|A_PTL  1.36
L_PTL_G6_2|_TX|P1 _PTL_G6_2|_TX|2 0  5.254e-13
L_PTL_G6_2|_TX|P2 _PTL_G6_2|_TX|5 0  5.141e-13
R_PTL_G6_2|_TX|B1 _PTL_G6_2|_TX|1 _PTL_G6_2|_TX|101  2.7439617672
R_PTL_G6_2|_TX|B2 _PTL_G6_2|_TX|4 _PTL_G6_2|_TX|104  2.7439617672
L_PTL_G6_2|_TX|RB1 _PTL_G6_2|_TX|101 0  1.550338398468e-12
L_PTL_G6_2|_TX|RB2 _PTL_G6_2|_TX|104 0  1.550338398468e-12
B_PTL_G6_2|_RX|1 _PTL_G6_2|_RX|1 _PTL_G6_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G6_2|_RX|2 _PTL_G6_2|_RX|4 _PTL_G6_2|_RX|5 JJMIT AREA=2.0
B_PTL_G6_2|_RX|3 _PTL_G6_2|_RX|7 _PTL_G6_2|_RX|8 JJMIT AREA=2.5
I_PTL_G6_2|_RX|B1 0 _PTL_G6_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G6_2|_RX|B1 _PTL_G6_2|_RX|1 _PTL_G6_2|_RX|3  2.777e-12
I_PTL_G6_2|_RX|B2 0 _PTL_G6_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G6_2|_RX|B2 _PTL_G6_2|_RX|4 _PTL_G6_2|_RX|6  2.685e-12
I_PTL_G6_2|_RX|B3 0 _PTL_G6_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G6_2|_RX|B3 _PTL_G6_2|_RX|7 _PTL_G6_2|_RX|9  2.764e-12
L_PTL_G6_2|_RX|1 _PTL_G6_2|A_PTL _PTL_G6_2|_RX|1  1.346e-12
L_PTL_G6_2|_RX|2 _PTL_G6_2|_RX|1 _PTL_G6_2|_RX|4  6.348e-12
L_PTL_G6_2|_RX|3 _PTL_G6_2|_RX|4 _PTL_G6_2|_RX|7  5.197e-12
L_PTL_G6_2|_RX|4 _PTL_G6_2|_RX|7 G6_2_TO6  2.058e-12
L_PTL_G6_2|_RX|P1 _PTL_G6_2|_RX|2 0  4.795e-13
L_PTL_G6_2|_RX|P2 _PTL_G6_2|_RX|5 0  5.431e-13
L_PTL_G6_2|_RX|P3 _PTL_G6_2|_RX|8 0  5.339e-13
R_PTL_G6_2|_RX|B1 _PTL_G6_2|_RX|1 _PTL_G6_2|_RX|101  4.225701121488
R_PTL_G6_2|_RX|B2 _PTL_G6_2|_RX|4 _PTL_G6_2|_RX|104  3.429952209
R_PTL_G6_2|_RX|B3 _PTL_G6_2|_RX|7 _PTL_G6_2|_RX|107  2.7439617672
L_PTL_G6_2|_RX|RB1 _PTL_G6_2|_RX|101 0  2.38752113364072e-12
L_PTL_G6_2|_RX|RB2 _PTL_G6_2|_RX|104 0  1.937922998085e-12
L_PTL_G6_2|_RX|RB3 _PTL_G6_2|_RX|107 0  1.550338398468e-12
B_PTL_IP7_2|_TX|1 _PTL_IP7_2|_TX|1 _PTL_IP7_2|_TX|2 JJMIT AREA=2.5
B_PTL_IP7_2|_TX|2 _PTL_IP7_2|_TX|4 _PTL_IP7_2|_TX|5 JJMIT AREA=2.5
I_PTL_IP7_2|_TX|B1 0 _PTL_IP7_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP7_2|_TX|B2 0 _PTL_IP7_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_2|_TX|B1 _PTL_IP7_2|_TX|1 _PTL_IP7_2|_TX|3  1.684e-12
L_PTL_IP7_2|_TX|B2 _PTL_IP7_2|_TX|4 _PTL_IP7_2|_TX|6  3.596e-12
L_PTL_IP7_2|_TX|1 IP7_2_OUT_TX _PTL_IP7_2|_TX|1  2.063e-12
L_PTL_IP7_2|_TX|2 _PTL_IP7_2|_TX|1 _PTL_IP7_2|_TX|4  4.123e-12
L_PTL_IP7_2|_TX|3 _PTL_IP7_2|_TX|4 _PTL_IP7_2|_TX|7  2.193e-12
R_PTL_IP7_2|_TX|D _PTL_IP7_2|_TX|7 _PTL_IP7_2|A_PTL  1.36
L_PTL_IP7_2|_TX|P1 _PTL_IP7_2|_TX|2 0  5.254e-13
L_PTL_IP7_2|_TX|P2 _PTL_IP7_2|_TX|5 0  5.141e-13
R_PTL_IP7_2|_TX|B1 _PTL_IP7_2|_TX|1 _PTL_IP7_2|_TX|101  2.7439617672
R_PTL_IP7_2|_TX|B2 _PTL_IP7_2|_TX|4 _PTL_IP7_2|_TX|104  2.7439617672
L_PTL_IP7_2|_TX|RB1 _PTL_IP7_2|_TX|101 0  1.550338398468e-12
L_PTL_IP7_2|_TX|RB2 _PTL_IP7_2|_TX|104 0  1.550338398468e-12
B_PTL_IP7_2|_RX|1 _PTL_IP7_2|_RX|1 _PTL_IP7_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP7_2|_RX|2 _PTL_IP7_2|_RX|4 _PTL_IP7_2|_RX|5 JJMIT AREA=2.0
B_PTL_IP7_2|_RX|3 _PTL_IP7_2|_RX|7 _PTL_IP7_2|_RX|8 JJMIT AREA=2.5
I_PTL_IP7_2|_RX|B1 0 _PTL_IP7_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP7_2|_RX|B1 _PTL_IP7_2|_RX|1 _PTL_IP7_2|_RX|3  2.777e-12
I_PTL_IP7_2|_RX|B2 0 _PTL_IP7_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP7_2|_RX|B2 _PTL_IP7_2|_RX|4 _PTL_IP7_2|_RX|6  2.685e-12
I_PTL_IP7_2|_RX|B3 0 _PTL_IP7_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_2|_RX|B3 _PTL_IP7_2|_RX|7 _PTL_IP7_2|_RX|9  2.764e-12
L_PTL_IP7_2|_RX|1 _PTL_IP7_2|A_PTL _PTL_IP7_2|_RX|1  1.346e-12
L_PTL_IP7_2|_RX|2 _PTL_IP7_2|_RX|1 _PTL_IP7_2|_RX|4  6.348e-12
L_PTL_IP7_2|_RX|3 _PTL_IP7_2|_RX|4 _PTL_IP7_2|_RX|7  5.197e-12
L_PTL_IP7_2|_RX|4 _PTL_IP7_2|_RX|7 IP7_2_OUT  2.058e-12
L_PTL_IP7_2|_RX|P1 _PTL_IP7_2|_RX|2 0  4.795e-13
L_PTL_IP7_2|_RX|P2 _PTL_IP7_2|_RX|5 0  5.431e-13
L_PTL_IP7_2|_RX|P3 _PTL_IP7_2|_RX|8 0  5.339e-13
R_PTL_IP7_2|_RX|B1 _PTL_IP7_2|_RX|1 _PTL_IP7_2|_RX|101  4.225701121488
R_PTL_IP7_2|_RX|B2 _PTL_IP7_2|_RX|4 _PTL_IP7_2|_RX|104  3.429952209
R_PTL_IP7_2|_RX|B3 _PTL_IP7_2|_RX|7 _PTL_IP7_2|_RX|107  2.7439617672
L_PTL_IP7_2|_RX|RB1 _PTL_IP7_2|_RX|101 0  2.38752113364072e-12
L_PTL_IP7_2|_RX|RB2 _PTL_IP7_2|_RX|104 0  1.937922998085e-12
L_PTL_IP7_2|_RX|RB3 _PTL_IP7_2|_RX|107 0  1.550338398468e-12
B_PTL_P7_2|_TX|1 _PTL_P7_2|_TX|1 _PTL_P7_2|_TX|2 JJMIT AREA=2.5
B_PTL_P7_2|_TX|2 _PTL_P7_2|_TX|4 _PTL_P7_2|_TX|5 JJMIT AREA=2.5
I_PTL_P7_2|_TX|B1 0 _PTL_P7_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P7_2|_TX|B2 0 _PTL_P7_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P7_2|_TX|B1 _PTL_P7_2|_TX|1 _PTL_P7_2|_TX|3  1.684e-12
L_PTL_P7_2|_TX|B2 _PTL_P7_2|_TX|4 _PTL_P7_2|_TX|6  3.596e-12
L_PTL_P7_2|_TX|1 P7_2_TX _PTL_P7_2|_TX|1  2.063e-12
L_PTL_P7_2|_TX|2 _PTL_P7_2|_TX|1 _PTL_P7_2|_TX|4  4.123e-12
L_PTL_P7_2|_TX|3 _PTL_P7_2|_TX|4 _PTL_P7_2|_TX|7  2.193e-12
R_PTL_P7_2|_TX|D _PTL_P7_2|_TX|7 _PTL_P7_2|A_PTL  1.36
L_PTL_P7_2|_TX|P1 _PTL_P7_2|_TX|2 0  5.254e-13
L_PTL_P7_2|_TX|P2 _PTL_P7_2|_TX|5 0  5.141e-13
R_PTL_P7_2|_TX|B1 _PTL_P7_2|_TX|1 _PTL_P7_2|_TX|101  2.7439617672
R_PTL_P7_2|_TX|B2 _PTL_P7_2|_TX|4 _PTL_P7_2|_TX|104  2.7439617672
L_PTL_P7_2|_TX|RB1 _PTL_P7_2|_TX|101 0  1.550338398468e-12
L_PTL_P7_2|_TX|RB2 _PTL_P7_2|_TX|104 0  1.550338398468e-12
B_PTL_P7_2|_RX|1 _PTL_P7_2|_RX|1 _PTL_P7_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P7_2|_RX|2 _PTL_P7_2|_RX|4 _PTL_P7_2|_RX|5 JJMIT AREA=2.0
B_PTL_P7_2|_RX|3 _PTL_P7_2|_RX|7 _PTL_P7_2|_RX|8 JJMIT AREA=2.5
I_PTL_P7_2|_RX|B1 0 _PTL_P7_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P7_2|_RX|B1 _PTL_P7_2|_RX|1 _PTL_P7_2|_RX|3  2.777e-12
I_PTL_P7_2|_RX|B2 0 _PTL_P7_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P7_2|_RX|B2 _PTL_P7_2|_RX|4 _PTL_P7_2|_RX|6  2.685e-12
I_PTL_P7_2|_RX|B3 0 _PTL_P7_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P7_2|_RX|B3 _PTL_P7_2|_RX|7 _PTL_P7_2|_RX|9  2.764e-12
L_PTL_P7_2|_RX|1 _PTL_P7_2|A_PTL _PTL_P7_2|_RX|1  1.346e-12
L_PTL_P7_2|_RX|2 _PTL_P7_2|_RX|1 _PTL_P7_2|_RX|4  6.348e-12
L_PTL_P7_2|_RX|3 _PTL_P7_2|_RX|4 _PTL_P7_2|_RX|7  5.197e-12
L_PTL_P7_2|_RX|4 _PTL_P7_2|_RX|7 P7_2_TO7  2.058e-12
L_PTL_P7_2|_RX|P1 _PTL_P7_2|_RX|2 0  4.795e-13
L_PTL_P7_2|_RX|P2 _PTL_P7_2|_RX|5 0  5.431e-13
L_PTL_P7_2|_RX|P3 _PTL_P7_2|_RX|8 0  5.339e-13
R_PTL_P7_2|_RX|B1 _PTL_P7_2|_RX|1 _PTL_P7_2|_RX|101  4.225701121488
R_PTL_P7_2|_RX|B2 _PTL_P7_2|_RX|4 _PTL_P7_2|_RX|104  3.429952209
R_PTL_P7_2|_RX|B3 _PTL_P7_2|_RX|7 _PTL_P7_2|_RX|107  2.7439617672
L_PTL_P7_2|_RX|RB1 _PTL_P7_2|_RX|101 0  2.38752113364072e-12
L_PTL_P7_2|_RX|RB2 _PTL_P7_2|_RX|104 0  1.937922998085e-12
L_PTL_P7_2|_RX|RB3 _PTL_P7_2|_RX|107 0  1.550338398468e-12
B_PTL_G7_2|_TX|1 _PTL_G7_2|_TX|1 _PTL_G7_2|_TX|2 JJMIT AREA=2.5
B_PTL_G7_2|_TX|2 _PTL_G7_2|_TX|4 _PTL_G7_2|_TX|5 JJMIT AREA=2.5
I_PTL_G7_2|_TX|B1 0 _PTL_G7_2|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G7_2|_TX|B2 0 _PTL_G7_2|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G7_2|_TX|B1 _PTL_G7_2|_TX|1 _PTL_G7_2|_TX|3  1.684e-12
L_PTL_G7_2|_TX|B2 _PTL_G7_2|_TX|4 _PTL_G7_2|_TX|6  3.596e-12
L_PTL_G7_2|_TX|1 G7_2_TX _PTL_G7_2|_TX|1  2.063e-12
L_PTL_G7_2|_TX|2 _PTL_G7_2|_TX|1 _PTL_G7_2|_TX|4  4.123e-12
L_PTL_G7_2|_TX|3 _PTL_G7_2|_TX|4 _PTL_G7_2|_TX|7  2.193e-12
R_PTL_G7_2|_TX|D _PTL_G7_2|_TX|7 _PTL_G7_2|A_PTL  1.36
L_PTL_G7_2|_TX|P1 _PTL_G7_2|_TX|2 0  5.254e-13
L_PTL_G7_2|_TX|P2 _PTL_G7_2|_TX|5 0  5.141e-13
R_PTL_G7_2|_TX|B1 _PTL_G7_2|_TX|1 _PTL_G7_2|_TX|101  2.7439617672
R_PTL_G7_2|_TX|B2 _PTL_G7_2|_TX|4 _PTL_G7_2|_TX|104  2.7439617672
L_PTL_G7_2|_TX|RB1 _PTL_G7_2|_TX|101 0  1.550338398468e-12
L_PTL_G7_2|_TX|RB2 _PTL_G7_2|_TX|104 0  1.550338398468e-12
B_PTL_G7_2|_RX|1 _PTL_G7_2|_RX|1 _PTL_G7_2|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G7_2|_RX|2 _PTL_G7_2|_RX|4 _PTL_G7_2|_RX|5 JJMIT AREA=2.0
B_PTL_G7_2|_RX|3 _PTL_G7_2|_RX|7 _PTL_G7_2|_RX|8 JJMIT AREA=2.5
I_PTL_G7_2|_RX|B1 0 _PTL_G7_2|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G7_2|_RX|B1 _PTL_G7_2|_RX|1 _PTL_G7_2|_RX|3  2.777e-12
I_PTL_G7_2|_RX|B2 0 _PTL_G7_2|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G7_2|_RX|B2 _PTL_G7_2|_RX|4 _PTL_G7_2|_RX|6  2.685e-12
I_PTL_G7_2|_RX|B3 0 _PTL_G7_2|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G7_2|_RX|B3 _PTL_G7_2|_RX|7 _PTL_G7_2|_RX|9  2.764e-12
L_PTL_G7_2|_RX|1 _PTL_G7_2|A_PTL _PTL_G7_2|_RX|1  1.346e-12
L_PTL_G7_2|_RX|2 _PTL_G7_2|_RX|1 _PTL_G7_2|_RX|4  6.348e-12
L_PTL_G7_2|_RX|3 _PTL_G7_2|_RX|4 _PTL_G7_2|_RX|7  5.197e-12
L_PTL_G7_2|_RX|4 _PTL_G7_2|_RX|7 G7_2_TO7  2.058e-12
L_PTL_G7_2|_RX|P1 _PTL_G7_2|_RX|2 0  4.795e-13
L_PTL_G7_2|_RX|P2 _PTL_G7_2|_RX|5 0  5.431e-13
L_PTL_G7_2|_RX|P3 _PTL_G7_2|_RX|8 0  5.339e-13
R_PTL_G7_2|_RX|B1 _PTL_G7_2|_RX|1 _PTL_G7_2|_RX|101  4.225701121488
R_PTL_G7_2|_RX|B2 _PTL_G7_2|_RX|4 _PTL_G7_2|_RX|104  3.429952209
R_PTL_G7_2|_RX|B3 _PTL_G7_2|_RX|7 _PTL_G7_2|_RX|107  2.7439617672
L_PTL_G7_2|_RX|RB1 _PTL_G7_2|_RX|101 0  2.38752113364072e-12
L_PTL_G7_2|_RX|RB2 _PTL_G7_2|_RX|104 0  1.937922998085e-12
L_PTL_G7_2|_RX|RB3 _PTL_G7_2|_RX|107 0  1.550338398468e-12
L_S0_23|I_1|B _S0_23|A1 _S0_23|I_1|MID  2e-12
I_S0_23|I_1|B 0 _S0_23|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0_23|I_3|B _S0_23|A3 _S0_23|I_3|MID  2e-12
I_S0_23|I_3|B 0 _S0_23|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0_23|I_T|B _S0_23|T1 _S0_23|I_T|MID  2e-12
I_S0_23|I_T|B 0 _S0_23|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0_23|I_6|B _S0_23|Q1 _S0_23|I_6|MID  2e-12
I_S0_23|I_6|B 0 _S0_23|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0_23|1|1 _S0_23|A1 _S0_23|1|MID_SERIES JJMIT AREA=2.5
L_S0_23|1|P _S0_23|1|MID_SERIES 0  2e-13
R_S0_23|1|B _S0_23|A1 _S0_23|1|MID_SHUNT  2.7439617672
L_S0_23|1|RB _S0_23|1|MID_SHUNT 0  1.550338398468e-12
B_S0_23|23|1 _S0_23|A2 _S0_23|A3 JJMIT AREA=1.7857142857142858
R_S0_23|23|B _S0_23|A2 _S0_23|23|MID_SHUNT  3.84154647408
L_S0_23|23|RB _S0_23|23|MID_SHUNT _S0_23|A3  2.1704737578552e-12
B_S0_23|3|1 _S0_23|A3 _S0_23|3|MID_SERIES JJMIT AREA=2.5
L_S0_23|3|P _S0_23|3|MID_SERIES 0  2e-13
R_S0_23|3|B _S0_23|A3 _S0_23|3|MID_SHUNT  2.7439617672
L_S0_23|3|RB _S0_23|3|MID_SHUNT 0  1.550338398468e-12
B_S0_23|4|1 _S0_23|A4 _S0_23|4|MID_SERIES JJMIT AREA=2.5
L_S0_23|4|P _S0_23|4|MID_SERIES 0  2e-13
R_S0_23|4|B _S0_23|A4 _S0_23|4|MID_SHUNT  2.7439617672
L_S0_23|4|RB _S0_23|4|MID_SHUNT 0  1.550338398468e-12
B_S0_23|T|1 _S0_23|T1 _S0_23|T|MID_SERIES JJMIT AREA=2.5
L_S0_23|T|P _S0_23|T|MID_SERIES 0  2e-13
R_S0_23|T|B _S0_23|T1 _S0_23|T|MID_SHUNT  2.7439617672
L_S0_23|T|RB _S0_23|T|MID_SHUNT 0  1.550338398468e-12
B_S0_23|45|1 _S0_23|T2 _S0_23|A4 JJMIT AREA=1.7857142857142858
R_S0_23|45|B _S0_23|T2 _S0_23|45|MID_SHUNT  3.84154647408
L_S0_23|45|RB _S0_23|45|MID_SHUNT _S0_23|A4  2.1704737578552e-12
B_S0_23|6|1 _S0_23|Q1 _S0_23|6|MID_SERIES JJMIT AREA=2.5
L_S0_23|6|P _S0_23|6|MID_SERIES 0  2e-13
R_S0_23|6|B _S0_23|Q1 _S0_23|6|MID_SHUNT  2.7439617672
L_S0_23|6|RB _S0_23|6|MID_SHUNT 0  1.550338398468e-12
L_S1_23|I_1|B _S1_23|A1 _S1_23|I_1|MID  2e-12
I_S1_23|I_1|B 0 _S1_23|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S1_23|I_3|B _S1_23|A3 _S1_23|I_3|MID  2e-12
I_S1_23|I_3|B 0 _S1_23|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S1_23|I_T|B _S1_23|T1 _S1_23|I_T|MID  2e-12
I_S1_23|I_T|B 0 _S1_23|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S1_23|I_6|B _S1_23|Q1 _S1_23|I_6|MID  2e-12
I_S1_23|I_6|B 0 _S1_23|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S1_23|1|1 _S1_23|A1 _S1_23|1|MID_SERIES JJMIT AREA=2.5
L_S1_23|1|P _S1_23|1|MID_SERIES 0  2e-13
R_S1_23|1|B _S1_23|A1 _S1_23|1|MID_SHUNT  2.7439617672
L_S1_23|1|RB _S1_23|1|MID_SHUNT 0  1.550338398468e-12
B_S1_23|23|1 _S1_23|A2 _S1_23|A3 JJMIT AREA=1.7857142857142858
R_S1_23|23|B _S1_23|A2 _S1_23|23|MID_SHUNT  3.84154647408
L_S1_23|23|RB _S1_23|23|MID_SHUNT _S1_23|A3  2.1704737578552e-12
B_S1_23|3|1 _S1_23|A3 _S1_23|3|MID_SERIES JJMIT AREA=2.5
L_S1_23|3|P _S1_23|3|MID_SERIES 0  2e-13
R_S1_23|3|B _S1_23|A3 _S1_23|3|MID_SHUNT  2.7439617672
L_S1_23|3|RB _S1_23|3|MID_SHUNT 0  1.550338398468e-12
B_S1_23|4|1 _S1_23|A4 _S1_23|4|MID_SERIES JJMIT AREA=2.5
L_S1_23|4|P _S1_23|4|MID_SERIES 0  2e-13
R_S1_23|4|B _S1_23|A4 _S1_23|4|MID_SHUNT  2.7439617672
L_S1_23|4|RB _S1_23|4|MID_SHUNT 0  1.550338398468e-12
B_S1_23|T|1 _S1_23|T1 _S1_23|T|MID_SERIES JJMIT AREA=2.5
L_S1_23|T|P _S1_23|T|MID_SERIES 0  2e-13
R_S1_23|T|B _S1_23|T1 _S1_23|T|MID_SHUNT  2.7439617672
L_S1_23|T|RB _S1_23|T|MID_SHUNT 0  1.550338398468e-12
B_S1_23|45|1 _S1_23|T2 _S1_23|A4 JJMIT AREA=1.7857142857142858
R_S1_23|45|B _S1_23|T2 _S1_23|45|MID_SHUNT  3.84154647408
L_S1_23|45|RB _S1_23|45|MID_SHUNT _S1_23|A4  2.1704737578552e-12
B_S1_23|6|1 _S1_23|Q1 _S1_23|6|MID_SERIES JJMIT AREA=2.5
L_S1_23|6|P _S1_23|6|MID_SERIES 0  2e-13
R_S1_23|6|B _S1_23|Q1 _S1_23|6|MID_SHUNT  2.7439617672
L_S1_23|6|RB _S1_23|6|MID_SHUNT 0  1.550338398468e-12
L_S2_23|I_1|B _S2_23|A1 _S2_23|I_1|MID  2e-12
I_S2_23|I_1|B 0 _S2_23|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S2_23|I_3|B _S2_23|A3 _S2_23|I_3|MID  2e-12
I_S2_23|I_3|B 0 _S2_23|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S2_23|I_T|B _S2_23|T1 _S2_23|I_T|MID  2e-12
I_S2_23|I_T|B 0 _S2_23|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S2_23|I_6|B _S2_23|Q1 _S2_23|I_6|MID  2e-12
I_S2_23|I_6|B 0 _S2_23|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S2_23|1|1 _S2_23|A1 _S2_23|1|MID_SERIES JJMIT AREA=2.5
L_S2_23|1|P _S2_23|1|MID_SERIES 0  2e-13
R_S2_23|1|B _S2_23|A1 _S2_23|1|MID_SHUNT  2.7439617672
L_S2_23|1|RB _S2_23|1|MID_SHUNT 0  1.550338398468e-12
B_S2_23|23|1 _S2_23|A2 _S2_23|A3 JJMIT AREA=1.7857142857142858
R_S2_23|23|B _S2_23|A2 _S2_23|23|MID_SHUNT  3.84154647408
L_S2_23|23|RB _S2_23|23|MID_SHUNT _S2_23|A3  2.1704737578552e-12
B_S2_23|3|1 _S2_23|A3 _S2_23|3|MID_SERIES JJMIT AREA=2.5
L_S2_23|3|P _S2_23|3|MID_SERIES 0  2e-13
R_S2_23|3|B _S2_23|A3 _S2_23|3|MID_SHUNT  2.7439617672
L_S2_23|3|RB _S2_23|3|MID_SHUNT 0  1.550338398468e-12
B_S2_23|4|1 _S2_23|A4 _S2_23|4|MID_SERIES JJMIT AREA=2.5
L_S2_23|4|P _S2_23|4|MID_SERIES 0  2e-13
R_S2_23|4|B _S2_23|A4 _S2_23|4|MID_SHUNT  2.7439617672
L_S2_23|4|RB _S2_23|4|MID_SHUNT 0  1.550338398468e-12
B_S2_23|T|1 _S2_23|T1 _S2_23|T|MID_SERIES JJMIT AREA=2.5
L_S2_23|T|P _S2_23|T|MID_SERIES 0  2e-13
R_S2_23|T|B _S2_23|T1 _S2_23|T|MID_SHUNT  2.7439617672
L_S2_23|T|RB _S2_23|T|MID_SHUNT 0  1.550338398468e-12
B_S2_23|45|1 _S2_23|T2 _S2_23|A4 JJMIT AREA=1.7857142857142858
R_S2_23|45|B _S2_23|T2 _S2_23|45|MID_SHUNT  3.84154647408
L_S2_23|45|RB _S2_23|45|MID_SHUNT _S2_23|A4  2.1704737578552e-12
B_S2_23|6|1 _S2_23|Q1 _S2_23|6|MID_SERIES JJMIT AREA=2.5
L_S2_23|6|P _S2_23|6|MID_SERIES 0  2e-13
R_S2_23|6|B _S2_23|Q1 _S2_23|6|MID_SHUNT  2.7439617672
L_S2_23|6|RB _S2_23|6|MID_SHUNT 0  1.550338398468e-12
L_S3_23|I_A1|B _S3_23|A1 _S3_23|I_A1|MID  2e-12
I_S3_23|I_A1|B 0 _S3_23|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S3_23|I_A3|B _S3_23|A3 _S3_23|I_A3|MID  2e-12
I_S3_23|I_A3|B 0 _S3_23|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S3_23|I_B1|B _S3_23|B1 _S3_23|I_B1|MID  2e-12
I_S3_23|I_B1|B 0 _S3_23|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S3_23|I_B3|B _S3_23|B3 _S3_23|I_B3|MID  2e-12
I_S3_23|I_B3|B 0 _S3_23|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S3_23|I_Q1|B _S3_23|Q1 _S3_23|I_Q1|MID  2e-12
I_S3_23|I_Q1|B 0 _S3_23|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S3_23|A1|1 _S3_23|A1 _S3_23|A1|MID_SERIES JJMIT AREA=2.5
L_S3_23|A1|P _S3_23|A1|MID_SERIES 0  5e-13
R_S3_23|A1|B _S3_23|A1 _S3_23|A1|MID_SHUNT  2.7439617672
L_S3_23|A1|RB _S3_23|A1|MID_SHUNT 0  2.050338398468e-12
B_S3_23|A2|1 _S3_23|A2 _S3_23|A2|MID_SERIES JJMIT AREA=2.5
L_S3_23|A2|P _S3_23|A2|MID_SERIES 0  5e-13
R_S3_23|A2|B _S3_23|A2 _S3_23|A2|MID_SHUNT  2.7439617672
L_S3_23|A2|RB _S3_23|A2|MID_SHUNT 0  2.050338398468e-12
B_S3_23|A3|1 _S3_23|A2 _S3_23|A3|MID_SERIES JJMIT AREA=2.5
L_S3_23|A3|P _S3_23|A3|MID_SERIES _S3_23|A3  1.2e-12
R_S3_23|A3|B _S3_23|A2 _S3_23|A3|MID_SHUNT  2.7439617672
L_S3_23|A3|RB _S3_23|A3|MID_SHUNT _S3_23|A3  2.050338398468e-12
B_S3_23|B1|1 _S3_23|B1 _S3_23|B1|MID_SERIES JJMIT AREA=2.5
L_S3_23|B1|P _S3_23|B1|MID_SERIES 0  5e-13
R_S3_23|B1|B _S3_23|B1 _S3_23|B1|MID_SHUNT  2.7439617672
L_S3_23|B1|RB _S3_23|B1|MID_SHUNT 0  2.050338398468e-12
B_S3_23|B2|1 _S3_23|B2 _S3_23|B2|MID_SERIES JJMIT AREA=2.5
L_S3_23|B2|P _S3_23|B2|MID_SERIES 0  5e-13
R_S3_23|B2|B _S3_23|B2 _S3_23|B2|MID_SHUNT  2.7439617672
L_S3_23|B2|RB _S3_23|B2|MID_SHUNT 0  2.050338398468e-12
B_S3_23|B3|1 _S3_23|B2 _S3_23|B3|MID_SERIES JJMIT AREA=2.5
L_S3_23|B3|P _S3_23|B3|MID_SERIES _S3_23|B3  1.2e-12
R_S3_23|B3|B _S3_23|B2 _S3_23|B3|MID_SHUNT  2.7439617672
L_S3_23|B3|RB _S3_23|B3|MID_SHUNT _S3_23|B3  2.050338398468e-12
B_S3_23|T1|1 _S3_23|T1 _S3_23|T1|MID_SERIES JJMIT AREA=2.5
L_S3_23|T1|P _S3_23|T1|MID_SERIES 0  5e-13
R_S3_23|T1|B _S3_23|T1 _S3_23|T1|MID_SHUNT  2.7439617672
L_S3_23|T1|RB _S3_23|T1|MID_SHUNT 0  2.050338398468e-12
B_S3_23|T2|1 _S3_23|T2 _S3_23|ABTQ JJMIT AREA=2.0
R_S3_23|T2|B _S3_23|T2 _S3_23|T2|MID_SHUNT  3.429952209
L_S3_23|T2|RB _S3_23|T2|MID_SHUNT _S3_23|ABTQ  2.437922998085e-12
B_S3_23|AB|1 _S3_23|AB _S3_23|AB|MID_SERIES JJMIT AREA=1.5
L_S3_23|AB|P _S3_23|AB|MID_SERIES _S3_23|ABTQ  1.2e-12
R_S3_23|AB|B _S3_23|AB _S3_23|AB|MID_SHUNT  4.573269612
L_S3_23|AB|RB _S3_23|AB|MID_SHUNT _S3_23|ABTQ  3.08389733078e-12
B_S3_23|ABTQ|1 _S3_23|ABTQ _S3_23|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S3_23|ABTQ|P _S3_23|ABTQ|MID_SERIES 0  5e-13
R_S3_23|ABTQ|B _S3_23|ABTQ _S3_23|ABTQ|MID_SHUNT  3.6586156896
L_S3_23|ABTQ|RB _S3_23|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S3_23|Q1|1 _S3_23|Q1 _S3_23|Q1|MID_SERIES JJMIT AREA=2.5
L_S3_23|Q1|P _S3_23|Q1|MID_SERIES 0  5e-13
R_S3_23|Q1|B _S3_23|Q1 _S3_23|Q1|MID_SHUNT  2.7439617672
L_S3_23|Q1|RB _S3_23|Q1|MID_SHUNT 0  2.050338398468e-12
L_S4_23|I_A1|B _S4_23|A1 _S4_23|I_A1|MID  2e-12
I_S4_23|I_A1|B 0 _S4_23|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S4_23|I_A3|B _S4_23|A3 _S4_23|I_A3|MID  2e-12
I_S4_23|I_A3|B 0 _S4_23|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S4_23|I_B1|B _S4_23|B1 _S4_23|I_B1|MID  2e-12
I_S4_23|I_B1|B 0 _S4_23|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S4_23|I_B3|B _S4_23|B3 _S4_23|I_B3|MID  2e-12
I_S4_23|I_B3|B 0 _S4_23|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S4_23|I_Q1|B _S4_23|Q1 _S4_23|I_Q1|MID  2e-12
I_S4_23|I_Q1|B 0 _S4_23|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S4_23|A1|1 _S4_23|A1 _S4_23|A1|MID_SERIES JJMIT AREA=2.5
L_S4_23|A1|P _S4_23|A1|MID_SERIES 0  5e-13
R_S4_23|A1|B _S4_23|A1 _S4_23|A1|MID_SHUNT  2.7439617672
L_S4_23|A1|RB _S4_23|A1|MID_SHUNT 0  2.050338398468e-12
B_S4_23|A2|1 _S4_23|A2 _S4_23|A2|MID_SERIES JJMIT AREA=2.5
L_S4_23|A2|P _S4_23|A2|MID_SERIES 0  5e-13
R_S4_23|A2|B _S4_23|A2 _S4_23|A2|MID_SHUNT  2.7439617672
L_S4_23|A2|RB _S4_23|A2|MID_SHUNT 0  2.050338398468e-12
B_S4_23|A3|1 _S4_23|A2 _S4_23|A3|MID_SERIES JJMIT AREA=2.5
L_S4_23|A3|P _S4_23|A3|MID_SERIES _S4_23|A3  1.2e-12
R_S4_23|A3|B _S4_23|A2 _S4_23|A3|MID_SHUNT  2.7439617672
L_S4_23|A3|RB _S4_23|A3|MID_SHUNT _S4_23|A3  2.050338398468e-12
B_S4_23|B1|1 _S4_23|B1 _S4_23|B1|MID_SERIES JJMIT AREA=2.5
L_S4_23|B1|P _S4_23|B1|MID_SERIES 0  5e-13
R_S4_23|B1|B _S4_23|B1 _S4_23|B1|MID_SHUNT  2.7439617672
L_S4_23|B1|RB _S4_23|B1|MID_SHUNT 0  2.050338398468e-12
B_S4_23|B2|1 _S4_23|B2 _S4_23|B2|MID_SERIES JJMIT AREA=2.5
L_S4_23|B2|P _S4_23|B2|MID_SERIES 0  5e-13
R_S4_23|B2|B _S4_23|B2 _S4_23|B2|MID_SHUNT  2.7439617672
L_S4_23|B2|RB _S4_23|B2|MID_SHUNT 0  2.050338398468e-12
B_S4_23|B3|1 _S4_23|B2 _S4_23|B3|MID_SERIES JJMIT AREA=2.5
L_S4_23|B3|P _S4_23|B3|MID_SERIES _S4_23|B3  1.2e-12
R_S4_23|B3|B _S4_23|B2 _S4_23|B3|MID_SHUNT  2.7439617672
L_S4_23|B3|RB _S4_23|B3|MID_SHUNT _S4_23|B3  2.050338398468e-12
B_S4_23|T1|1 _S4_23|T1 _S4_23|T1|MID_SERIES JJMIT AREA=2.5
L_S4_23|T1|P _S4_23|T1|MID_SERIES 0  5e-13
R_S4_23|T1|B _S4_23|T1 _S4_23|T1|MID_SHUNT  2.7439617672
L_S4_23|T1|RB _S4_23|T1|MID_SHUNT 0  2.050338398468e-12
B_S4_23|T2|1 _S4_23|T2 _S4_23|ABTQ JJMIT AREA=2.0
R_S4_23|T2|B _S4_23|T2 _S4_23|T2|MID_SHUNT  3.429952209
L_S4_23|T2|RB _S4_23|T2|MID_SHUNT _S4_23|ABTQ  2.437922998085e-12
B_S4_23|AB|1 _S4_23|AB _S4_23|AB|MID_SERIES JJMIT AREA=1.5
L_S4_23|AB|P _S4_23|AB|MID_SERIES _S4_23|ABTQ  1.2e-12
R_S4_23|AB|B _S4_23|AB _S4_23|AB|MID_SHUNT  4.573269612
L_S4_23|AB|RB _S4_23|AB|MID_SHUNT _S4_23|ABTQ  3.08389733078e-12
B_S4_23|ABTQ|1 _S4_23|ABTQ _S4_23|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S4_23|ABTQ|P _S4_23|ABTQ|MID_SERIES 0  5e-13
R_S4_23|ABTQ|B _S4_23|ABTQ _S4_23|ABTQ|MID_SHUNT  3.6586156896
L_S4_23|ABTQ|RB _S4_23|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S4_23|Q1|1 _S4_23|Q1 _S4_23|Q1|MID_SERIES JJMIT AREA=2.5
L_S4_23|Q1|P _S4_23|Q1|MID_SERIES 0  5e-13
R_S4_23|Q1|B _S4_23|Q1 _S4_23|Q1|MID_SHUNT  2.7439617672
L_S4_23|Q1|RB _S4_23|Q1|MID_SHUNT 0  2.050338398468e-12
L_PG4_23|_SPL_G1|1 G4_2_TO4 _PG4_23|_SPL_G1|D1  2e-12
L_PG4_23|_SPL_G1|2 _PG4_23|_SPL_G1|D1 _PG4_23|_SPL_G1|D2  4.135667696e-12
L_PG4_23|_SPL_G1|3 _PG4_23|_SPL_G1|D2 _PG4_23|_SPL_G1|JCT  9.84682784761905e-13
L_PG4_23|_SPL_G1|4 _PG4_23|_SPL_G1|JCT _PG4_23|_SPL_G1|QA1  9.84682784761905e-13
L_PG4_23|_SPL_G1|5 _PG4_23|_SPL_G1|QA1 _PG4_23|G1_COPY_1  2e-12
L_PG4_23|_SPL_G1|6 _PG4_23|_SPL_G1|JCT _PG4_23|_SPL_G1|QB1  9.84682784761905e-13
L_PG4_23|_SPL_G1|7 _PG4_23|_SPL_G1|QB1 _PG4_23|G1_COPY_2  2e-12
L_PG4_23|_SPL_P1|1 P4_2_TO4 _PG4_23|_SPL_P1|D1  2e-12
L_PG4_23|_SPL_P1|2 _PG4_23|_SPL_P1|D1 _PG4_23|_SPL_P1|D2  4.135667696e-12
L_PG4_23|_SPL_P1|3 _PG4_23|_SPL_P1|D2 _PG4_23|_SPL_P1|JCT  9.84682784761905e-13
L_PG4_23|_SPL_P1|4 _PG4_23|_SPL_P1|JCT _PG4_23|_SPL_P1|QA1  9.84682784761905e-13
L_PG4_23|_SPL_P1|5 _PG4_23|_SPL_P1|QA1 _PG4_23|P1_COPY_1  2e-12
L_PG4_23|_SPL_P1|6 _PG4_23|_SPL_P1|JCT _PG4_23|_SPL_P1|QB1  9.84682784761905e-13
L_PG4_23|_SPL_P1|7 _PG4_23|_SPL_P1|QB1 _PG4_23|P1_COPY_2  2e-12
L_PG4_23|_PG|A1 _PG4_23|P1_COPY_1 _PG4_23|_PG|A1  2.067833848e-12
L_PG4_23|_PG|A2 _PG4_23|_PG|A1 _PG4_23|_PG|A2  4.135667696e-12
L_PG4_23|_PG|A3 _PG4_23|_PG|A3 _PG4_23|_PG|Q3  1.2e-12
L_PG4_23|_PG|B1 _PG4_23|G1_COPY_1 _PG4_23|_PG|B1  2.067833848e-12
L_PG4_23|_PG|B2 _PG4_23|_PG|B1 _PG4_23|_PG|B2  4.135667696e-12
L_PG4_23|_PG|B3 _PG4_23|_PG|B3 _PG4_23|_PG|Q3  1.2e-12
L_PG4_23|_PG|Q3 _PG4_23|_PG|Q3 _PG4_23|_PG|Q2  4.135667696e-12
L_PG4_23|_PG|Q2 _PG4_23|_PG|Q2 _PG4_23|_PG|Q1  4.135667696e-12
L_PG4_23|_PG|Q1 _PG4_23|_PG|Q1 _PG4_23|PG  2.067833848e-12
L_PG4_23|_GG|A1 G3_2_TO4 _PG4_23|_GG|A1  2.067833848e-12
L_PG4_23|_GG|A2 _PG4_23|_GG|A1 _PG4_23|_GG|A2  4.135667696e-12
L_PG4_23|_GG|A3 _PG4_23|_GG|A3 _PG4_23|_GG|Q3  1.2e-12
L_PG4_23|_GG|B1 _PG4_23|G1_COPY_2 _PG4_23|_GG|B1  2.067833848e-12
L_PG4_23|_GG|B2 _PG4_23|_GG|B1 _PG4_23|_GG|B2  4.135667696e-12
L_PG4_23|_GG|B3 _PG4_23|_GG|B3 _PG4_23|_GG|Q3  1.2e-12
L_PG4_23|_GG|Q3 _PG4_23|_GG|Q3 _PG4_23|_GG|Q2  4.135667696e-12
L_PG4_23|_GG|Q2 _PG4_23|_GG|Q2 _PG4_23|_GG|Q1  4.135667696e-12
L_PG4_23|_GG|Q1 _PG4_23|_GG|Q1 _PG4_23|GG  2.067833848e-12
L_PG4_23|_DFF_P0|1 P3_2_TO4 _PG4_23|_DFF_P0|A1  2.067833848e-12
L_PG4_23|_DFF_P0|2 _PG4_23|_DFF_P0|A1 _PG4_23|_DFF_P0|A2  4.135667696e-12
L_PG4_23|_DFF_P0|3 _PG4_23|_DFF_P0|A3 _PG4_23|_DFF_P0|A4  8.271335392e-12
L_PG4_23|_DFF_P0|T T35 _PG4_23|_DFF_P0|T1  2.067833848e-12
L_PG4_23|_DFF_P0|4 _PG4_23|_DFF_P0|T1 _PG4_23|_DFF_P0|T2  4.135667696e-12
L_PG4_23|_DFF_P0|5 _PG4_23|_DFF_P0|A4 _PG4_23|_DFF_P0|Q1  4.135667696e-12
L_PG4_23|_DFF_P0|6 _PG4_23|_DFF_P0|Q1 _PG4_23|P0_SYNC  2.067833848e-12
L_PG4_23|_DFF_P1|1 _PG4_23|P1_COPY_2 _PG4_23|_DFF_P1|A1  2.067833848e-12
L_PG4_23|_DFF_P1|2 _PG4_23|_DFF_P1|A1 _PG4_23|_DFF_P1|A2  4.135667696e-12
L_PG4_23|_DFF_P1|3 _PG4_23|_DFF_P1|A3 _PG4_23|_DFF_P1|A4  8.271335392e-12
L_PG4_23|_DFF_P1|T T35 _PG4_23|_DFF_P1|T1  2.067833848e-12
L_PG4_23|_DFF_P1|4 _PG4_23|_DFF_P1|T1 _PG4_23|_DFF_P1|T2  4.135667696e-12
L_PG4_23|_DFF_P1|5 _PG4_23|_DFF_P1|A4 _PG4_23|_DFF_P1|Q1  4.135667696e-12
L_PG4_23|_DFF_P1|6 _PG4_23|_DFF_P1|Q1 _PG4_23|P1_SYNC  2.067833848e-12
L_PG4_23|_DFF_PG|1 _PG4_23|PG _PG4_23|_DFF_PG|A1  2.067833848e-12
L_PG4_23|_DFF_PG|2 _PG4_23|_DFF_PG|A1 _PG4_23|_DFF_PG|A2  4.135667696e-12
L_PG4_23|_DFF_PG|3 _PG4_23|_DFF_PG|A3 _PG4_23|_DFF_PG|A4  8.271335392e-12
L_PG4_23|_DFF_PG|T T35 _PG4_23|_DFF_PG|T1  2.067833848e-12
L_PG4_23|_DFF_PG|4 _PG4_23|_DFF_PG|T1 _PG4_23|_DFF_PG|T2  4.135667696e-12
L_PG4_23|_DFF_PG|5 _PG4_23|_DFF_PG|A4 _PG4_23|_DFF_PG|Q1  4.135667696e-12
L_PG4_23|_DFF_PG|6 _PG4_23|_DFF_PG|Q1 _PG4_23|PG_SYNC  2.067833848e-12
L_PG4_23|_DFF_GG|1 _PG4_23|GG _PG4_23|_DFF_GG|A1  2.067833848e-12
L_PG4_23|_DFF_GG|2 _PG4_23|_DFF_GG|A1 _PG4_23|_DFF_GG|A2  4.135667696e-12
L_PG4_23|_DFF_GG|3 _PG4_23|_DFF_GG|A3 _PG4_23|_DFF_GG|A4  8.271335392e-12
L_PG4_23|_DFF_GG|T T35 _PG4_23|_DFF_GG|T1  2.067833848e-12
L_PG4_23|_DFF_GG|4 _PG4_23|_DFF_GG|T1 _PG4_23|_DFF_GG|T2  4.135667696e-12
L_PG4_23|_DFF_GG|5 _PG4_23|_DFF_GG|A4 _PG4_23|_DFF_GG|Q1  4.135667696e-12
L_PG4_23|_DFF_GG|6 _PG4_23|_DFF_GG|Q1 _PG4_23|GG_SYNC  2.067833848e-12
L_PG4_23|_AND_G|A1 _PG4_23|PG_SYNC _PG4_23|_AND_G|A1  2.067833848e-12
L_PG4_23|_AND_G|A2 _PG4_23|_AND_G|A1 _PG4_23|_AND_G|A2  4.135667696e-12
L_PG4_23|_AND_G|A3 _PG4_23|_AND_G|A3 _PG4_23|_AND_G|Q3  1.2e-12
L_PG4_23|_AND_G|B1 _PG4_23|GG_SYNC _PG4_23|_AND_G|B1  2.067833848e-12
L_PG4_23|_AND_G|B2 _PG4_23|_AND_G|B1 _PG4_23|_AND_G|B2  4.135667696e-12
L_PG4_23|_AND_G|B3 _PG4_23|_AND_G|B3 _PG4_23|_AND_G|Q3  1.2e-12
L_PG4_23|_AND_G|Q3 _PG4_23|_AND_G|Q3 _PG4_23|_AND_G|Q2  4.135667696e-12
L_PG4_23|_AND_G|Q2 _PG4_23|_AND_G|Q2 _PG4_23|_AND_G|Q1  4.135667696e-12
L_PG4_23|_AND_G|Q1 _PG4_23|_AND_G|Q1 G4_3_TX  2.067833848e-12
L_PG4_23|_AND_P|A1 _PG4_23|P0_SYNC _PG4_23|_AND_P|A1  2.067833848e-12
L_PG4_23|_AND_P|A2 _PG4_23|_AND_P|A1 _PG4_23|_AND_P|A2  4.135667696e-12
L_PG4_23|_AND_P|A3 _PG4_23|_AND_P|A3 _PG4_23|_AND_P|Q3  1.2e-12
L_PG4_23|_AND_P|B1 _PG4_23|P1_SYNC _PG4_23|_AND_P|B1  2.067833848e-12
L_PG4_23|_AND_P|B2 _PG4_23|_AND_P|B1 _PG4_23|_AND_P|B2  4.135667696e-12
L_PG4_23|_AND_P|B3 _PG4_23|_AND_P|B3 _PG4_23|_AND_P|Q3  1.2e-12
L_PG4_23|_AND_P|Q3 _PG4_23|_AND_P|Q3 _PG4_23|_AND_P|Q2  4.135667696e-12
L_PG4_23|_AND_P|Q2 _PG4_23|_AND_P|Q2 _PG4_23|_AND_P|Q1  4.135667696e-12
L_PG4_23|_AND_P|Q1 _PG4_23|_AND_P|Q1 P4_3_TX  2.067833848e-12
L_IP5_23|I_1|B _IP5_23|A1 _IP5_23|I_1|MID  2e-12
I_IP5_23|I_1|B 0 _IP5_23|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP5_23|I_3|B _IP5_23|A3 _IP5_23|I_3|MID  2e-12
I_IP5_23|I_3|B 0 _IP5_23|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP5_23|I_T|B _IP5_23|T1 _IP5_23|I_T|MID  2e-12
I_IP5_23|I_T|B 0 _IP5_23|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP5_23|I_6|B _IP5_23|Q1 _IP5_23|I_6|MID  2e-12
I_IP5_23|I_6|B 0 _IP5_23|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP5_23|1|1 _IP5_23|A1 _IP5_23|1|MID_SERIES JJMIT AREA=2.5
L_IP5_23|1|P _IP5_23|1|MID_SERIES 0  2e-13
R_IP5_23|1|B _IP5_23|A1 _IP5_23|1|MID_SHUNT  2.7439617672
L_IP5_23|1|RB _IP5_23|1|MID_SHUNT 0  1.550338398468e-12
B_IP5_23|23|1 _IP5_23|A2 _IP5_23|A3 JJMIT AREA=1.7857142857142858
R_IP5_23|23|B _IP5_23|A2 _IP5_23|23|MID_SHUNT  3.84154647408
L_IP5_23|23|RB _IP5_23|23|MID_SHUNT _IP5_23|A3  2.1704737578552e-12
B_IP5_23|3|1 _IP5_23|A3 _IP5_23|3|MID_SERIES JJMIT AREA=2.5
L_IP5_23|3|P _IP5_23|3|MID_SERIES 0  2e-13
R_IP5_23|3|B _IP5_23|A3 _IP5_23|3|MID_SHUNT  2.7439617672
L_IP5_23|3|RB _IP5_23|3|MID_SHUNT 0  1.550338398468e-12
B_IP5_23|4|1 _IP5_23|A4 _IP5_23|4|MID_SERIES JJMIT AREA=2.5
L_IP5_23|4|P _IP5_23|4|MID_SERIES 0  2e-13
R_IP5_23|4|B _IP5_23|A4 _IP5_23|4|MID_SHUNT  2.7439617672
L_IP5_23|4|RB _IP5_23|4|MID_SHUNT 0  1.550338398468e-12
B_IP5_23|T|1 _IP5_23|T1 _IP5_23|T|MID_SERIES JJMIT AREA=2.5
L_IP5_23|T|P _IP5_23|T|MID_SERIES 0  2e-13
R_IP5_23|T|B _IP5_23|T1 _IP5_23|T|MID_SHUNT  2.7439617672
L_IP5_23|T|RB _IP5_23|T|MID_SHUNT 0  1.550338398468e-12
B_IP5_23|45|1 _IP5_23|T2 _IP5_23|A4 JJMIT AREA=1.7857142857142858
R_IP5_23|45|B _IP5_23|T2 _IP5_23|45|MID_SHUNT  3.84154647408
L_IP5_23|45|RB _IP5_23|45|MID_SHUNT _IP5_23|A4  2.1704737578552e-12
B_IP5_23|6|1 _IP5_23|Q1 _IP5_23|6|MID_SERIES JJMIT AREA=2.5
L_IP5_23|6|P _IP5_23|6|MID_SERIES 0  2e-13
R_IP5_23|6|B _IP5_23|Q1 _IP5_23|6|MID_SHUNT  2.7439617672
L_IP5_23|6|RB _IP5_23|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_SPL_G1|1 G5_2_TO5 _PG5_23|_SPL_G1|D1  2e-12
L_PG5_23|_SPL_G1|2 _PG5_23|_SPL_G1|D1 _PG5_23|_SPL_G1|D2  4.135667696e-12
L_PG5_23|_SPL_G1|3 _PG5_23|_SPL_G1|D2 _PG5_23|_SPL_G1|JCT  9.84682784761905e-13
L_PG5_23|_SPL_G1|4 _PG5_23|_SPL_G1|JCT _PG5_23|_SPL_G1|QA1  9.84682784761905e-13
L_PG5_23|_SPL_G1|5 _PG5_23|_SPL_G1|QA1 _PG5_23|G1_COPY_1  2e-12
L_PG5_23|_SPL_G1|6 _PG5_23|_SPL_G1|JCT _PG5_23|_SPL_G1|QB1  9.84682784761905e-13
L_PG5_23|_SPL_G1|7 _PG5_23|_SPL_G1|QB1 _PG5_23|G1_COPY_2  2e-12
L_PG5_23|_SPL_P1|1 P5_2_TO5 _PG5_23|_SPL_P1|D1  2e-12
L_PG5_23|_SPL_P1|2 _PG5_23|_SPL_P1|D1 _PG5_23|_SPL_P1|D2  4.135667696e-12
L_PG5_23|_SPL_P1|3 _PG5_23|_SPL_P1|D2 _PG5_23|_SPL_P1|JCT  9.84682784761905e-13
L_PG5_23|_SPL_P1|4 _PG5_23|_SPL_P1|JCT _PG5_23|_SPL_P1|QA1  9.84682784761905e-13
L_PG5_23|_SPL_P1|5 _PG5_23|_SPL_P1|QA1 _PG5_23|P1_COPY_1  2e-12
L_PG5_23|_SPL_P1|6 _PG5_23|_SPL_P1|JCT _PG5_23|_SPL_P1|QB1  9.84682784761905e-13
L_PG5_23|_SPL_P1|7 _PG5_23|_SPL_P1|QB1 _PG5_23|P1_COPY_2  2e-12
L_PG5_23|_PG|A1 _PG5_23|P1_COPY_1 _PG5_23|_PG|A1  2.067833848e-12
L_PG5_23|_PG|A2 _PG5_23|_PG|A1 _PG5_23|_PG|A2  4.135667696e-12
L_PG5_23|_PG|A3 _PG5_23|_PG|A3 _PG5_23|_PG|Q3  1.2e-12
L_PG5_23|_PG|B1 _PG5_23|G1_COPY_1 _PG5_23|_PG|B1  2.067833848e-12
L_PG5_23|_PG|B2 _PG5_23|_PG|B1 _PG5_23|_PG|B2  4.135667696e-12
L_PG5_23|_PG|B3 _PG5_23|_PG|B3 _PG5_23|_PG|Q3  1.2e-12
L_PG5_23|_PG|Q3 _PG5_23|_PG|Q3 _PG5_23|_PG|Q2  4.135667696e-12
L_PG5_23|_PG|Q2 _PG5_23|_PG|Q2 _PG5_23|_PG|Q1  4.135667696e-12
L_PG5_23|_PG|Q1 _PG5_23|_PG|Q1 _PG5_23|PG  2.067833848e-12
L_PG5_23|_GG|A1 G3_2_TO5 _PG5_23|_GG|A1  2.067833848e-12
L_PG5_23|_GG|A2 _PG5_23|_GG|A1 _PG5_23|_GG|A2  4.135667696e-12
L_PG5_23|_GG|A3 _PG5_23|_GG|A3 _PG5_23|_GG|Q3  1.2e-12
L_PG5_23|_GG|B1 _PG5_23|G1_COPY_2 _PG5_23|_GG|B1  2.067833848e-12
L_PG5_23|_GG|B2 _PG5_23|_GG|B1 _PG5_23|_GG|B2  4.135667696e-12
L_PG5_23|_GG|B3 _PG5_23|_GG|B3 _PG5_23|_GG|Q3  1.2e-12
L_PG5_23|_GG|Q3 _PG5_23|_GG|Q3 _PG5_23|_GG|Q2  4.135667696e-12
L_PG5_23|_GG|Q2 _PG5_23|_GG|Q2 _PG5_23|_GG|Q1  4.135667696e-12
L_PG5_23|_GG|Q1 _PG5_23|_GG|Q1 _PG5_23|GG  2.067833848e-12
L_PG5_23|_DFF_P0|1 P3_2_TO5 _PG5_23|_DFF_P0|A1  2.067833848e-12
L_PG5_23|_DFF_P0|2 _PG5_23|_DFF_P0|A1 _PG5_23|_DFF_P0|A2  4.135667696e-12
L_PG5_23|_DFF_P0|3 _PG5_23|_DFF_P0|A3 _PG5_23|_DFF_P0|A4  8.271335392e-12
L_PG5_23|_DFF_P0|T T37 _PG5_23|_DFF_P0|T1  2.067833848e-12
L_PG5_23|_DFF_P0|4 _PG5_23|_DFF_P0|T1 _PG5_23|_DFF_P0|T2  4.135667696e-12
L_PG5_23|_DFF_P0|5 _PG5_23|_DFF_P0|A4 _PG5_23|_DFF_P0|Q1  4.135667696e-12
L_PG5_23|_DFF_P0|6 _PG5_23|_DFF_P0|Q1 _PG5_23|P0_SYNC  2.067833848e-12
L_PG5_23|_DFF_P1|1 _PG5_23|P1_COPY_2 _PG5_23|_DFF_P1|A1  2.067833848e-12
L_PG5_23|_DFF_P1|2 _PG5_23|_DFF_P1|A1 _PG5_23|_DFF_P1|A2  4.135667696e-12
L_PG5_23|_DFF_P1|3 _PG5_23|_DFF_P1|A3 _PG5_23|_DFF_P1|A4  8.271335392e-12
L_PG5_23|_DFF_P1|T T37 _PG5_23|_DFF_P1|T1  2.067833848e-12
L_PG5_23|_DFF_P1|4 _PG5_23|_DFF_P1|T1 _PG5_23|_DFF_P1|T2  4.135667696e-12
L_PG5_23|_DFF_P1|5 _PG5_23|_DFF_P1|A4 _PG5_23|_DFF_P1|Q1  4.135667696e-12
L_PG5_23|_DFF_P1|6 _PG5_23|_DFF_P1|Q1 _PG5_23|P1_SYNC  2.067833848e-12
L_PG5_23|_DFF_PG|1 _PG5_23|PG _PG5_23|_DFF_PG|A1  2.067833848e-12
L_PG5_23|_DFF_PG|2 _PG5_23|_DFF_PG|A1 _PG5_23|_DFF_PG|A2  4.135667696e-12
L_PG5_23|_DFF_PG|3 _PG5_23|_DFF_PG|A3 _PG5_23|_DFF_PG|A4  8.271335392e-12
L_PG5_23|_DFF_PG|T T37 _PG5_23|_DFF_PG|T1  2.067833848e-12
L_PG5_23|_DFF_PG|4 _PG5_23|_DFF_PG|T1 _PG5_23|_DFF_PG|T2  4.135667696e-12
L_PG5_23|_DFF_PG|5 _PG5_23|_DFF_PG|A4 _PG5_23|_DFF_PG|Q1  4.135667696e-12
L_PG5_23|_DFF_PG|6 _PG5_23|_DFF_PG|Q1 _PG5_23|PG_SYNC  2.067833848e-12
L_PG5_23|_DFF_GG|1 _PG5_23|GG _PG5_23|_DFF_GG|A1  2.067833848e-12
L_PG5_23|_DFF_GG|2 _PG5_23|_DFF_GG|A1 _PG5_23|_DFF_GG|A2  4.135667696e-12
L_PG5_23|_DFF_GG|3 _PG5_23|_DFF_GG|A3 _PG5_23|_DFF_GG|A4  8.271335392e-12
L_PG5_23|_DFF_GG|T T37 _PG5_23|_DFF_GG|T1  2.067833848e-12
L_PG5_23|_DFF_GG|4 _PG5_23|_DFF_GG|T1 _PG5_23|_DFF_GG|T2  4.135667696e-12
L_PG5_23|_DFF_GG|5 _PG5_23|_DFF_GG|A4 _PG5_23|_DFF_GG|Q1  4.135667696e-12
L_PG5_23|_DFF_GG|6 _PG5_23|_DFF_GG|Q1 _PG5_23|GG_SYNC  2.067833848e-12
L_PG5_23|_AND_G|A1 _PG5_23|PG_SYNC _PG5_23|_AND_G|A1  2.067833848e-12
L_PG5_23|_AND_G|A2 _PG5_23|_AND_G|A1 _PG5_23|_AND_G|A2  4.135667696e-12
L_PG5_23|_AND_G|A3 _PG5_23|_AND_G|A3 _PG5_23|_AND_G|Q3  1.2e-12
L_PG5_23|_AND_G|B1 _PG5_23|GG_SYNC _PG5_23|_AND_G|B1  2.067833848e-12
L_PG5_23|_AND_G|B2 _PG5_23|_AND_G|B1 _PG5_23|_AND_G|B2  4.135667696e-12
L_PG5_23|_AND_G|B3 _PG5_23|_AND_G|B3 _PG5_23|_AND_G|Q3  1.2e-12
L_PG5_23|_AND_G|Q3 _PG5_23|_AND_G|Q3 _PG5_23|_AND_G|Q2  4.135667696e-12
L_PG5_23|_AND_G|Q2 _PG5_23|_AND_G|Q2 _PG5_23|_AND_G|Q1  4.135667696e-12
L_PG5_23|_AND_G|Q1 _PG5_23|_AND_G|Q1 G5_3_TX  2.067833848e-12
L_PG5_23|_AND_P|A1 _PG5_23|P0_SYNC _PG5_23|_AND_P|A1  2.067833848e-12
L_PG5_23|_AND_P|A2 _PG5_23|_AND_P|A1 _PG5_23|_AND_P|A2  4.135667696e-12
L_PG5_23|_AND_P|A3 _PG5_23|_AND_P|A3 _PG5_23|_AND_P|Q3  1.2e-12
L_PG5_23|_AND_P|B1 _PG5_23|P1_SYNC _PG5_23|_AND_P|B1  2.067833848e-12
L_PG5_23|_AND_P|B2 _PG5_23|_AND_P|B1 _PG5_23|_AND_P|B2  4.135667696e-12
L_PG5_23|_AND_P|B3 _PG5_23|_AND_P|B3 _PG5_23|_AND_P|Q3  1.2e-12
L_PG5_23|_AND_P|Q3 _PG5_23|_AND_P|Q3 _PG5_23|_AND_P|Q2  4.135667696e-12
L_PG5_23|_AND_P|Q2 _PG5_23|_AND_P|Q2 _PG5_23|_AND_P|Q1  4.135667696e-12
L_PG5_23|_AND_P|Q1 _PG5_23|_AND_P|Q1 P5_3_TX  2.067833848e-12
L_PG6_23|P|1 P6_2_TO6 _PG6_23|P|A1  2.067833848e-12
L_PG6_23|P|2 _PG6_23|P|A1 _PG6_23|P|A2  4.135667696e-12
L_PG6_23|P|3 _PG6_23|P|A3 _PG6_23|P|A4  8.271335392e-12
L_PG6_23|P|T T38 _PG6_23|P|T1  2.067833848e-12
L_PG6_23|P|4 _PG6_23|P|T1 _PG6_23|P|T2  4.135667696e-12
L_PG6_23|P|5 _PG6_23|P|A4 _PG6_23|P|Q1  4.135667696e-12
L_PG6_23|P|6 _PG6_23|P|Q1 P6_3_TX  2.067833848e-12
L_PG6_23|G|1 G6_2_TO6 _PG6_23|G|A1  2.067833848e-12
L_PG6_23|G|2 _PG6_23|G|A1 _PG6_23|G|A2  4.135667696e-12
L_PG6_23|G|3 _PG6_23|G|A3 _PG6_23|G|A4  8.271335392e-12
L_PG6_23|G|T T38 _PG6_23|G|T1  2.067833848e-12
L_PG6_23|G|4 _PG6_23|G|T1 _PG6_23|G|T2  4.135667696e-12
L_PG6_23|G|5 _PG6_23|G|A4 _PG6_23|G|Q1  4.135667696e-12
L_PG6_23|G|6 _PG6_23|G|Q1 G6_3_TX  2.067833848e-12
L_IP7_23|I_1|B _IP7_23|A1 _IP7_23|I_1|MID  2e-12
I_IP7_23|I_1|B 0 _IP7_23|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP7_23|I_3|B _IP7_23|A3 _IP7_23|I_3|MID  2e-12
I_IP7_23|I_3|B 0 _IP7_23|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP7_23|I_T|B _IP7_23|T1 _IP7_23|I_T|MID  2e-12
I_IP7_23|I_T|B 0 _IP7_23|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP7_23|I_6|B _IP7_23|Q1 _IP7_23|I_6|MID  2e-12
I_IP7_23|I_6|B 0 _IP7_23|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP7_23|1|1 _IP7_23|A1 _IP7_23|1|MID_SERIES JJMIT AREA=2.5
L_IP7_23|1|P _IP7_23|1|MID_SERIES 0  2e-13
R_IP7_23|1|B _IP7_23|A1 _IP7_23|1|MID_SHUNT  2.7439617672
L_IP7_23|1|RB _IP7_23|1|MID_SHUNT 0  1.550338398468e-12
B_IP7_23|23|1 _IP7_23|A2 _IP7_23|A3 JJMIT AREA=1.7857142857142858
R_IP7_23|23|B _IP7_23|A2 _IP7_23|23|MID_SHUNT  3.84154647408
L_IP7_23|23|RB _IP7_23|23|MID_SHUNT _IP7_23|A3  2.1704737578552e-12
B_IP7_23|3|1 _IP7_23|A3 _IP7_23|3|MID_SERIES JJMIT AREA=2.5
L_IP7_23|3|P _IP7_23|3|MID_SERIES 0  2e-13
R_IP7_23|3|B _IP7_23|A3 _IP7_23|3|MID_SHUNT  2.7439617672
L_IP7_23|3|RB _IP7_23|3|MID_SHUNT 0  1.550338398468e-12
B_IP7_23|4|1 _IP7_23|A4 _IP7_23|4|MID_SERIES JJMIT AREA=2.5
L_IP7_23|4|P _IP7_23|4|MID_SERIES 0  2e-13
R_IP7_23|4|B _IP7_23|A4 _IP7_23|4|MID_SHUNT  2.7439617672
L_IP7_23|4|RB _IP7_23|4|MID_SHUNT 0  1.550338398468e-12
B_IP7_23|T|1 _IP7_23|T1 _IP7_23|T|MID_SERIES JJMIT AREA=2.5
L_IP7_23|T|P _IP7_23|T|MID_SERIES 0  2e-13
R_IP7_23|T|B _IP7_23|T1 _IP7_23|T|MID_SHUNT  2.7439617672
L_IP7_23|T|RB _IP7_23|T|MID_SHUNT 0  1.550338398468e-12
B_IP7_23|45|1 _IP7_23|T2 _IP7_23|A4 JJMIT AREA=1.7857142857142858
R_IP7_23|45|B _IP7_23|T2 _IP7_23|45|MID_SHUNT  3.84154647408
L_IP7_23|45|RB _IP7_23|45|MID_SHUNT _IP7_23|A4  2.1704737578552e-12
B_IP7_23|6|1 _IP7_23|Q1 _IP7_23|6|MID_SERIES JJMIT AREA=2.5
L_IP7_23|6|P _IP7_23|6|MID_SERIES 0  2e-13
R_IP7_23|6|B _IP7_23|Q1 _IP7_23|6|MID_SHUNT  2.7439617672
L_IP7_23|6|RB _IP7_23|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_SPL_G1|1 G7_2_TO7 _PG7_23|_SPL_G1|D1  2e-12
L_PG7_23|_SPL_G1|2 _PG7_23|_SPL_G1|D1 _PG7_23|_SPL_G1|D2  4.135667696e-12
L_PG7_23|_SPL_G1|3 _PG7_23|_SPL_G1|D2 _PG7_23|_SPL_G1|JCT  9.84682784761905e-13
L_PG7_23|_SPL_G1|4 _PG7_23|_SPL_G1|JCT _PG7_23|_SPL_G1|QA1  9.84682784761905e-13
L_PG7_23|_SPL_G1|5 _PG7_23|_SPL_G1|QA1 _PG7_23|G1_COPY_1  2e-12
L_PG7_23|_SPL_G1|6 _PG7_23|_SPL_G1|JCT _PG7_23|_SPL_G1|QB1  9.84682784761905e-13
L_PG7_23|_SPL_G1|7 _PG7_23|_SPL_G1|QB1 _PG7_23|G1_COPY_2  2e-12
L_PG7_23|_SPL_P1|1 P7_2_TO7 _PG7_23|_SPL_P1|D1  2e-12
L_PG7_23|_SPL_P1|2 _PG7_23|_SPL_P1|D1 _PG7_23|_SPL_P1|D2  4.135667696e-12
L_PG7_23|_SPL_P1|3 _PG7_23|_SPL_P1|D2 _PG7_23|_SPL_P1|JCT  9.84682784761905e-13
L_PG7_23|_SPL_P1|4 _PG7_23|_SPL_P1|JCT _PG7_23|_SPL_P1|QA1  9.84682784761905e-13
L_PG7_23|_SPL_P1|5 _PG7_23|_SPL_P1|QA1 _PG7_23|P1_COPY_1  2e-12
L_PG7_23|_SPL_P1|6 _PG7_23|_SPL_P1|JCT _PG7_23|_SPL_P1|QB1  9.84682784761905e-13
L_PG7_23|_SPL_P1|7 _PG7_23|_SPL_P1|QB1 _PG7_23|P1_COPY_2  2e-12
L_PG7_23|_PG|A1 _PG7_23|P1_COPY_1 _PG7_23|_PG|A1  2.067833848e-12
L_PG7_23|_PG|A2 _PG7_23|_PG|A1 _PG7_23|_PG|A2  4.135667696e-12
L_PG7_23|_PG|A3 _PG7_23|_PG|A3 _PG7_23|_PG|Q3  1.2e-12
L_PG7_23|_PG|B1 _PG7_23|G1_COPY_1 _PG7_23|_PG|B1  2.067833848e-12
L_PG7_23|_PG|B2 _PG7_23|_PG|B1 _PG7_23|_PG|B2  4.135667696e-12
L_PG7_23|_PG|B3 _PG7_23|_PG|B3 _PG7_23|_PG|Q3  1.2e-12
L_PG7_23|_PG|Q3 _PG7_23|_PG|Q3 _PG7_23|_PG|Q2  4.135667696e-12
L_PG7_23|_PG|Q2 _PG7_23|_PG|Q2 _PG7_23|_PG|Q1  4.135667696e-12
L_PG7_23|_PG|Q1 _PG7_23|_PG|Q1 _PG7_23|PG  2.067833848e-12
L_PG7_23|_GG|A1 G3_2_TO7 _PG7_23|_GG|A1  2.067833848e-12
L_PG7_23|_GG|A2 _PG7_23|_GG|A1 _PG7_23|_GG|A2  4.135667696e-12
L_PG7_23|_GG|A3 _PG7_23|_GG|A3 _PG7_23|_GG|Q3  1.2e-12
L_PG7_23|_GG|B1 _PG7_23|G1_COPY_2 _PG7_23|_GG|B1  2.067833848e-12
L_PG7_23|_GG|B2 _PG7_23|_GG|B1 _PG7_23|_GG|B2  4.135667696e-12
L_PG7_23|_GG|B3 _PG7_23|_GG|B3 _PG7_23|_GG|Q3  1.2e-12
L_PG7_23|_GG|Q3 _PG7_23|_GG|Q3 _PG7_23|_GG|Q2  4.135667696e-12
L_PG7_23|_GG|Q2 _PG7_23|_GG|Q2 _PG7_23|_GG|Q1  4.135667696e-12
L_PG7_23|_GG|Q1 _PG7_23|_GG|Q1 _PG7_23|GG  2.067833848e-12
L_PG7_23|_DFF_P0|1 P3_2_TO7 _PG7_23|_DFF_P0|A1  2.067833848e-12
L_PG7_23|_DFF_P0|2 _PG7_23|_DFF_P0|A1 _PG7_23|_DFF_P0|A2  4.135667696e-12
L_PG7_23|_DFF_P0|3 _PG7_23|_DFF_P0|A3 _PG7_23|_DFF_P0|A4  8.271335392e-12
L_PG7_23|_DFF_P0|T T3A _PG7_23|_DFF_P0|T1  2.067833848e-12
L_PG7_23|_DFF_P0|4 _PG7_23|_DFF_P0|T1 _PG7_23|_DFF_P0|T2  4.135667696e-12
L_PG7_23|_DFF_P0|5 _PG7_23|_DFF_P0|A4 _PG7_23|_DFF_P0|Q1  4.135667696e-12
L_PG7_23|_DFF_P0|6 _PG7_23|_DFF_P0|Q1 _PG7_23|P0_SYNC  2.067833848e-12
L_PG7_23|_DFF_P1|1 _PG7_23|P1_COPY_2 _PG7_23|_DFF_P1|A1  2.067833848e-12
L_PG7_23|_DFF_P1|2 _PG7_23|_DFF_P1|A1 _PG7_23|_DFF_P1|A2  4.135667696e-12
L_PG7_23|_DFF_P1|3 _PG7_23|_DFF_P1|A3 _PG7_23|_DFF_P1|A4  8.271335392e-12
L_PG7_23|_DFF_P1|T T3A _PG7_23|_DFF_P1|T1  2.067833848e-12
L_PG7_23|_DFF_P1|4 _PG7_23|_DFF_P1|T1 _PG7_23|_DFF_P1|T2  4.135667696e-12
L_PG7_23|_DFF_P1|5 _PG7_23|_DFF_P1|A4 _PG7_23|_DFF_P1|Q1  4.135667696e-12
L_PG7_23|_DFF_P1|6 _PG7_23|_DFF_P1|Q1 _PG7_23|P1_SYNC  2.067833848e-12
L_PG7_23|_DFF_PG|1 _PG7_23|PG _PG7_23|_DFF_PG|A1  2.067833848e-12
L_PG7_23|_DFF_PG|2 _PG7_23|_DFF_PG|A1 _PG7_23|_DFF_PG|A2  4.135667696e-12
L_PG7_23|_DFF_PG|3 _PG7_23|_DFF_PG|A3 _PG7_23|_DFF_PG|A4  8.271335392e-12
L_PG7_23|_DFF_PG|T T3A _PG7_23|_DFF_PG|T1  2.067833848e-12
L_PG7_23|_DFF_PG|4 _PG7_23|_DFF_PG|T1 _PG7_23|_DFF_PG|T2  4.135667696e-12
L_PG7_23|_DFF_PG|5 _PG7_23|_DFF_PG|A4 _PG7_23|_DFF_PG|Q1  4.135667696e-12
L_PG7_23|_DFF_PG|6 _PG7_23|_DFF_PG|Q1 _PG7_23|PG_SYNC  2.067833848e-12
L_PG7_23|_DFF_GG|1 _PG7_23|GG _PG7_23|_DFF_GG|A1  2.067833848e-12
L_PG7_23|_DFF_GG|2 _PG7_23|_DFF_GG|A1 _PG7_23|_DFF_GG|A2  4.135667696e-12
L_PG7_23|_DFF_GG|3 _PG7_23|_DFF_GG|A3 _PG7_23|_DFF_GG|A4  8.271335392e-12
L_PG7_23|_DFF_GG|T T3A _PG7_23|_DFF_GG|T1  2.067833848e-12
L_PG7_23|_DFF_GG|4 _PG7_23|_DFF_GG|T1 _PG7_23|_DFF_GG|T2  4.135667696e-12
L_PG7_23|_DFF_GG|5 _PG7_23|_DFF_GG|A4 _PG7_23|_DFF_GG|Q1  4.135667696e-12
L_PG7_23|_DFF_GG|6 _PG7_23|_DFF_GG|Q1 _PG7_23|GG_SYNC  2.067833848e-12
L_PG7_23|_AND_G|A1 _PG7_23|PG_SYNC _PG7_23|_AND_G|A1  2.067833848e-12
L_PG7_23|_AND_G|A2 _PG7_23|_AND_G|A1 _PG7_23|_AND_G|A2  4.135667696e-12
L_PG7_23|_AND_G|A3 _PG7_23|_AND_G|A3 _PG7_23|_AND_G|Q3  1.2e-12
L_PG7_23|_AND_G|B1 _PG7_23|GG_SYNC _PG7_23|_AND_G|B1  2.067833848e-12
L_PG7_23|_AND_G|B2 _PG7_23|_AND_G|B1 _PG7_23|_AND_G|B2  4.135667696e-12
L_PG7_23|_AND_G|B3 _PG7_23|_AND_G|B3 _PG7_23|_AND_G|Q3  1.2e-12
L_PG7_23|_AND_G|Q3 _PG7_23|_AND_G|Q3 _PG7_23|_AND_G|Q2  4.135667696e-12
L_PG7_23|_AND_G|Q2 _PG7_23|_AND_G|Q2 _PG7_23|_AND_G|Q1  4.135667696e-12
L_PG7_23|_AND_G|Q1 _PG7_23|_AND_G|Q1 S8_3_TX  2.067833848e-12
L_PG7_23|_AND_P|A1 _PG7_23|P0_SYNC _PG7_23|_AND_P|A1  2.067833848e-12
L_PG7_23|_AND_P|A2 _PG7_23|_AND_P|A1 _PG7_23|_AND_P|A2  4.135667696e-12
L_PG7_23|_AND_P|A3 _PG7_23|_AND_P|A3 _PG7_23|_AND_P|Q3  1.2e-12
L_PG7_23|_AND_P|B1 _PG7_23|P1_SYNC _PG7_23|_AND_P|B1  2.067833848e-12
L_PG7_23|_AND_P|B2 _PG7_23|_AND_P|B1 _PG7_23|_AND_P|B2  4.135667696e-12
L_PG7_23|_AND_P|B3 _PG7_23|_AND_P|B3 _PG7_23|_AND_P|Q3  1.2e-12
L_PG7_23|_AND_P|Q3 _PG7_23|_AND_P|Q3 _PG7_23|_AND_P|Q2  4.135667696e-12
L_PG7_23|_AND_P|Q2 _PG7_23|_AND_P|Q2 _PG7_23|_AND_P|Q1  4.135667696e-12
L_PG7_23|_AND_P|Q1 _PG7_23|_AND_P|Q1 P7_3_TX  2.067833848e-12
B_PTL_S0_3|_TX|1 _PTL_S0_3|_TX|1 _PTL_S0_3|_TX|2 JJMIT AREA=2.5
B_PTL_S0_3|_TX|2 _PTL_S0_3|_TX|4 _PTL_S0_3|_TX|5 JJMIT AREA=2.5
I_PTL_S0_3|_TX|B1 0 _PTL_S0_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S0_3|_TX|B2 0 _PTL_S0_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S0_3|_TX|B1 _PTL_S0_3|_TX|1 _PTL_S0_3|_TX|3  1.684e-12
L_PTL_S0_3|_TX|B2 _PTL_S0_3|_TX|4 _PTL_S0_3|_TX|6  3.596e-12
L_PTL_S0_3|_TX|1 S0_3_TX _PTL_S0_3|_TX|1  2.063e-12
L_PTL_S0_3|_TX|2 _PTL_S0_3|_TX|1 _PTL_S0_3|_TX|4  4.123e-12
L_PTL_S0_3|_TX|3 _PTL_S0_3|_TX|4 _PTL_S0_3|_TX|7  2.193e-12
R_PTL_S0_3|_TX|D _PTL_S0_3|_TX|7 _PTL_S0_3|A_PTL  1.36
L_PTL_S0_3|_TX|P1 _PTL_S0_3|_TX|2 0  5.254e-13
L_PTL_S0_3|_TX|P2 _PTL_S0_3|_TX|5 0  5.141e-13
R_PTL_S0_3|_TX|B1 _PTL_S0_3|_TX|1 _PTL_S0_3|_TX|101  2.7439617672
R_PTL_S0_3|_TX|B2 _PTL_S0_3|_TX|4 _PTL_S0_3|_TX|104  2.7439617672
L_PTL_S0_3|_TX|RB1 _PTL_S0_3|_TX|101 0  1.550338398468e-12
L_PTL_S0_3|_TX|RB2 _PTL_S0_3|_TX|104 0  1.550338398468e-12
B_PTL_S0_3|_RX|1 _PTL_S0_3|_RX|1 _PTL_S0_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S0_3|_RX|2 _PTL_S0_3|_RX|4 _PTL_S0_3|_RX|5 JJMIT AREA=2.0
B_PTL_S0_3|_RX|3 _PTL_S0_3|_RX|7 _PTL_S0_3|_RX|8 JJMIT AREA=2.5
I_PTL_S0_3|_RX|B1 0 _PTL_S0_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S0_3|_RX|B1 _PTL_S0_3|_RX|1 _PTL_S0_3|_RX|3  2.777e-12
I_PTL_S0_3|_RX|B2 0 _PTL_S0_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S0_3|_RX|B2 _PTL_S0_3|_RX|4 _PTL_S0_3|_RX|6  2.685e-12
I_PTL_S0_3|_RX|B3 0 _PTL_S0_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S0_3|_RX|B3 _PTL_S0_3|_RX|7 _PTL_S0_3|_RX|9  2.764e-12
L_PTL_S0_3|_RX|1 _PTL_S0_3|A_PTL _PTL_S0_3|_RX|1  1.346e-12
L_PTL_S0_3|_RX|2 _PTL_S0_3|_RX|1 _PTL_S0_3|_RX|4  6.348e-12
L_PTL_S0_3|_RX|3 _PTL_S0_3|_RX|4 _PTL_S0_3|_RX|7  5.197e-12
L_PTL_S0_3|_RX|4 _PTL_S0_3|_RX|7 S0_3  2.058e-12
L_PTL_S0_3|_RX|P1 _PTL_S0_3|_RX|2 0  4.795e-13
L_PTL_S0_3|_RX|P2 _PTL_S0_3|_RX|5 0  5.431e-13
L_PTL_S0_3|_RX|P3 _PTL_S0_3|_RX|8 0  5.339e-13
R_PTL_S0_3|_RX|B1 _PTL_S0_3|_RX|1 _PTL_S0_3|_RX|101  4.225701121488
R_PTL_S0_3|_RX|B2 _PTL_S0_3|_RX|4 _PTL_S0_3|_RX|104  3.429952209
R_PTL_S0_3|_RX|B3 _PTL_S0_3|_RX|7 _PTL_S0_3|_RX|107  2.7439617672
L_PTL_S0_3|_RX|RB1 _PTL_S0_3|_RX|101 0  2.38752113364072e-12
L_PTL_S0_3|_RX|RB2 _PTL_S0_3|_RX|104 0  1.937922998085e-12
L_PTL_S0_3|_RX|RB3 _PTL_S0_3|_RX|107 0  1.550338398468e-12
B_PTL_S1_3|_TX|1 _PTL_S1_3|_TX|1 _PTL_S1_3|_TX|2 JJMIT AREA=2.5
B_PTL_S1_3|_TX|2 _PTL_S1_3|_TX|4 _PTL_S1_3|_TX|5 JJMIT AREA=2.5
I_PTL_S1_3|_TX|B1 0 _PTL_S1_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S1_3|_TX|B2 0 _PTL_S1_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S1_3|_TX|B1 _PTL_S1_3|_TX|1 _PTL_S1_3|_TX|3  1.684e-12
L_PTL_S1_3|_TX|B2 _PTL_S1_3|_TX|4 _PTL_S1_3|_TX|6  3.596e-12
L_PTL_S1_3|_TX|1 S1_3_TX _PTL_S1_3|_TX|1  2.063e-12
L_PTL_S1_3|_TX|2 _PTL_S1_3|_TX|1 _PTL_S1_3|_TX|4  4.123e-12
L_PTL_S1_3|_TX|3 _PTL_S1_3|_TX|4 _PTL_S1_3|_TX|7  2.193e-12
R_PTL_S1_3|_TX|D _PTL_S1_3|_TX|7 _PTL_S1_3|A_PTL  1.36
L_PTL_S1_3|_TX|P1 _PTL_S1_3|_TX|2 0  5.254e-13
L_PTL_S1_3|_TX|P2 _PTL_S1_3|_TX|5 0  5.141e-13
R_PTL_S1_3|_TX|B1 _PTL_S1_3|_TX|1 _PTL_S1_3|_TX|101  2.7439617672
R_PTL_S1_3|_TX|B2 _PTL_S1_3|_TX|4 _PTL_S1_3|_TX|104  2.7439617672
L_PTL_S1_3|_TX|RB1 _PTL_S1_3|_TX|101 0  1.550338398468e-12
L_PTL_S1_3|_TX|RB2 _PTL_S1_3|_TX|104 0  1.550338398468e-12
B_PTL_S1_3|_RX|1 _PTL_S1_3|_RX|1 _PTL_S1_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S1_3|_RX|2 _PTL_S1_3|_RX|4 _PTL_S1_3|_RX|5 JJMIT AREA=2.0
B_PTL_S1_3|_RX|3 _PTL_S1_3|_RX|7 _PTL_S1_3|_RX|8 JJMIT AREA=2.5
I_PTL_S1_3|_RX|B1 0 _PTL_S1_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S1_3|_RX|B1 _PTL_S1_3|_RX|1 _PTL_S1_3|_RX|3  2.777e-12
I_PTL_S1_3|_RX|B2 0 _PTL_S1_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S1_3|_RX|B2 _PTL_S1_3|_RX|4 _PTL_S1_3|_RX|6  2.685e-12
I_PTL_S1_3|_RX|B3 0 _PTL_S1_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S1_3|_RX|B3 _PTL_S1_3|_RX|7 _PTL_S1_3|_RX|9  2.764e-12
L_PTL_S1_3|_RX|1 _PTL_S1_3|A_PTL _PTL_S1_3|_RX|1  1.346e-12
L_PTL_S1_3|_RX|2 _PTL_S1_3|_RX|1 _PTL_S1_3|_RX|4  6.348e-12
L_PTL_S1_3|_RX|3 _PTL_S1_3|_RX|4 _PTL_S1_3|_RX|7  5.197e-12
L_PTL_S1_3|_RX|4 _PTL_S1_3|_RX|7 S1_3  2.058e-12
L_PTL_S1_3|_RX|P1 _PTL_S1_3|_RX|2 0  4.795e-13
L_PTL_S1_3|_RX|P2 _PTL_S1_3|_RX|5 0  5.431e-13
L_PTL_S1_3|_RX|P3 _PTL_S1_3|_RX|8 0  5.339e-13
R_PTL_S1_3|_RX|B1 _PTL_S1_3|_RX|1 _PTL_S1_3|_RX|101  4.225701121488
R_PTL_S1_3|_RX|B2 _PTL_S1_3|_RX|4 _PTL_S1_3|_RX|104  3.429952209
R_PTL_S1_3|_RX|B3 _PTL_S1_3|_RX|7 _PTL_S1_3|_RX|107  2.7439617672
L_PTL_S1_3|_RX|RB1 _PTL_S1_3|_RX|101 0  2.38752113364072e-12
L_PTL_S1_3|_RX|RB2 _PTL_S1_3|_RX|104 0  1.937922998085e-12
L_PTL_S1_3|_RX|RB3 _PTL_S1_3|_RX|107 0  1.550338398468e-12
B_PTL_S2_3|_TX|1 _PTL_S2_3|_TX|1 _PTL_S2_3|_TX|2 JJMIT AREA=2.5
B_PTL_S2_3|_TX|2 _PTL_S2_3|_TX|4 _PTL_S2_3|_TX|5 JJMIT AREA=2.5
I_PTL_S2_3|_TX|B1 0 _PTL_S2_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S2_3|_TX|B2 0 _PTL_S2_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S2_3|_TX|B1 _PTL_S2_3|_TX|1 _PTL_S2_3|_TX|3  1.684e-12
L_PTL_S2_3|_TX|B2 _PTL_S2_3|_TX|4 _PTL_S2_3|_TX|6  3.596e-12
L_PTL_S2_3|_TX|1 S2_3_TX _PTL_S2_3|_TX|1  2.063e-12
L_PTL_S2_3|_TX|2 _PTL_S2_3|_TX|1 _PTL_S2_3|_TX|4  4.123e-12
L_PTL_S2_3|_TX|3 _PTL_S2_3|_TX|4 _PTL_S2_3|_TX|7  2.193e-12
R_PTL_S2_3|_TX|D _PTL_S2_3|_TX|7 _PTL_S2_3|A_PTL  1.36
L_PTL_S2_3|_TX|P1 _PTL_S2_3|_TX|2 0  5.254e-13
L_PTL_S2_3|_TX|P2 _PTL_S2_3|_TX|5 0  5.141e-13
R_PTL_S2_3|_TX|B1 _PTL_S2_3|_TX|1 _PTL_S2_3|_TX|101  2.7439617672
R_PTL_S2_3|_TX|B2 _PTL_S2_3|_TX|4 _PTL_S2_3|_TX|104  2.7439617672
L_PTL_S2_3|_TX|RB1 _PTL_S2_3|_TX|101 0  1.550338398468e-12
L_PTL_S2_3|_TX|RB2 _PTL_S2_3|_TX|104 0  1.550338398468e-12
B_PTL_S2_3|_RX|1 _PTL_S2_3|_RX|1 _PTL_S2_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S2_3|_RX|2 _PTL_S2_3|_RX|4 _PTL_S2_3|_RX|5 JJMIT AREA=2.0
B_PTL_S2_3|_RX|3 _PTL_S2_3|_RX|7 _PTL_S2_3|_RX|8 JJMIT AREA=2.5
I_PTL_S2_3|_RX|B1 0 _PTL_S2_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S2_3|_RX|B1 _PTL_S2_3|_RX|1 _PTL_S2_3|_RX|3  2.777e-12
I_PTL_S2_3|_RX|B2 0 _PTL_S2_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S2_3|_RX|B2 _PTL_S2_3|_RX|4 _PTL_S2_3|_RX|6  2.685e-12
I_PTL_S2_3|_RX|B3 0 _PTL_S2_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S2_3|_RX|B3 _PTL_S2_3|_RX|7 _PTL_S2_3|_RX|9  2.764e-12
L_PTL_S2_3|_RX|1 _PTL_S2_3|A_PTL _PTL_S2_3|_RX|1  1.346e-12
L_PTL_S2_3|_RX|2 _PTL_S2_3|_RX|1 _PTL_S2_3|_RX|4  6.348e-12
L_PTL_S2_3|_RX|3 _PTL_S2_3|_RX|4 _PTL_S2_3|_RX|7  5.197e-12
L_PTL_S2_3|_RX|4 _PTL_S2_3|_RX|7 S2_3  2.058e-12
L_PTL_S2_3|_RX|P1 _PTL_S2_3|_RX|2 0  4.795e-13
L_PTL_S2_3|_RX|P2 _PTL_S2_3|_RX|5 0  5.431e-13
L_PTL_S2_3|_RX|P3 _PTL_S2_3|_RX|8 0  5.339e-13
R_PTL_S2_3|_RX|B1 _PTL_S2_3|_RX|1 _PTL_S2_3|_RX|101  4.225701121488
R_PTL_S2_3|_RX|B2 _PTL_S2_3|_RX|4 _PTL_S2_3|_RX|104  3.429952209
R_PTL_S2_3|_RX|B3 _PTL_S2_3|_RX|7 _PTL_S2_3|_RX|107  2.7439617672
L_PTL_S2_3|_RX|RB1 _PTL_S2_3|_RX|101 0  2.38752113364072e-12
L_PTL_S2_3|_RX|RB2 _PTL_S2_3|_RX|104 0  1.937922998085e-12
L_PTL_S2_3|_RX|RB3 _PTL_S2_3|_RX|107 0  1.550338398468e-12
B_PTL_S3_3|_TX|1 _PTL_S3_3|_TX|1 _PTL_S3_3|_TX|2 JJMIT AREA=2.5
B_PTL_S3_3|_TX|2 _PTL_S3_3|_TX|4 _PTL_S3_3|_TX|5 JJMIT AREA=2.5
I_PTL_S3_3|_TX|B1 0 _PTL_S3_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S3_3|_TX|B2 0 _PTL_S3_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S3_3|_TX|B1 _PTL_S3_3|_TX|1 _PTL_S3_3|_TX|3  1.684e-12
L_PTL_S3_3|_TX|B2 _PTL_S3_3|_TX|4 _PTL_S3_3|_TX|6  3.596e-12
L_PTL_S3_3|_TX|1 S3_3_TX _PTL_S3_3|_TX|1  2.063e-12
L_PTL_S3_3|_TX|2 _PTL_S3_3|_TX|1 _PTL_S3_3|_TX|4  4.123e-12
L_PTL_S3_3|_TX|3 _PTL_S3_3|_TX|4 _PTL_S3_3|_TX|7  2.193e-12
R_PTL_S3_3|_TX|D _PTL_S3_3|_TX|7 _PTL_S3_3|A_PTL  1.36
L_PTL_S3_3|_TX|P1 _PTL_S3_3|_TX|2 0  5.254e-13
L_PTL_S3_3|_TX|P2 _PTL_S3_3|_TX|5 0  5.141e-13
R_PTL_S3_3|_TX|B1 _PTL_S3_3|_TX|1 _PTL_S3_3|_TX|101  2.7439617672
R_PTL_S3_3|_TX|B2 _PTL_S3_3|_TX|4 _PTL_S3_3|_TX|104  2.7439617672
L_PTL_S3_3|_TX|RB1 _PTL_S3_3|_TX|101 0  1.550338398468e-12
L_PTL_S3_3|_TX|RB2 _PTL_S3_3|_TX|104 0  1.550338398468e-12
B_PTL_S3_3|_RX|1 _PTL_S3_3|_RX|1 _PTL_S3_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S3_3|_RX|2 _PTL_S3_3|_RX|4 _PTL_S3_3|_RX|5 JJMIT AREA=2.0
B_PTL_S3_3|_RX|3 _PTL_S3_3|_RX|7 _PTL_S3_3|_RX|8 JJMIT AREA=2.5
I_PTL_S3_3|_RX|B1 0 _PTL_S3_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S3_3|_RX|B1 _PTL_S3_3|_RX|1 _PTL_S3_3|_RX|3  2.777e-12
I_PTL_S3_3|_RX|B2 0 _PTL_S3_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S3_3|_RX|B2 _PTL_S3_3|_RX|4 _PTL_S3_3|_RX|6  2.685e-12
I_PTL_S3_3|_RX|B3 0 _PTL_S3_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S3_3|_RX|B3 _PTL_S3_3|_RX|7 _PTL_S3_3|_RX|9  2.764e-12
L_PTL_S3_3|_RX|1 _PTL_S3_3|A_PTL _PTL_S3_3|_RX|1  1.346e-12
L_PTL_S3_3|_RX|2 _PTL_S3_3|_RX|1 _PTL_S3_3|_RX|4  6.348e-12
L_PTL_S3_3|_RX|3 _PTL_S3_3|_RX|4 _PTL_S3_3|_RX|7  5.197e-12
L_PTL_S3_3|_RX|4 _PTL_S3_3|_RX|7 S3_3  2.058e-12
L_PTL_S3_3|_RX|P1 _PTL_S3_3|_RX|2 0  4.795e-13
L_PTL_S3_3|_RX|P2 _PTL_S3_3|_RX|5 0  5.431e-13
L_PTL_S3_3|_RX|P3 _PTL_S3_3|_RX|8 0  5.339e-13
R_PTL_S3_3|_RX|B1 _PTL_S3_3|_RX|1 _PTL_S3_3|_RX|101  4.225701121488
R_PTL_S3_3|_RX|B2 _PTL_S3_3|_RX|4 _PTL_S3_3|_RX|104  3.429952209
R_PTL_S3_3|_RX|B3 _PTL_S3_3|_RX|7 _PTL_S3_3|_RX|107  2.7439617672
L_PTL_S3_3|_RX|RB1 _PTL_S3_3|_RX|101 0  2.38752113364072e-12
L_PTL_S3_3|_RX|RB2 _PTL_S3_3|_RX|104 0  1.937922998085e-12
L_PTL_S3_3|_RX|RB3 _PTL_S3_3|_RX|107 0  1.550338398468e-12
B_PTL_S4_3|_TX|1 _PTL_S4_3|_TX|1 _PTL_S4_3|_TX|2 JJMIT AREA=2.5
B_PTL_S4_3|_TX|2 _PTL_S4_3|_TX|4 _PTL_S4_3|_TX|5 JJMIT AREA=2.5
I_PTL_S4_3|_TX|B1 0 _PTL_S4_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S4_3|_TX|B2 0 _PTL_S4_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S4_3|_TX|B1 _PTL_S4_3|_TX|1 _PTL_S4_3|_TX|3  1.684e-12
L_PTL_S4_3|_TX|B2 _PTL_S4_3|_TX|4 _PTL_S4_3|_TX|6  3.596e-12
L_PTL_S4_3|_TX|1 S4_3_TX _PTL_S4_3|_TX|1  2.063e-12
L_PTL_S4_3|_TX|2 _PTL_S4_3|_TX|1 _PTL_S4_3|_TX|4  4.123e-12
L_PTL_S4_3|_TX|3 _PTL_S4_3|_TX|4 _PTL_S4_3|_TX|7  2.193e-12
R_PTL_S4_3|_TX|D _PTL_S4_3|_TX|7 _PTL_S4_3|A_PTL  1.36
L_PTL_S4_3|_TX|P1 _PTL_S4_3|_TX|2 0  5.254e-13
L_PTL_S4_3|_TX|P2 _PTL_S4_3|_TX|5 0  5.141e-13
R_PTL_S4_3|_TX|B1 _PTL_S4_3|_TX|1 _PTL_S4_3|_TX|101  2.7439617672
R_PTL_S4_3|_TX|B2 _PTL_S4_3|_TX|4 _PTL_S4_3|_TX|104  2.7439617672
L_PTL_S4_3|_TX|RB1 _PTL_S4_3|_TX|101 0  1.550338398468e-12
L_PTL_S4_3|_TX|RB2 _PTL_S4_3|_TX|104 0  1.550338398468e-12
B_PTL_S4_3|_RX|1 _PTL_S4_3|_RX|1 _PTL_S4_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S4_3|_RX|2 _PTL_S4_3|_RX|4 _PTL_S4_3|_RX|5 JJMIT AREA=2.0
B_PTL_S4_3|_RX|3 _PTL_S4_3|_RX|7 _PTL_S4_3|_RX|8 JJMIT AREA=2.5
I_PTL_S4_3|_RX|B1 0 _PTL_S4_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S4_3|_RX|B1 _PTL_S4_3|_RX|1 _PTL_S4_3|_RX|3  2.777e-12
I_PTL_S4_3|_RX|B2 0 _PTL_S4_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S4_3|_RX|B2 _PTL_S4_3|_RX|4 _PTL_S4_3|_RX|6  2.685e-12
I_PTL_S4_3|_RX|B3 0 _PTL_S4_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S4_3|_RX|B3 _PTL_S4_3|_RX|7 _PTL_S4_3|_RX|9  2.764e-12
L_PTL_S4_3|_RX|1 _PTL_S4_3|A_PTL _PTL_S4_3|_RX|1  1.346e-12
L_PTL_S4_3|_RX|2 _PTL_S4_3|_RX|1 _PTL_S4_3|_RX|4  6.348e-12
L_PTL_S4_3|_RX|3 _PTL_S4_3|_RX|4 _PTL_S4_3|_RX|7  5.197e-12
L_PTL_S4_3|_RX|4 _PTL_S4_3|_RX|7 S4_3  2.058e-12
L_PTL_S4_3|_RX|P1 _PTL_S4_3|_RX|2 0  4.795e-13
L_PTL_S4_3|_RX|P2 _PTL_S4_3|_RX|5 0  5.431e-13
L_PTL_S4_3|_RX|P3 _PTL_S4_3|_RX|8 0  5.339e-13
R_PTL_S4_3|_RX|B1 _PTL_S4_3|_RX|1 _PTL_S4_3|_RX|101  4.225701121488
R_PTL_S4_3|_RX|B2 _PTL_S4_3|_RX|4 _PTL_S4_3|_RX|104  3.429952209
R_PTL_S4_3|_RX|B3 _PTL_S4_3|_RX|7 _PTL_S4_3|_RX|107  2.7439617672
L_PTL_S4_3|_RX|RB1 _PTL_S4_3|_RX|101 0  2.38752113364072e-12
L_PTL_S4_3|_RX|RB2 _PTL_S4_3|_RX|104 0  1.937922998085e-12
L_PTL_S4_3|_RX|RB3 _PTL_S4_3|_RX|107 0  1.550338398468e-12
B_PTL_G4_3|_TX|1 _PTL_G4_3|_TX|1 _PTL_G4_3|_TX|2 JJMIT AREA=2.5
B_PTL_G4_3|_TX|2 _PTL_G4_3|_TX|4 _PTL_G4_3|_TX|5 JJMIT AREA=2.5
I_PTL_G4_3|_TX|B1 0 _PTL_G4_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G4_3|_TX|B2 0 _PTL_G4_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G4_3|_TX|B1 _PTL_G4_3|_TX|1 _PTL_G4_3|_TX|3  1.684e-12
L_PTL_G4_3|_TX|B2 _PTL_G4_3|_TX|4 _PTL_G4_3|_TX|6  3.596e-12
L_PTL_G4_3|_TX|1 G4_3_TX _PTL_G4_3|_TX|1  2.063e-12
L_PTL_G4_3|_TX|2 _PTL_G4_3|_TX|1 _PTL_G4_3|_TX|4  4.123e-12
L_PTL_G4_3|_TX|3 _PTL_G4_3|_TX|4 _PTL_G4_3|_TX|7  2.193e-12
R_PTL_G4_3|_TX|D _PTL_G4_3|_TX|7 _PTL_G4_3|A_PTL  1.36
L_PTL_G4_3|_TX|P1 _PTL_G4_3|_TX|2 0  5.254e-13
L_PTL_G4_3|_TX|P2 _PTL_G4_3|_TX|5 0  5.141e-13
R_PTL_G4_3|_TX|B1 _PTL_G4_3|_TX|1 _PTL_G4_3|_TX|101  2.7439617672
R_PTL_G4_3|_TX|B2 _PTL_G4_3|_TX|4 _PTL_G4_3|_TX|104  2.7439617672
L_PTL_G4_3|_TX|RB1 _PTL_G4_3|_TX|101 0  1.550338398468e-12
L_PTL_G4_3|_TX|RB2 _PTL_G4_3|_TX|104 0  1.550338398468e-12
B_PTL_G4_3|_RX|1 _PTL_G4_3|_RX|1 _PTL_G4_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G4_3|_RX|2 _PTL_G4_3|_RX|4 _PTL_G4_3|_RX|5 JJMIT AREA=2.0
B_PTL_G4_3|_RX|3 _PTL_G4_3|_RX|7 _PTL_G4_3|_RX|8 JJMIT AREA=2.5
I_PTL_G4_3|_RX|B1 0 _PTL_G4_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G4_3|_RX|B1 _PTL_G4_3|_RX|1 _PTL_G4_3|_RX|3  2.777e-12
I_PTL_G4_3|_RX|B2 0 _PTL_G4_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G4_3|_RX|B2 _PTL_G4_3|_RX|4 _PTL_G4_3|_RX|6  2.685e-12
I_PTL_G4_3|_RX|B3 0 _PTL_G4_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G4_3|_RX|B3 _PTL_G4_3|_RX|7 _PTL_G4_3|_RX|9  2.764e-12
L_PTL_G4_3|_RX|1 _PTL_G4_3|A_PTL _PTL_G4_3|_RX|1  1.346e-12
L_PTL_G4_3|_RX|2 _PTL_G4_3|_RX|1 _PTL_G4_3|_RX|4  6.348e-12
L_PTL_G4_3|_RX|3 _PTL_G4_3|_RX|4 _PTL_G4_3|_RX|7  5.197e-12
L_PTL_G4_3|_RX|4 _PTL_G4_3|_RX|7 G4_3_OUT  2.058e-12
L_PTL_G4_3|_RX|P1 _PTL_G4_3|_RX|2 0  4.795e-13
L_PTL_G4_3|_RX|P2 _PTL_G4_3|_RX|5 0  5.431e-13
L_PTL_G4_3|_RX|P3 _PTL_G4_3|_RX|8 0  5.339e-13
R_PTL_G4_3|_RX|B1 _PTL_G4_3|_RX|1 _PTL_G4_3|_RX|101  4.225701121488
R_PTL_G4_3|_RX|B2 _PTL_G4_3|_RX|4 _PTL_G4_3|_RX|104  3.429952209
R_PTL_G4_3|_RX|B3 _PTL_G4_3|_RX|7 _PTL_G4_3|_RX|107  2.7439617672
L_PTL_G4_3|_RX|RB1 _PTL_G4_3|_RX|101 0  2.38752113364072e-12
L_PTL_G4_3|_RX|RB2 _PTL_G4_3|_RX|104 0  1.937922998085e-12
L_PTL_G4_3|_RX|RB3 _PTL_G4_3|_RX|107 0  1.550338398468e-12
B_PTL_IP5_3|_TX|1 _PTL_IP5_3|_TX|1 _PTL_IP5_3|_TX|2 JJMIT AREA=2.5
B_PTL_IP5_3|_TX|2 _PTL_IP5_3|_TX|4 _PTL_IP5_3|_TX|5 JJMIT AREA=2.5
I_PTL_IP5_3|_TX|B1 0 _PTL_IP5_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP5_3|_TX|B2 0 _PTL_IP5_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_3|_TX|B1 _PTL_IP5_3|_TX|1 _PTL_IP5_3|_TX|3  1.684e-12
L_PTL_IP5_3|_TX|B2 _PTL_IP5_3|_TX|4 _PTL_IP5_3|_TX|6  3.596e-12
L_PTL_IP5_3|_TX|1 IP5_3_OUT_TX _PTL_IP5_3|_TX|1  2.063e-12
L_PTL_IP5_3|_TX|2 _PTL_IP5_3|_TX|1 _PTL_IP5_3|_TX|4  4.123e-12
L_PTL_IP5_3|_TX|3 _PTL_IP5_3|_TX|4 _PTL_IP5_3|_TX|7  2.193e-12
R_PTL_IP5_3|_TX|D _PTL_IP5_3|_TX|7 _PTL_IP5_3|A_PTL  1.36
L_PTL_IP5_3|_TX|P1 _PTL_IP5_3|_TX|2 0  5.254e-13
L_PTL_IP5_3|_TX|P2 _PTL_IP5_3|_TX|5 0  5.141e-13
R_PTL_IP5_3|_TX|B1 _PTL_IP5_3|_TX|1 _PTL_IP5_3|_TX|101  2.7439617672
R_PTL_IP5_3|_TX|B2 _PTL_IP5_3|_TX|4 _PTL_IP5_3|_TX|104  2.7439617672
L_PTL_IP5_3|_TX|RB1 _PTL_IP5_3|_TX|101 0  1.550338398468e-12
L_PTL_IP5_3|_TX|RB2 _PTL_IP5_3|_TX|104 0  1.550338398468e-12
B_PTL_IP5_3|_RX|1 _PTL_IP5_3|_RX|1 _PTL_IP5_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP5_3|_RX|2 _PTL_IP5_3|_RX|4 _PTL_IP5_3|_RX|5 JJMIT AREA=2.0
B_PTL_IP5_3|_RX|3 _PTL_IP5_3|_RX|7 _PTL_IP5_3|_RX|8 JJMIT AREA=2.5
I_PTL_IP5_3|_RX|B1 0 _PTL_IP5_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP5_3|_RX|B1 _PTL_IP5_3|_RX|1 _PTL_IP5_3|_RX|3  2.777e-12
I_PTL_IP5_3|_RX|B2 0 _PTL_IP5_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP5_3|_RX|B2 _PTL_IP5_3|_RX|4 _PTL_IP5_3|_RX|6  2.685e-12
I_PTL_IP5_3|_RX|B3 0 _PTL_IP5_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_3|_RX|B3 _PTL_IP5_3|_RX|7 _PTL_IP5_3|_RX|9  2.764e-12
L_PTL_IP5_3|_RX|1 _PTL_IP5_3|A_PTL _PTL_IP5_3|_RX|1  1.346e-12
L_PTL_IP5_3|_RX|2 _PTL_IP5_3|_RX|1 _PTL_IP5_3|_RX|4  6.348e-12
L_PTL_IP5_3|_RX|3 _PTL_IP5_3|_RX|4 _PTL_IP5_3|_RX|7  5.197e-12
L_PTL_IP5_3|_RX|4 _PTL_IP5_3|_RX|7 IP5_3_OUT  2.058e-12
L_PTL_IP5_3|_RX|P1 _PTL_IP5_3|_RX|2 0  4.795e-13
L_PTL_IP5_3|_RX|P2 _PTL_IP5_3|_RX|5 0  5.431e-13
L_PTL_IP5_3|_RX|P3 _PTL_IP5_3|_RX|8 0  5.339e-13
R_PTL_IP5_3|_RX|B1 _PTL_IP5_3|_RX|1 _PTL_IP5_3|_RX|101  4.225701121488
R_PTL_IP5_3|_RX|B2 _PTL_IP5_3|_RX|4 _PTL_IP5_3|_RX|104  3.429952209
R_PTL_IP5_3|_RX|B3 _PTL_IP5_3|_RX|7 _PTL_IP5_3|_RX|107  2.7439617672
L_PTL_IP5_3|_RX|RB1 _PTL_IP5_3|_RX|101 0  2.38752113364072e-12
L_PTL_IP5_3|_RX|RB2 _PTL_IP5_3|_RX|104 0  1.937922998085e-12
L_PTL_IP5_3|_RX|RB3 _PTL_IP5_3|_RX|107 0  1.550338398468e-12
B_PTL_P5_3|_TX|1 _PTL_P5_3|_TX|1 _PTL_P5_3|_TX|2 JJMIT AREA=2.5
B_PTL_P5_3|_TX|2 _PTL_P5_3|_TX|4 _PTL_P5_3|_TX|5 JJMIT AREA=2.5
I_PTL_P5_3|_TX|B1 0 _PTL_P5_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P5_3|_TX|B2 0 _PTL_P5_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P5_3|_TX|B1 _PTL_P5_3|_TX|1 _PTL_P5_3|_TX|3  1.684e-12
L_PTL_P5_3|_TX|B2 _PTL_P5_3|_TX|4 _PTL_P5_3|_TX|6  3.596e-12
L_PTL_P5_3|_TX|1 P5_3_TX _PTL_P5_3|_TX|1  2.063e-12
L_PTL_P5_3|_TX|2 _PTL_P5_3|_TX|1 _PTL_P5_3|_TX|4  4.123e-12
L_PTL_P5_3|_TX|3 _PTL_P5_3|_TX|4 _PTL_P5_3|_TX|7  2.193e-12
R_PTL_P5_3|_TX|D _PTL_P5_3|_TX|7 _PTL_P5_3|A_PTL  1.36
L_PTL_P5_3|_TX|P1 _PTL_P5_3|_TX|2 0  5.254e-13
L_PTL_P5_3|_TX|P2 _PTL_P5_3|_TX|5 0  5.141e-13
R_PTL_P5_3|_TX|B1 _PTL_P5_3|_TX|1 _PTL_P5_3|_TX|101  2.7439617672
R_PTL_P5_3|_TX|B2 _PTL_P5_3|_TX|4 _PTL_P5_3|_TX|104  2.7439617672
L_PTL_P5_3|_TX|RB1 _PTL_P5_3|_TX|101 0  1.550338398468e-12
L_PTL_P5_3|_TX|RB2 _PTL_P5_3|_TX|104 0  1.550338398468e-12
B_PTL_P5_3|_RX|1 _PTL_P5_3|_RX|1 _PTL_P5_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P5_3|_RX|2 _PTL_P5_3|_RX|4 _PTL_P5_3|_RX|5 JJMIT AREA=2.0
B_PTL_P5_3|_RX|3 _PTL_P5_3|_RX|7 _PTL_P5_3|_RX|8 JJMIT AREA=2.5
I_PTL_P5_3|_RX|B1 0 _PTL_P5_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P5_3|_RX|B1 _PTL_P5_3|_RX|1 _PTL_P5_3|_RX|3  2.777e-12
I_PTL_P5_3|_RX|B2 0 _PTL_P5_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P5_3|_RX|B2 _PTL_P5_3|_RX|4 _PTL_P5_3|_RX|6  2.685e-12
I_PTL_P5_3|_RX|B3 0 _PTL_P5_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P5_3|_RX|B3 _PTL_P5_3|_RX|7 _PTL_P5_3|_RX|9  2.764e-12
L_PTL_P5_3|_RX|1 _PTL_P5_3|A_PTL _PTL_P5_3|_RX|1  1.346e-12
L_PTL_P5_3|_RX|2 _PTL_P5_3|_RX|1 _PTL_P5_3|_RX|4  6.348e-12
L_PTL_P5_3|_RX|3 _PTL_P5_3|_RX|4 _PTL_P5_3|_RX|7  5.197e-12
L_PTL_P5_3|_RX|4 _PTL_P5_3|_RX|7 P5_3_TO6  2.058e-12
L_PTL_P5_3|_RX|P1 _PTL_P5_3|_RX|2 0  4.795e-13
L_PTL_P5_3|_RX|P2 _PTL_P5_3|_RX|5 0  5.431e-13
L_PTL_P5_3|_RX|P3 _PTL_P5_3|_RX|8 0  5.339e-13
R_PTL_P5_3|_RX|B1 _PTL_P5_3|_RX|1 _PTL_P5_3|_RX|101  4.225701121488
R_PTL_P5_3|_RX|B2 _PTL_P5_3|_RX|4 _PTL_P5_3|_RX|104  3.429952209
R_PTL_P5_3|_RX|B3 _PTL_P5_3|_RX|7 _PTL_P5_3|_RX|107  2.7439617672
L_PTL_P5_3|_RX|RB1 _PTL_P5_3|_RX|101 0  2.38752113364072e-12
L_PTL_P5_3|_RX|RB2 _PTL_P5_3|_RX|104 0  1.937922998085e-12
L_PTL_P5_3|_RX|RB3 _PTL_P5_3|_RX|107 0  1.550338398468e-12
B_PTL_G5_3|_TX|1 _PTL_G5_3|_TX|1 _PTL_G5_3|_TX|2 JJMIT AREA=2.5
B_PTL_G5_3|_TX|2 _PTL_G5_3|_TX|4 _PTL_G5_3|_TX|5 JJMIT AREA=2.5
I_PTL_G5_3|_TX|B1 0 _PTL_G5_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G5_3|_TX|B2 0 _PTL_G5_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G5_3|_TX|B1 _PTL_G5_3|_TX|1 _PTL_G5_3|_TX|3  1.684e-12
L_PTL_G5_3|_TX|B2 _PTL_G5_3|_TX|4 _PTL_G5_3|_TX|6  3.596e-12
L_PTL_G5_3|_TX|1 G5_3_TX _PTL_G5_3|_TX|1  2.063e-12
L_PTL_G5_3|_TX|2 _PTL_G5_3|_TX|1 _PTL_G5_3|_TX|4  4.123e-12
L_PTL_G5_3|_TX|3 _PTL_G5_3|_TX|4 _PTL_G5_3|_TX|7  2.193e-12
R_PTL_G5_3|_TX|D _PTL_G5_3|_TX|7 _PTL_G5_3|A_PTL  1.36
L_PTL_G5_3|_TX|P1 _PTL_G5_3|_TX|2 0  5.254e-13
L_PTL_G5_3|_TX|P2 _PTL_G5_3|_TX|5 0  5.141e-13
R_PTL_G5_3|_TX|B1 _PTL_G5_3|_TX|1 _PTL_G5_3|_TX|101  2.7439617672
R_PTL_G5_3|_TX|B2 _PTL_G5_3|_TX|4 _PTL_G5_3|_TX|104  2.7439617672
L_PTL_G5_3|_TX|RB1 _PTL_G5_3|_TX|101 0  1.550338398468e-12
L_PTL_G5_3|_TX|RB2 _PTL_G5_3|_TX|104 0  1.550338398468e-12
B_PTL_G5_3|_RX|1 _PTL_G5_3|_RX|1 _PTL_G5_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G5_3|_RX|2 _PTL_G5_3|_RX|4 _PTL_G5_3|_RX|5 JJMIT AREA=2.0
B_PTL_G5_3|_RX|3 _PTL_G5_3|_RX|7 _PTL_G5_3|_RX|8 JJMIT AREA=2.5
I_PTL_G5_3|_RX|B1 0 _PTL_G5_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G5_3|_RX|B1 _PTL_G5_3|_RX|1 _PTL_G5_3|_RX|3  2.777e-12
I_PTL_G5_3|_RX|B2 0 _PTL_G5_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G5_3|_RX|B2 _PTL_G5_3|_RX|4 _PTL_G5_3|_RX|6  2.685e-12
I_PTL_G5_3|_RX|B3 0 _PTL_G5_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G5_3|_RX|B3 _PTL_G5_3|_RX|7 _PTL_G5_3|_RX|9  2.764e-12
L_PTL_G5_3|_RX|1 _PTL_G5_3|A_PTL _PTL_G5_3|_RX|1  1.346e-12
L_PTL_G5_3|_RX|2 _PTL_G5_3|_RX|1 _PTL_G5_3|_RX|4  6.348e-12
L_PTL_G5_3|_RX|3 _PTL_G5_3|_RX|4 _PTL_G5_3|_RX|7  5.197e-12
L_PTL_G5_3|_RX|4 _PTL_G5_3|_RX|7 _PTL_G5_3|D  2.058e-12
L_PTL_G5_3|_RX|P1 _PTL_G5_3|_RX|2 0  4.795e-13
L_PTL_G5_3|_RX|P2 _PTL_G5_3|_RX|5 0  5.431e-13
L_PTL_G5_3|_RX|P3 _PTL_G5_3|_RX|8 0  5.339e-13
R_PTL_G5_3|_RX|B1 _PTL_G5_3|_RX|1 _PTL_G5_3|_RX|101  4.225701121488
R_PTL_G5_3|_RX|B2 _PTL_G5_3|_RX|4 _PTL_G5_3|_RX|104  3.429952209
R_PTL_G5_3|_RX|B3 _PTL_G5_3|_RX|7 _PTL_G5_3|_RX|107  2.7439617672
L_PTL_G5_3|_RX|RB1 _PTL_G5_3|_RX|101 0  2.38752113364072e-12
L_PTL_G5_3|_RX|RB2 _PTL_G5_3|_RX|104 0  1.937922998085e-12
L_PTL_G5_3|_RX|RB3 _PTL_G5_3|_RX|107 0  1.550338398468e-12
L_PTL_G5_3|_SPL|1 _PTL_G5_3|D _PTL_G5_3|_SPL|D1  2e-12
L_PTL_G5_3|_SPL|2 _PTL_G5_3|_SPL|D1 _PTL_G5_3|_SPL|D2  4.135667696e-12
L_PTL_G5_3|_SPL|3 _PTL_G5_3|_SPL|D2 _PTL_G5_3|_SPL|JCT  9.84682784761905e-13
L_PTL_G5_3|_SPL|4 _PTL_G5_3|_SPL|JCT _PTL_G5_3|_SPL|QA1  9.84682784761905e-13
L_PTL_G5_3|_SPL|5 _PTL_G5_3|_SPL|QA1 G5_3_TO6  2e-12
L_PTL_G5_3|_SPL|6 _PTL_G5_3|_SPL|JCT _PTL_G5_3|_SPL|QB1  9.84682784761905e-13
L_PTL_G5_3|_SPL|7 _PTL_G5_3|_SPL|QB1 G5_3_OUT  2e-12
B_PTL_P6_3|_TX|1 _PTL_P6_3|_TX|1 _PTL_P6_3|_TX|2 JJMIT AREA=2.5
B_PTL_P6_3|_TX|2 _PTL_P6_3|_TX|4 _PTL_P6_3|_TX|5 JJMIT AREA=2.5
I_PTL_P6_3|_TX|B1 0 _PTL_P6_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_P6_3|_TX|B2 0 _PTL_P6_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_P6_3|_TX|B1 _PTL_P6_3|_TX|1 _PTL_P6_3|_TX|3  1.684e-12
L_PTL_P6_3|_TX|B2 _PTL_P6_3|_TX|4 _PTL_P6_3|_TX|6  3.596e-12
L_PTL_P6_3|_TX|1 P6_3_TX _PTL_P6_3|_TX|1  2.063e-12
L_PTL_P6_3|_TX|2 _PTL_P6_3|_TX|1 _PTL_P6_3|_TX|4  4.123e-12
L_PTL_P6_3|_TX|3 _PTL_P6_3|_TX|4 _PTL_P6_3|_TX|7  2.193e-12
R_PTL_P6_3|_TX|D _PTL_P6_3|_TX|7 _PTL_P6_3|A_PTL  1.36
L_PTL_P6_3|_TX|P1 _PTL_P6_3|_TX|2 0  5.254e-13
L_PTL_P6_3|_TX|P2 _PTL_P6_3|_TX|5 0  5.141e-13
R_PTL_P6_3|_TX|B1 _PTL_P6_3|_TX|1 _PTL_P6_3|_TX|101  2.7439617672
R_PTL_P6_3|_TX|B2 _PTL_P6_3|_TX|4 _PTL_P6_3|_TX|104  2.7439617672
L_PTL_P6_3|_TX|RB1 _PTL_P6_3|_TX|101 0  1.550338398468e-12
L_PTL_P6_3|_TX|RB2 _PTL_P6_3|_TX|104 0  1.550338398468e-12
B_PTL_P6_3|_RX|1 _PTL_P6_3|_RX|1 _PTL_P6_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_P6_3|_RX|2 _PTL_P6_3|_RX|4 _PTL_P6_3|_RX|5 JJMIT AREA=2.0
B_PTL_P6_3|_RX|3 _PTL_P6_3|_RX|7 _PTL_P6_3|_RX|8 JJMIT AREA=2.5
I_PTL_P6_3|_RX|B1 0 _PTL_P6_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_P6_3|_RX|B1 _PTL_P6_3|_RX|1 _PTL_P6_3|_RX|3  2.777e-12
I_PTL_P6_3|_RX|B2 0 _PTL_P6_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_P6_3|_RX|B2 _PTL_P6_3|_RX|4 _PTL_P6_3|_RX|6  2.685e-12
I_PTL_P6_3|_RX|B3 0 _PTL_P6_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_P6_3|_RX|B3 _PTL_P6_3|_RX|7 _PTL_P6_3|_RX|9  2.764e-12
L_PTL_P6_3|_RX|1 _PTL_P6_3|A_PTL _PTL_P6_3|_RX|1  1.346e-12
L_PTL_P6_3|_RX|2 _PTL_P6_3|_RX|1 _PTL_P6_3|_RX|4  6.348e-12
L_PTL_P6_3|_RX|3 _PTL_P6_3|_RX|4 _PTL_P6_3|_RX|7  5.197e-12
L_PTL_P6_3|_RX|4 _PTL_P6_3|_RX|7 _PTL_P6_3|D  2.058e-12
L_PTL_P6_3|_RX|P1 _PTL_P6_3|_RX|2 0  4.795e-13
L_PTL_P6_3|_RX|P2 _PTL_P6_3|_RX|5 0  5.431e-13
L_PTL_P6_3|_RX|P3 _PTL_P6_3|_RX|8 0  5.339e-13
R_PTL_P6_3|_RX|B1 _PTL_P6_3|_RX|1 _PTL_P6_3|_RX|101  4.225701121488
R_PTL_P6_3|_RX|B2 _PTL_P6_3|_RX|4 _PTL_P6_3|_RX|104  3.429952209
R_PTL_P6_3|_RX|B3 _PTL_P6_3|_RX|7 _PTL_P6_3|_RX|107  2.7439617672
L_PTL_P6_3|_RX|RB1 _PTL_P6_3|_RX|101 0  2.38752113364072e-12
L_PTL_P6_3|_RX|RB2 _PTL_P6_3|_RX|104 0  1.937922998085e-12
L_PTL_P6_3|_RX|RB3 _PTL_P6_3|_RX|107 0  1.550338398468e-12
L_PTL_P6_3|_SPL|1 _PTL_P6_3|D _PTL_P6_3|_SPL|D1  2e-12
L_PTL_P6_3|_SPL|2 _PTL_P6_3|_SPL|D1 _PTL_P6_3|_SPL|D2  4.135667696e-12
L_PTL_P6_3|_SPL|3 _PTL_P6_3|_SPL|D2 _PTL_P6_3|_SPL|JCT  9.84682784761905e-13
L_PTL_P6_3|_SPL|4 _PTL_P6_3|_SPL|JCT _PTL_P6_3|_SPL|QA1  9.84682784761905e-13
L_PTL_P6_3|_SPL|5 _PTL_P6_3|_SPL|QA1 P6_3_TO6  2e-12
L_PTL_P6_3|_SPL|6 _PTL_P6_3|_SPL|JCT _PTL_P6_3|_SPL|QB1  9.84682784761905e-13
L_PTL_P6_3|_SPL|7 _PTL_P6_3|_SPL|QB1 P6_3_OUT  2e-12
B_PTL_G6_3|_TX|1 _PTL_G6_3|_TX|1 _PTL_G6_3|_TX|2 JJMIT AREA=2.5
B_PTL_G6_3|_TX|2 _PTL_G6_3|_TX|4 _PTL_G6_3|_TX|5 JJMIT AREA=2.5
I_PTL_G6_3|_TX|B1 0 _PTL_G6_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G6_3|_TX|B2 0 _PTL_G6_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G6_3|_TX|B1 _PTL_G6_3|_TX|1 _PTL_G6_3|_TX|3  1.684e-12
L_PTL_G6_3|_TX|B2 _PTL_G6_3|_TX|4 _PTL_G6_3|_TX|6  3.596e-12
L_PTL_G6_3|_TX|1 G6_3_TX _PTL_G6_3|_TX|1  2.063e-12
L_PTL_G6_3|_TX|2 _PTL_G6_3|_TX|1 _PTL_G6_3|_TX|4  4.123e-12
L_PTL_G6_3|_TX|3 _PTL_G6_3|_TX|4 _PTL_G6_3|_TX|7  2.193e-12
R_PTL_G6_3|_TX|D _PTL_G6_3|_TX|7 _PTL_G6_3|A_PTL  1.36
L_PTL_G6_3|_TX|P1 _PTL_G6_3|_TX|2 0  5.254e-13
L_PTL_G6_3|_TX|P2 _PTL_G6_3|_TX|5 0  5.141e-13
R_PTL_G6_3|_TX|B1 _PTL_G6_3|_TX|1 _PTL_G6_3|_TX|101  2.7439617672
R_PTL_G6_3|_TX|B2 _PTL_G6_3|_TX|4 _PTL_G6_3|_TX|104  2.7439617672
L_PTL_G6_3|_TX|RB1 _PTL_G6_3|_TX|101 0  1.550338398468e-12
L_PTL_G6_3|_TX|RB2 _PTL_G6_3|_TX|104 0  1.550338398468e-12
B_PTL_G6_3|_RX|1 _PTL_G6_3|_RX|1 _PTL_G6_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G6_3|_RX|2 _PTL_G6_3|_RX|4 _PTL_G6_3|_RX|5 JJMIT AREA=2.0
B_PTL_G6_3|_RX|3 _PTL_G6_3|_RX|7 _PTL_G6_3|_RX|8 JJMIT AREA=2.5
I_PTL_G6_3|_RX|B1 0 _PTL_G6_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G6_3|_RX|B1 _PTL_G6_3|_RX|1 _PTL_G6_3|_RX|3  2.777e-12
I_PTL_G6_3|_RX|B2 0 _PTL_G6_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G6_3|_RX|B2 _PTL_G6_3|_RX|4 _PTL_G6_3|_RX|6  2.685e-12
I_PTL_G6_3|_RX|B3 0 _PTL_G6_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G6_3|_RX|B3 _PTL_G6_3|_RX|7 _PTL_G6_3|_RX|9  2.764e-12
L_PTL_G6_3|_RX|1 _PTL_G6_3|A_PTL _PTL_G6_3|_RX|1  1.346e-12
L_PTL_G6_3|_RX|2 _PTL_G6_3|_RX|1 _PTL_G6_3|_RX|4  6.348e-12
L_PTL_G6_3|_RX|3 _PTL_G6_3|_RX|4 _PTL_G6_3|_RX|7  5.197e-12
L_PTL_G6_3|_RX|4 _PTL_G6_3|_RX|7 G6_3_TO6  2.058e-12
L_PTL_G6_3|_RX|P1 _PTL_G6_3|_RX|2 0  4.795e-13
L_PTL_G6_3|_RX|P2 _PTL_G6_3|_RX|5 0  5.431e-13
L_PTL_G6_3|_RX|P3 _PTL_G6_3|_RX|8 0  5.339e-13
R_PTL_G6_3|_RX|B1 _PTL_G6_3|_RX|1 _PTL_G6_3|_RX|101  4.225701121488
R_PTL_G6_3|_RX|B2 _PTL_G6_3|_RX|4 _PTL_G6_3|_RX|104  3.429952209
R_PTL_G6_3|_RX|B3 _PTL_G6_3|_RX|7 _PTL_G6_3|_RX|107  2.7439617672
L_PTL_G6_3|_RX|RB1 _PTL_G6_3|_RX|101 0  2.38752113364072e-12
L_PTL_G6_3|_RX|RB2 _PTL_G6_3|_RX|104 0  1.937922998085e-12
L_PTL_G6_3|_RX|RB3 _PTL_G6_3|_RX|107 0  1.550338398468e-12
B_PTL_IP7_3|_TX|1 _PTL_IP7_3|_TX|1 _PTL_IP7_3|_TX|2 JJMIT AREA=2.5
B_PTL_IP7_3|_TX|2 _PTL_IP7_3|_TX|4 _PTL_IP7_3|_TX|5 JJMIT AREA=2.5
I_PTL_IP7_3|_TX|B1 0 _PTL_IP7_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP7_3|_TX|B2 0 _PTL_IP7_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_3|_TX|B1 _PTL_IP7_3|_TX|1 _PTL_IP7_3|_TX|3  1.684e-12
L_PTL_IP7_3|_TX|B2 _PTL_IP7_3|_TX|4 _PTL_IP7_3|_TX|6  3.596e-12
L_PTL_IP7_3|_TX|1 IP7_3_OUT_TX _PTL_IP7_3|_TX|1  2.063e-12
L_PTL_IP7_3|_TX|2 _PTL_IP7_3|_TX|1 _PTL_IP7_3|_TX|4  4.123e-12
L_PTL_IP7_3|_TX|3 _PTL_IP7_3|_TX|4 _PTL_IP7_3|_TX|7  2.193e-12
R_PTL_IP7_3|_TX|D _PTL_IP7_3|_TX|7 _PTL_IP7_3|A_PTL  1.36
L_PTL_IP7_3|_TX|P1 _PTL_IP7_3|_TX|2 0  5.254e-13
L_PTL_IP7_3|_TX|P2 _PTL_IP7_3|_TX|5 0  5.141e-13
R_PTL_IP7_3|_TX|B1 _PTL_IP7_3|_TX|1 _PTL_IP7_3|_TX|101  2.7439617672
R_PTL_IP7_3|_TX|B2 _PTL_IP7_3|_TX|4 _PTL_IP7_3|_TX|104  2.7439617672
L_PTL_IP7_3|_TX|RB1 _PTL_IP7_3|_TX|101 0  1.550338398468e-12
L_PTL_IP7_3|_TX|RB2 _PTL_IP7_3|_TX|104 0  1.550338398468e-12
B_PTL_IP7_3|_RX|1 _PTL_IP7_3|_RX|1 _PTL_IP7_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP7_3|_RX|2 _PTL_IP7_3|_RX|4 _PTL_IP7_3|_RX|5 JJMIT AREA=2.0
B_PTL_IP7_3|_RX|3 _PTL_IP7_3|_RX|7 _PTL_IP7_3|_RX|8 JJMIT AREA=2.5
I_PTL_IP7_3|_RX|B1 0 _PTL_IP7_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP7_3|_RX|B1 _PTL_IP7_3|_RX|1 _PTL_IP7_3|_RX|3  2.777e-12
I_PTL_IP7_3|_RX|B2 0 _PTL_IP7_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP7_3|_RX|B2 _PTL_IP7_3|_RX|4 _PTL_IP7_3|_RX|6  2.685e-12
I_PTL_IP7_3|_RX|B3 0 _PTL_IP7_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_3|_RX|B3 _PTL_IP7_3|_RX|7 _PTL_IP7_3|_RX|9  2.764e-12
L_PTL_IP7_3|_RX|1 _PTL_IP7_3|A_PTL _PTL_IP7_3|_RX|1  1.346e-12
L_PTL_IP7_3|_RX|2 _PTL_IP7_3|_RX|1 _PTL_IP7_3|_RX|4  6.348e-12
L_PTL_IP7_3|_RX|3 _PTL_IP7_3|_RX|4 _PTL_IP7_3|_RX|7  5.197e-12
L_PTL_IP7_3|_RX|4 _PTL_IP7_3|_RX|7 IP7_3_OUT  2.058e-12
L_PTL_IP7_3|_RX|P1 _PTL_IP7_3|_RX|2 0  4.795e-13
L_PTL_IP7_3|_RX|P2 _PTL_IP7_3|_RX|5 0  5.431e-13
L_PTL_IP7_3|_RX|P3 _PTL_IP7_3|_RX|8 0  5.339e-13
R_PTL_IP7_3|_RX|B1 _PTL_IP7_3|_RX|1 _PTL_IP7_3|_RX|101  4.225701121488
R_PTL_IP7_3|_RX|B2 _PTL_IP7_3|_RX|4 _PTL_IP7_3|_RX|104  3.429952209
R_PTL_IP7_3|_RX|B3 _PTL_IP7_3|_RX|7 _PTL_IP7_3|_RX|107  2.7439617672
L_PTL_IP7_3|_RX|RB1 _PTL_IP7_3|_RX|101 0  2.38752113364072e-12
L_PTL_IP7_3|_RX|RB2 _PTL_IP7_3|_RX|104 0  1.937922998085e-12
L_PTL_IP7_3|_RX|RB3 _PTL_IP7_3|_RX|107 0  1.550338398468e-12
B_PTL_S8_3|_TX|1 _PTL_S8_3|_TX|1 _PTL_S8_3|_TX|2 JJMIT AREA=2.5
B_PTL_S8_3|_TX|2 _PTL_S8_3|_TX|4 _PTL_S8_3|_TX|5 JJMIT AREA=2.5
I_PTL_S8_3|_TX|B1 0 _PTL_S8_3|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S8_3|_TX|B2 0 _PTL_S8_3|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S8_3|_TX|B1 _PTL_S8_3|_TX|1 _PTL_S8_3|_TX|3  1.684e-12
L_PTL_S8_3|_TX|B2 _PTL_S8_3|_TX|4 _PTL_S8_3|_TX|6  3.596e-12
L_PTL_S8_3|_TX|1 S8_3_TX _PTL_S8_3|_TX|1  2.063e-12
L_PTL_S8_3|_TX|2 _PTL_S8_3|_TX|1 _PTL_S8_3|_TX|4  4.123e-12
L_PTL_S8_3|_TX|3 _PTL_S8_3|_TX|4 _PTL_S8_3|_TX|7  2.193e-12
R_PTL_S8_3|_TX|D _PTL_S8_3|_TX|7 _PTL_S8_3|A_PTL  1.36
L_PTL_S8_3|_TX|P1 _PTL_S8_3|_TX|2 0  5.254e-13
L_PTL_S8_3|_TX|P2 _PTL_S8_3|_TX|5 0  5.141e-13
R_PTL_S8_3|_TX|B1 _PTL_S8_3|_TX|1 _PTL_S8_3|_TX|101  2.7439617672
R_PTL_S8_3|_TX|B2 _PTL_S8_3|_TX|4 _PTL_S8_3|_TX|104  2.7439617672
L_PTL_S8_3|_TX|RB1 _PTL_S8_3|_TX|101 0  1.550338398468e-12
L_PTL_S8_3|_TX|RB2 _PTL_S8_3|_TX|104 0  1.550338398468e-12
B_PTL_S8_3|_RX|1 _PTL_S8_3|_RX|1 _PTL_S8_3|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S8_3|_RX|2 _PTL_S8_3|_RX|4 _PTL_S8_3|_RX|5 JJMIT AREA=2.0
B_PTL_S8_3|_RX|3 _PTL_S8_3|_RX|7 _PTL_S8_3|_RX|8 JJMIT AREA=2.5
I_PTL_S8_3|_RX|B1 0 _PTL_S8_3|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S8_3|_RX|B1 _PTL_S8_3|_RX|1 _PTL_S8_3|_RX|3  2.777e-12
I_PTL_S8_3|_RX|B2 0 _PTL_S8_3|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S8_3|_RX|B2 _PTL_S8_3|_RX|4 _PTL_S8_3|_RX|6  2.685e-12
I_PTL_S8_3|_RX|B3 0 _PTL_S8_3|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S8_3|_RX|B3 _PTL_S8_3|_RX|7 _PTL_S8_3|_RX|9  2.764e-12
L_PTL_S8_3|_RX|1 _PTL_S8_3|A_PTL _PTL_S8_3|_RX|1  1.346e-12
L_PTL_S8_3|_RX|2 _PTL_S8_3|_RX|1 _PTL_S8_3|_RX|4  6.348e-12
L_PTL_S8_3|_RX|3 _PTL_S8_3|_RX|4 _PTL_S8_3|_RX|7  5.197e-12
L_PTL_S8_3|_RX|4 _PTL_S8_3|_RX|7 S8_3  2.058e-12
L_PTL_S8_3|_RX|P1 _PTL_S8_3|_RX|2 0  4.795e-13
L_PTL_S8_3|_RX|P2 _PTL_S8_3|_RX|5 0  5.431e-13
L_PTL_S8_3|_RX|P3 _PTL_S8_3|_RX|8 0  5.339e-13
R_PTL_S8_3|_RX|B1 _PTL_S8_3|_RX|1 _PTL_S8_3|_RX|101  4.225701121488
R_PTL_S8_3|_RX|B2 _PTL_S8_3|_RX|4 _PTL_S8_3|_RX|104  3.429952209
R_PTL_S8_3|_RX|B3 _PTL_S8_3|_RX|7 _PTL_S8_3|_RX|107  2.7439617672
L_PTL_S8_3|_RX|RB1 _PTL_S8_3|_RX|101 0  2.38752113364072e-12
L_PTL_S8_3|_RX|RB2 _PTL_S8_3|_RX|104 0  1.937922998085e-12
L_PTL_S8_3|_RX|RB3 _PTL_S8_3|_RX|107 0  1.550338398468e-12
L_S0_34|I_1|B _S0_34|A1 _S0_34|I_1|MID  2e-12
I_S0_34|I_1|B 0 _S0_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0_34|I_3|B _S0_34|A3 _S0_34|I_3|MID  2e-12
I_S0_34|I_3|B 0 _S0_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0_34|I_T|B _S0_34|T1 _S0_34|I_T|MID  2e-12
I_S0_34|I_T|B 0 _S0_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0_34|I_6|B _S0_34|Q1 _S0_34|I_6|MID  2e-12
I_S0_34|I_6|B 0 _S0_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0_34|1|1 _S0_34|A1 _S0_34|1|MID_SERIES JJMIT AREA=2.5
L_S0_34|1|P _S0_34|1|MID_SERIES 0  2e-13
R_S0_34|1|B _S0_34|A1 _S0_34|1|MID_SHUNT  2.7439617672
L_S0_34|1|RB _S0_34|1|MID_SHUNT 0  1.550338398468e-12
B_S0_34|23|1 _S0_34|A2 _S0_34|A3 JJMIT AREA=1.7857142857142858
R_S0_34|23|B _S0_34|A2 _S0_34|23|MID_SHUNT  3.84154647408
L_S0_34|23|RB _S0_34|23|MID_SHUNT _S0_34|A3  2.1704737578552e-12
B_S0_34|3|1 _S0_34|A3 _S0_34|3|MID_SERIES JJMIT AREA=2.5
L_S0_34|3|P _S0_34|3|MID_SERIES 0  2e-13
R_S0_34|3|B _S0_34|A3 _S0_34|3|MID_SHUNT  2.7439617672
L_S0_34|3|RB _S0_34|3|MID_SHUNT 0  1.550338398468e-12
B_S0_34|4|1 _S0_34|A4 _S0_34|4|MID_SERIES JJMIT AREA=2.5
L_S0_34|4|P _S0_34|4|MID_SERIES 0  2e-13
R_S0_34|4|B _S0_34|A4 _S0_34|4|MID_SHUNT  2.7439617672
L_S0_34|4|RB _S0_34|4|MID_SHUNT 0  1.550338398468e-12
B_S0_34|T|1 _S0_34|T1 _S0_34|T|MID_SERIES JJMIT AREA=2.5
L_S0_34|T|P _S0_34|T|MID_SERIES 0  2e-13
R_S0_34|T|B _S0_34|T1 _S0_34|T|MID_SHUNT  2.7439617672
L_S0_34|T|RB _S0_34|T|MID_SHUNT 0  1.550338398468e-12
B_S0_34|45|1 _S0_34|T2 _S0_34|A4 JJMIT AREA=1.7857142857142858
R_S0_34|45|B _S0_34|T2 _S0_34|45|MID_SHUNT  3.84154647408
L_S0_34|45|RB _S0_34|45|MID_SHUNT _S0_34|A4  2.1704737578552e-12
B_S0_34|6|1 _S0_34|Q1 _S0_34|6|MID_SERIES JJMIT AREA=2.5
L_S0_34|6|P _S0_34|6|MID_SERIES 0  2e-13
R_S0_34|6|B _S0_34|Q1 _S0_34|6|MID_SHUNT  2.7439617672
L_S0_34|6|RB _S0_34|6|MID_SHUNT 0  1.550338398468e-12
L_S1_34|I_1|B _S1_34|A1 _S1_34|I_1|MID  2e-12
I_S1_34|I_1|B 0 _S1_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S1_34|I_3|B _S1_34|A3 _S1_34|I_3|MID  2e-12
I_S1_34|I_3|B 0 _S1_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S1_34|I_T|B _S1_34|T1 _S1_34|I_T|MID  2e-12
I_S1_34|I_T|B 0 _S1_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S1_34|I_6|B _S1_34|Q1 _S1_34|I_6|MID  2e-12
I_S1_34|I_6|B 0 _S1_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S1_34|1|1 _S1_34|A1 _S1_34|1|MID_SERIES JJMIT AREA=2.5
L_S1_34|1|P _S1_34|1|MID_SERIES 0  2e-13
R_S1_34|1|B _S1_34|A1 _S1_34|1|MID_SHUNT  2.7439617672
L_S1_34|1|RB _S1_34|1|MID_SHUNT 0  1.550338398468e-12
B_S1_34|23|1 _S1_34|A2 _S1_34|A3 JJMIT AREA=1.7857142857142858
R_S1_34|23|B _S1_34|A2 _S1_34|23|MID_SHUNT  3.84154647408
L_S1_34|23|RB _S1_34|23|MID_SHUNT _S1_34|A3  2.1704737578552e-12
B_S1_34|3|1 _S1_34|A3 _S1_34|3|MID_SERIES JJMIT AREA=2.5
L_S1_34|3|P _S1_34|3|MID_SERIES 0  2e-13
R_S1_34|3|B _S1_34|A3 _S1_34|3|MID_SHUNT  2.7439617672
L_S1_34|3|RB _S1_34|3|MID_SHUNT 0  1.550338398468e-12
B_S1_34|4|1 _S1_34|A4 _S1_34|4|MID_SERIES JJMIT AREA=2.5
L_S1_34|4|P _S1_34|4|MID_SERIES 0  2e-13
R_S1_34|4|B _S1_34|A4 _S1_34|4|MID_SHUNT  2.7439617672
L_S1_34|4|RB _S1_34|4|MID_SHUNT 0  1.550338398468e-12
B_S1_34|T|1 _S1_34|T1 _S1_34|T|MID_SERIES JJMIT AREA=2.5
L_S1_34|T|P _S1_34|T|MID_SERIES 0  2e-13
R_S1_34|T|B _S1_34|T1 _S1_34|T|MID_SHUNT  2.7439617672
L_S1_34|T|RB _S1_34|T|MID_SHUNT 0  1.550338398468e-12
B_S1_34|45|1 _S1_34|T2 _S1_34|A4 JJMIT AREA=1.7857142857142858
R_S1_34|45|B _S1_34|T2 _S1_34|45|MID_SHUNT  3.84154647408
L_S1_34|45|RB _S1_34|45|MID_SHUNT _S1_34|A4  2.1704737578552e-12
B_S1_34|6|1 _S1_34|Q1 _S1_34|6|MID_SERIES JJMIT AREA=2.5
L_S1_34|6|P _S1_34|6|MID_SERIES 0  2e-13
R_S1_34|6|B _S1_34|Q1 _S1_34|6|MID_SHUNT  2.7439617672
L_S1_34|6|RB _S1_34|6|MID_SHUNT 0  1.550338398468e-12
L_S2_34|I_1|B _S2_34|A1 _S2_34|I_1|MID  2e-12
I_S2_34|I_1|B 0 _S2_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S2_34|I_3|B _S2_34|A3 _S2_34|I_3|MID  2e-12
I_S2_34|I_3|B 0 _S2_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S2_34|I_T|B _S2_34|T1 _S2_34|I_T|MID  2e-12
I_S2_34|I_T|B 0 _S2_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S2_34|I_6|B _S2_34|Q1 _S2_34|I_6|MID  2e-12
I_S2_34|I_6|B 0 _S2_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S2_34|1|1 _S2_34|A1 _S2_34|1|MID_SERIES JJMIT AREA=2.5
L_S2_34|1|P _S2_34|1|MID_SERIES 0  2e-13
R_S2_34|1|B _S2_34|A1 _S2_34|1|MID_SHUNT  2.7439617672
L_S2_34|1|RB _S2_34|1|MID_SHUNT 0  1.550338398468e-12
B_S2_34|23|1 _S2_34|A2 _S2_34|A3 JJMIT AREA=1.7857142857142858
R_S2_34|23|B _S2_34|A2 _S2_34|23|MID_SHUNT  3.84154647408
L_S2_34|23|RB _S2_34|23|MID_SHUNT _S2_34|A3  2.1704737578552e-12
B_S2_34|3|1 _S2_34|A3 _S2_34|3|MID_SERIES JJMIT AREA=2.5
L_S2_34|3|P _S2_34|3|MID_SERIES 0  2e-13
R_S2_34|3|B _S2_34|A3 _S2_34|3|MID_SHUNT  2.7439617672
L_S2_34|3|RB _S2_34|3|MID_SHUNT 0  1.550338398468e-12
B_S2_34|4|1 _S2_34|A4 _S2_34|4|MID_SERIES JJMIT AREA=2.5
L_S2_34|4|P _S2_34|4|MID_SERIES 0  2e-13
R_S2_34|4|B _S2_34|A4 _S2_34|4|MID_SHUNT  2.7439617672
L_S2_34|4|RB _S2_34|4|MID_SHUNT 0  1.550338398468e-12
B_S2_34|T|1 _S2_34|T1 _S2_34|T|MID_SERIES JJMIT AREA=2.5
L_S2_34|T|P _S2_34|T|MID_SERIES 0  2e-13
R_S2_34|T|B _S2_34|T1 _S2_34|T|MID_SHUNT  2.7439617672
L_S2_34|T|RB _S2_34|T|MID_SHUNT 0  1.550338398468e-12
B_S2_34|45|1 _S2_34|T2 _S2_34|A4 JJMIT AREA=1.7857142857142858
R_S2_34|45|B _S2_34|T2 _S2_34|45|MID_SHUNT  3.84154647408
L_S2_34|45|RB _S2_34|45|MID_SHUNT _S2_34|A4  2.1704737578552e-12
B_S2_34|6|1 _S2_34|Q1 _S2_34|6|MID_SERIES JJMIT AREA=2.5
L_S2_34|6|P _S2_34|6|MID_SERIES 0  2e-13
R_S2_34|6|B _S2_34|Q1 _S2_34|6|MID_SHUNT  2.7439617672
L_S2_34|6|RB _S2_34|6|MID_SHUNT 0  1.550338398468e-12
L_S3_34|I_1|B _S3_34|A1 _S3_34|I_1|MID  2e-12
I_S3_34|I_1|B 0 _S3_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S3_34|I_3|B _S3_34|A3 _S3_34|I_3|MID  2e-12
I_S3_34|I_3|B 0 _S3_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S3_34|I_T|B _S3_34|T1 _S3_34|I_T|MID  2e-12
I_S3_34|I_T|B 0 _S3_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S3_34|I_6|B _S3_34|Q1 _S3_34|I_6|MID  2e-12
I_S3_34|I_6|B 0 _S3_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S3_34|1|1 _S3_34|A1 _S3_34|1|MID_SERIES JJMIT AREA=2.5
L_S3_34|1|P _S3_34|1|MID_SERIES 0  2e-13
R_S3_34|1|B _S3_34|A1 _S3_34|1|MID_SHUNT  2.7439617672
L_S3_34|1|RB _S3_34|1|MID_SHUNT 0  1.550338398468e-12
B_S3_34|23|1 _S3_34|A2 _S3_34|A3 JJMIT AREA=1.7857142857142858
R_S3_34|23|B _S3_34|A2 _S3_34|23|MID_SHUNT  3.84154647408
L_S3_34|23|RB _S3_34|23|MID_SHUNT _S3_34|A3  2.1704737578552e-12
B_S3_34|3|1 _S3_34|A3 _S3_34|3|MID_SERIES JJMIT AREA=2.5
L_S3_34|3|P _S3_34|3|MID_SERIES 0  2e-13
R_S3_34|3|B _S3_34|A3 _S3_34|3|MID_SHUNT  2.7439617672
L_S3_34|3|RB _S3_34|3|MID_SHUNT 0  1.550338398468e-12
B_S3_34|4|1 _S3_34|A4 _S3_34|4|MID_SERIES JJMIT AREA=2.5
L_S3_34|4|P _S3_34|4|MID_SERIES 0  2e-13
R_S3_34|4|B _S3_34|A4 _S3_34|4|MID_SHUNT  2.7439617672
L_S3_34|4|RB _S3_34|4|MID_SHUNT 0  1.550338398468e-12
B_S3_34|T|1 _S3_34|T1 _S3_34|T|MID_SERIES JJMIT AREA=2.5
L_S3_34|T|P _S3_34|T|MID_SERIES 0  2e-13
R_S3_34|T|B _S3_34|T1 _S3_34|T|MID_SHUNT  2.7439617672
L_S3_34|T|RB _S3_34|T|MID_SHUNT 0  1.550338398468e-12
B_S3_34|45|1 _S3_34|T2 _S3_34|A4 JJMIT AREA=1.7857142857142858
R_S3_34|45|B _S3_34|T2 _S3_34|45|MID_SHUNT  3.84154647408
L_S3_34|45|RB _S3_34|45|MID_SHUNT _S3_34|A4  2.1704737578552e-12
B_S3_34|6|1 _S3_34|Q1 _S3_34|6|MID_SERIES JJMIT AREA=2.5
L_S3_34|6|P _S3_34|6|MID_SERIES 0  2e-13
R_S3_34|6|B _S3_34|Q1 _S3_34|6|MID_SHUNT  2.7439617672
L_S3_34|6|RB _S3_34|6|MID_SHUNT 0  1.550338398468e-12
L_S4_34|I_1|B _S4_34|A1 _S4_34|I_1|MID  2e-12
I_S4_34|I_1|B 0 _S4_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S4_34|I_3|B _S4_34|A3 _S4_34|I_3|MID  2e-12
I_S4_34|I_3|B 0 _S4_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S4_34|I_T|B _S4_34|T1 _S4_34|I_T|MID  2e-12
I_S4_34|I_T|B 0 _S4_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S4_34|I_6|B _S4_34|Q1 _S4_34|I_6|MID  2e-12
I_S4_34|I_6|B 0 _S4_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S4_34|1|1 _S4_34|A1 _S4_34|1|MID_SERIES JJMIT AREA=2.5
L_S4_34|1|P _S4_34|1|MID_SERIES 0  2e-13
R_S4_34|1|B _S4_34|A1 _S4_34|1|MID_SHUNT  2.7439617672
L_S4_34|1|RB _S4_34|1|MID_SHUNT 0  1.550338398468e-12
B_S4_34|23|1 _S4_34|A2 _S4_34|A3 JJMIT AREA=1.7857142857142858
R_S4_34|23|B _S4_34|A2 _S4_34|23|MID_SHUNT  3.84154647408
L_S4_34|23|RB _S4_34|23|MID_SHUNT _S4_34|A3  2.1704737578552e-12
B_S4_34|3|1 _S4_34|A3 _S4_34|3|MID_SERIES JJMIT AREA=2.5
L_S4_34|3|P _S4_34|3|MID_SERIES 0  2e-13
R_S4_34|3|B _S4_34|A3 _S4_34|3|MID_SHUNT  2.7439617672
L_S4_34|3|RB _S4_34|3|MID_SHUNT 0  1.550338398468e-12
B_S4_34|4|1 _S4_34|A4 _S4_34|4|MID_SERIES JJMIT AREA=2.5
L_S4_34|4|P _S4_34|4|MID_SERIES 0  2e-13
R_S4_34|4|B _S4_34|A4 _S4_34|4|MID_SHUNT  2.7439617672
L_S4_34|4|RB _S4_34|4|MID_SHUNT 0  1.550338398468e-12
B_S4_34|T|1 _S4_34|T1 _S4_34|T|MID_SERIES JJMIT AREA=2.5
L_S4_34|T|P _S4_34|T|MID_SERIES 0  2e-13
R_S4_34|T|B _S4_34|T1 _S4_34|T|MID_SHUNT  2.7439617672
L_S4_34|T|RB _S4_34|T|MID_SHUNT 0  1.550338398468e-12
B_S4_34|45|1 _S4_34|T2 _S4_34|A4 JJMIT AREA=1.7857142857142858
R_S4_34|45|B _S4_34|T2 _S4_34|45|MID_SHUNT  3.84154647408
L_S4_34|45|RB _S4_34|45|MID_SHUNT _S4_34|A4  2.1704737578552e-12
B_S4_34|6|1 _S4_34|Q1 _S4_34|6|MID_SERIES JJMIT AREA=2.5
L_S4_34|6|P _S4_34|6|MID_SERIES 0  2e-13
R_S4_34|6|B _S4_34|Q1 _S4_34|6|MID_SHUNT  2.7439617672
L_S4_34|6|RB _S4_34|6|MID_SHUNT 0  1.550338398468e-12
L_S5_34|I_A1|B _S5_34|A1 _S5_34|I_A1|MID  2e-12
I_S5_34|I_A1|B 0 _S5_34|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S5_34|I_A3|B _S5_34|A3 _S5_34|I_A3|MID  2e-12
I_S5_34|I_A3|B 0 _S5_34|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S5_34|I_B1|B _S5_34|B1 _S5_34|I_B1|MID  2e-12
I_S5_34|I_B1|B 0 _S5_34|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S5_34|I_B3|B _S5_34|B3 _S5_34|I_B3|MID  2e-12
I_S5_34|I_B3|B 0 _S5_34|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S5_34|I_Q1|B _S5_34|Q1 _S5_34|I_Q1|MID  2e-12
I_S5_34|I_Q1|B 0 _S5_34|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S5_34|A1|1 _S5_34|A1 _S5_34|A1|MID_SERIES JJMIT AREA=2.5
L_S5_34|A1|P _S5_34|A1|MID_SERIES 0  5e-13
R_S5_34|A1|B _S5_34|A1 _S5_34|A1|MID_SHUNT  2.7439617672
L_S5_34|A1|RB _S5_34|A1|MID_SHUNT 0  2.050338398468e-12
B_S5_34|A2|1 _S5_34|A2 _S5_34|A2|MID_SERIES JJMIT AREA=2.5
L_S5_34|A2|P _S5_34|A2|MID_SERIES 0  5e-13
R_S5_34|A2|B _S5_34|A2 _S5_34|A2|MID_SHUNT  2.7439617672
L_S5_34|A2|RB _S5_34|A2|MID_SHUNT 0  2.050338398468e-12
B_S5_34|A3|1 _S5_34|A2 _S5_34|A3|MID_SERIES JJMIT AREA=2.5
L_S5_34|A3|P _S5_34|A3|MID_SERIES _S5_34|A3  1.2e-12
R_S5_34|A3|B _S5_34|A2 _S5_34|A3|MID_SHUNT  2.7439617672
L_S5_34|A3|RB _S5_34|A3|MID_SHUNT _S5_34|A3  2.050338398468e-12
B_S5_34|B1|1 _S5_34|B1 _S5_34|B1|MID_SERIES JJMIT AREA=2.5
L_S5_34|B1|P _S5_34|B1|MID_SERIES 0  5e-13
R_S5_34|B1|B _S5_34|B1 _S5_34|B1|MID_SHUNT  2.7439617672
L_S5_34|B1|RB _S5_34|B1|MID_SHUNT 0  2.050338398468e-12
B_S5_34|B2|1 _S5_34|B2 _S5_34|B2|MID_SERIES JJMIT AREA=2.5
L_S5_34|B2|P _S5_34|B2|MID_SERIES 0  5e-13
R_S5_34|B2|B _S5_34|B2 _S5_34|B2|MID_SHUNT  2.7439617672
L_S5_34|B2|RB _S5_34|B2|MID_SHUNT 0  2.050338398468e-12
B_S5_34|B3|1 _S5_34|B2 _S5_34|B3|MID_SERIES JJMIT AREA=2.5
L_S5_34|B3|P _S5_34|B3|MID_SERIES _S5_34|B3  1.2e-12
R_S5_34|B3|B _S5_34|B2 _S5_34|B3|MID_SHUNT  2.7439617672
L_S5_34|B3|RB _S5_34|B3|MID_SHUNT _S5_34|B3  2.050338398468e-12
B_S5_34|T1|1 _S5_34|T1 _S5_34|T1|MID_SERIES JJMIT AREA=2.5
L_S5_34|T1|P _S5_34|T1|MID_SERIES 0  5e-13
R_S5_34|T1|B _S5_34|T1 _S5_34|T1|MID_SHUNT  2.7439617672
L_S5_34|T1|RB _S5_34|T1|MID_SHUNT 0  2.050338398468e-12
B_S5_34|T2|1 _S5_34|T2 _S5_34|ABTQ JJMIT AREA=2.0
R_S5_34|T2|B _S5_34|T2 _S5_34|T2|MID_SHUNT  3.429952209
L_S5_34|T2|RB _S5_34|T2|MID_SHUNT _S5_34|ABTQ  2.437922998085e-12
B_S5_34|AB|1 _S5_34|AB _S5_34|AB|MID_SERIES JJMIT AREA=1.5
L_S5_34|AB|P _S5_34|AB|MID_SERIES _S5_34|ABTQ  1.2e-12
R_S5_34|AB|B _S5_34|AB _S5_34|AB|MID_SHUNT  4.573269612
L_S5_34|AB|RB _S5_34|AB|MID_SHUNT _S5_34|ABTQ  3.08389733078e-12
B_S5_34|ABTQ|1 _S5_34|ABTQ _S5_34|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S5_34|ABTQ|P _S5_34|ABTQ|MID_SERIES 0  5e-13
R_S5_34|ABTQ|B _S5_34|ABTQ _S5_34|ABTQ|MID_SHUNT  3.6586156896
L_S5_34|ABTQ|RB _S5_34|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S5_34|Q1|1 _S5_34|Q1 _S5_34|Q1|MID_SERIES JJMIT AREA=2.5
L_S5_34|Q1|P _S5_34|Q1|MID_SERIES 0  5e-13
R_S5_34|Q1|B _S5_34|Q1 _S5_34|Q1|MID_SHUNT  2.7439617672
L_S5_34|Q1|RB _S5_34|Q1|MID_SHUNT 0  2.050338398468e-12
L_S6_34|I_A1|B _S6_34|A1 _S6_34|I_A1|MID  2e-12
I_S6_34|I_A1|B 0 _S6_34|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S6_34|I_A3|B _S6_34|A3 _S6_34|I_A3|MID  2e-12
I_S6_34|I_A3|B 0 _S6_34|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S6_34|I_B1|B _S6_34|B1 _S6_34|I_B1|MID  2e-12
I_S6_34|I_B1|B 0 _S6_34|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S6_34|I_B3|B _S6_34|B3 _S6_34|I_B3|MID  2e-12
I_S6_34|I_B3|B 0 _S6_34|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S6_34|I_Q1|B _S6_34|Q1 _S6_34|I_Q1|MID  2e-12
I_S6_34|I_Q1|B 0 _S6_34|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S6_34|A1|1 _S6_34|A1 _S6_34|A1|MID_SERIES JJMIT AREA=2.5
L_S6_34|A1|P _S6_34|A1|MID_SERIES 0  5e-13
R_S6_34|A1|B _S6_34|A1 _S6_34|A1|MID_SHUNT  2.7439617672
L_S6_34|A1|RB _S6_34|A1|MID_SHUNT 0  2.050338398468e-12
B_S6_34|A2|1 _S6_34|A2 _S6_34|A2|MID_SERIES JJMIT AREA=2.5
L_S6_34|A2|P _S6_34|A2|MID_SERIES 0  5e-13
R_S6_34|A2|B _S6_34|A2 _S6_34|A2|MID_SHUNT  2.7439617672
L_S6_34|A2|RB _S6_34|A2|MID_SHUNT 0  2.050338398468e-12
B_S6_34|A3|1 _S6_34|A2 _S6_34|A3|MID_SERIES JJMIT AREA=2.5
L_S6_34|A3|P _S6_34|A3|MID_SERIES _S6_34|A3  1.2e-12
R_S6_34|A3|B _S6_34|A2 _S6_34|A3|MID_SHUNT  2.7439617672
L_S6_34|A3|RB _S6_34|A3|MID_SHUNT _S6_34|A3  2.050338398468e-12
B_S6_34|B1|1 _S6_34|B1 _S6_34|B1|MID_SERIES JJMIT AREA=2.5
L_S6_34|B1|P _S6_34|B1|MID_SERIES 0  5e-13
R_S6_34|B1|B _S6_34|B1 _S6_34|B1|MID_SHUNT  2.7439617672
L_S6_34|B1|RB _S6_34|B1|MID_SHUNT 0  2.050338398468e-12
B_S6_34|B2|1 _S6_34|B2 _S6_34|B2|MID_SERIES JJMIT AREA=2.5
L_S6_34|B2|P _S6_34|B2|MID_SERIES 0  5e-13
R_S6_34|B2|B _S6_34|B2 _S6_34|B2|MID_SHUNT  2.7439617672
L_S6_34|B2|RB _S6_34|B2|MID_SHUNT 0  2.050338398468e-12
B_S6_34|B3|1 _S6_34|B2 _S6_34|B3|MID_SERIES JJMIT AREA=2.5
L_S6_34|B3|P _S6_34|B3|MID_SERIES _S6_34|B3  1.2e-12
R_S6_34|B3|B _S6_34|B2 _S6_34|B3|MID_SHUNT  2.7439617672
L_S6_34|B3|RB _S6_34|B3|MID_SHUNT _S6_34|B3  2.050338398468e-12
B_S6_34|T1|1 _S6_34|T1 _S6_34|T1|MID_SERIES JJMIT AREA=2.5
L_S6_34|T1|P _S6_34|T1|MID_SERIES 0  5e-13
R_S6_34|T1|B _S6_34|T1 _S6_34|T1|MID_SHUNT  2.7439617672
L_S6_34|T1|RB _S6_34|T1|MID_SHUNT 0  2.050338398468e-12
B_S6_34|T2|1 _S6_34|T2 _S6_34|ABTQ JJMIT AREA=2.0
R_S6_34|T2|B _S6_34|T2 _S6_34|T2|MID_SHUNT  3.429952209
L_S6_34|T2|RB _S6_34|T2|MID_SHUNT _S6_34|ABTQ  2.437922998085e-12
B_S6_34|AB|1 _S6_34|AB _S6_34|AB|MID_SERIES JJMIT AREA=1.5
L_S6_34|AB|P _S6_34|AB|MID_SERIES _S6_34|ABTQ  1.2e-12
R_S6_34|AB|B _S6_34|AB _S6_34|AB|MID_SHUNT  4.573269612
L_S6_34|AB|RB _S6_34|AB|MID_SHUNT _S6_34|ABTQ  3.08389733078e-12
B_S6_34|ABTQ|1 _S6_34|ABTQ _S6_34|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S6_34|ABTQ|P _S6_34|ABTQ|MID_SERIES 0  5e-13
R_S6_34|ABTQ|B _S6_34|ABTQ _S6_34|ABTQ|MID_SHUNT  3.6586156896
L_S6_34|ABTQ|RB _S6_34|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S6_34|Q1|1 _S6_34|Q1 _S6_34|Q1|MID_SERIES JJMIT AREA=2.5
L_S6_34|Q1|P _S6_34|Q1|MID_SERIES 0  5e-13
R_S6_34|Q1|B _S6_34|Q1 _S6_34|Q1|MID_SHUNT  2.7439617672
L_S6_34|Q1|RB _S6_34|Q1|MID_SHUNT 0  2.050338398468e-12
L_PG6_34|_SPL_G1|1 G6_3_TO6 _PG6_34|_SPL_G1|D1  2e-12
L_PG6_34|_SPL_G1|2 _PG6_34|_SPL_G1|D1 _PG6_34|_SPL_G1|D2  4.135667696e-12
L_PG6_34|_SPL_G1|3 _PG6_34|_SPL_G1|D2 _PG6_34|_SPL_G1|JCT  9.84682784761905e-13
L_PG6_34|_SPL_G1|4 _PG6_34|_SPL_G1|JCT _PG6_34|_SPL_G1|QA1  9.84682784761905e-13
L_PG6_34|_SPL_G1|5 _PG6_34|_SPL_G1|QA1 _PG6_34|G1_COPY_1  2e-12
L_PG6_34|_SPL_G1|6 _PG6_34|_SPL_G1|JCT _PG6_34|_SPL_G1|QB1  9.84682784761905e-13
L_PG6_34|_SPL_G1|7 _PG6_34|_SPL_G1|QB1 _PG6_34|G1_COPY_2  2e-12
L_PG6_34|_SPL_P1|1 P6_3_TO6 _PG6_34|_SPL_P1|D1  2e-12
L_PG6_34|_SPL_P1|2 _PG6_34|_SPL_P1|D1 _PG6_34|_SPL_P1|D2  4.135667696e-12
L_PG6_34|_SPL_P1|3 _PG6_34|_SPL_P1|D2 _PG6_34|_SPL_P1|JCT  9.84682784761905e-13
L_PG6_34|_SPL_P1|4 _PG6_34|_SPL_P1|JCT _PG6_34|_SPL_P1|QA1  9.84682784761905e-13
L_PG6_34|_SPL_P1|5 _PG6_34|_SPL_P1|QA1 _PG6_34|P1_COPY_1  2e-12
L_PG6_34|_SPL_P1|6 _PG6_34|_SPL_P1|JCT _PG6_34|_SPL_P1|QB1  9.84682784761905e-13
L_PG6_34|_SPL_P1|7 _PG6_34|_SPL_P1|QB1 _PG6_34|P1_COPY_2  2e-12
L_PG6_34|_PG|A1 _PG6_34|P1_COPY_1 _PG6_34|_PG|A1  2.067833848e-12
L_PG6_34|_PG|A2 _PG6_34|_PG|A1 _PG6_34|_PG|A2  4.135667696e-12
L_PG6_34|_PG|A3 _PG6_34|_PG|A3 _PG6_34|_PG|Q3  1.2e-12
L_PG6_34|_PG|B1 _PG6_34|G1_COPY_1 _PG6_34|_PG|B1  2.067833848e-12
L_PG6_34|_PG|B2 _PG6_34|_PG|B1 _PG6_34|_PG|B2  4.135667696e-12
L_PG6_34|_PG|B3 _PG6_34|_PG|B3 _PG6_34|_PG|Q3  1.2e-12
L_PG6_34|_PG|Q3 _PG6_34|_PG|Q3 _PG6_34|_PG|Q2  4.135667696e-12
L_PG6_34|_PG|Q2 _PG6_34|_PG|Q2 _PG6_34|_PG|Q1  4.135667696e-12
L_PG6_34|_PG|Q1 _PG6_34|_PG|Q1 _PG6_34|PG  2.067833848e-12
L_PG6_34|_GG|A1 G5_3_TO6 _PG6_34|_GG|A1  2.067833848e-12
L_PG6_34|_GG|A2 _PG6_34|_GG|A1 _PG6_34|_GG|A2  4.135667696e-12
L_PG6_34|_GG|A3 _PG6_34|_GG|A3 _PG6_34|_GG|Q3  1.2e-12
L_PG6_34|_GG|B1 _PG6_34|G1_COPY_2 _PG6_34|_GG|B1  2.067833848e-12
L_PG6_34|_GG|B2 _PG6_34|_GG|B1 _PG6_34|_GG|B2  4.135667696e-12
L_PG6_34|_GG|B3 _PG6_34|_GG|B3 _PG6_34|_GG|Q3  1.2e-12
L_PG6_34|_GG|Q3 _PG6_34|_GG|Q3 _PG6_34|_GG|Q2  4.135667696e-12
L_PG6_34|_GG|Q2 _PG6_34|_GG|Q2 _PG6_34|_GG|Q1  4.135667696e-12
L_PG6_34|_GG|Q1 _PG6_34|_GG|Q1 _PG6_34|GG  2.067833848e-12
L_PG6_34|_DFF_P0|1 P5_3_TO6 _PG6_34|_DFF_P0|A1  2.067833848e-12
L_PG6_34|_DFF_P0|2 _PG6_34|_DFF_P0|A1 _PG6_34|_DFF_P0|A2  4.135667696e-12
L_PG6_34|_DFF_P0|3 _PG6_34|_DFF_P0|A3 _PG6_34|_DFF_P0|A4  8.271335392e-12
L_PG6_34|_DFF_P0|T T47 _PG6_34|_DFF_P0|T1  2.067833848e-12
L_PG6_34|_DFF_P0|4 _PG6_34|_DFF_P0|T1 _PG6_34|_DFF_P0|T2  4.135667696e-12
L_PG6_34|_DFF_P0|5 _PG6_34|_DFF_P0|A4 _PG6_34|_DFF_P0|Q1  4.135667696e-12
L_PG6_34|_DFF_P0|6 _PG6_34|_DFF_P0|Q1 _PG6_34|P0_SYNC  2.067833848e-12
L_PG6_34|_DFF_P1|1 _PG6_34|P1_COPY_2 _PG6_34|_DFF_P1|A1  2.067833848e-12
L_PG6_34|_DFF_P1|2 _PG6_34|_DFF_P1|A1 _PG6_34|_DFF_P1|A2  4.135667696e-12
L_PG6_34|_DFF_P1|3 _PG6_34|_DFF_P1|A3 _PG6_34|_DFF_P1|A4  8.271335392e-12
L_PG6_34|_DFF_P1|T T47 _PG6_34|_DFF_P1|T1  2.067833848e-12
L_PG6_34|_DFF_P1|4 _PG6_34|_DFF_P1|T1 _PG6_34|_DFF_P1|T2  4.135667696e-12
L_PG6_34|_DFF_P1|5 _PG6_34|_DFF_P1|A4 _PG6_34|_DFF_P1|Q1  4.135667696e-12
L_PG6_34|_DFF_P1|6 _PG6_34|_DFF_P1|Q1 _PG6_34|P1_SYNC  2.067833848e-12
L_PG6_34|_DFF_PG|1 _PG6_34|PG _PG6_34|_DFF_PG|A1  2.067833848e-12
L_PG6_34|_DFF_PG|2 _PG6_34|_DFF_PG|A1 _PG6_34|_DFF_PG|A2  4.135667696e-12
L_PG6_34|_DFF_PG|3 _PG6_34|_DFF_PG|A3 _PG6_34|_DFF_PG|A4  8.271335392e-12
L_PG6_34|_DFF_PG|T T47 _PG6_34|_DFF_PG|T1  2.067833848e-12
L_PG6_34|_DFF_PG|4 _PG6_34|_DFF_PG|T1 _PG6_34|_DFF_PG|T2  4.135667696e-12
L_PG6_34|_DFF_PG|5 _PG6_34|_DFF_PG|A4 _PG6_34|_DFF_PG|Q1  4.135667696e-12
L_PG6_34|_DFF_PG|6 _PG6_34|_DFF_PG|Q1 _PG6_34|PG_SYNC  2.067833848e-12
L_PG6_34|_DFF_GG|1 _PG6_34|GG _PG6_34|_DFF_GG|A1  2.067833848e-12
L_PG6_34|_DFF_GG|2 _PG6_34|_DFF_GG|A1 _PG6_34|_DFF_GG|A2  4.135667696e-12
L_PG6_34|_DFF_GG|3 _PG6_34|_DFF_GG|A3 _PG6_34|_DFF_GG|A4  8.271335392e-12
L_PG6_34|_DFF_GG|T T47 _PG6_34|_DFF_GG|T1  2.067833848e-12
L_PG6_34|_DFF_GG|4 _PG6_34|_DFF_GG|T1 _PG6_34|_DFF_GG|T2  4.135667696e-12
L_PG6_34|_DFF_GG|5 _PG6_34|_DFF_GG|A4 _PG6_34|_DFF_GG|Q1  4.135667696e-12
L_PG6_34|_DFF_GG|6 _PG6_34|_DFF_GG|Q1 _PG6_34|GG_SYNC  2.067833848e-12
L_PG6_34|_AND_G|A1 _PG6_34|PG_SYNC _PG6_34|_AND_G|A1  2.067833848e-12
L_PG6_34|_AND_G|A2 _PG6_34|_AND_G|A1 _PG6_34|_AND_G|A2  4.135667696e-12
L_PG6_34|_AND_G|A3 _PG6_34|_AND_G|A3 _PG6_34|_AND_G|Q3  1.2e-12
L_PG6_34|_AND_G|B1 _PG6_34|GG_SYNC _PG6_34|_AND_G|B1  2.067833848e-12
L_PG6_34|_AND_G|B2 _PG6_34|_AND_G|B1 _PG6_34|_AND_G|B2  4.135667696e-12
L_PG6_34|_AND_G|B3 _PG6_34|_AND_G|B3 _PG6_34|_AND_G|Q3  1.2e-12
L_PG6_34|_AND_G|Q3 _PG6_34|_AND_G|Q3 _PG6_34|_AND_G|Q2  4.135667696e-12
L_PG6_34|_AND_G|Q2 _PG6_34|_AND_G|Q2 _PG6_34|_AND_G|Q1  4.135667696e-12
L_PG6_34|_AND_G|Q1 _PG6_34|_AND_G|Q1 G6_4_TX  2.067833848e-12
L_PG6_34|_AND_P|A1 _PG6_34|P0_SYNC _PG6_34|_AND_P|A1  2.067833848e-12
L_PG6_34|_AND_P|A2 _PG6_34|_AND_P|A1 _PG6_34|_AND_P|A2  4.135667696e-12
L_PG6_34|_AND_P|A3 _PG6_34|_AND_P|A3 _PG6_34|_AND_P|Q3  1.2e-12
L_PG6_34|_AND_P|B1 _PG6_34|P1_SYNC _PG6_34|_AND_P|B1  2.067833848e-12
L_PG6_34|_AND_P|B2 _PG6_34|_AND_P|B1 _PG6_34|_AND_P|B2  4.135667696e-12
L_PG6_34|_AND_P|B3 _PG6_34|_AND_P|B3 _PG6_34|_AND_P|Q3  1.2e-12
L_PG6_34|_AND_P|Q3 _PG6_34|_AND_P|Q3 _PG6_34|_AND_P|Q2  4.135667696e-12
L_PG6_34|_AND_P|Q2 _PG6_34|_AND_P|Q2 _PG6_34|_AND_P|Q1  4.135667696e-12
L_PG6_34|_AND_P|Q1 _PG6_34|_AND_P|Q1 P6_4_TX  2.067833848e-12
L_IP7_34|I_1|B _IP7_34|A1 _IP7_34|I_1|MID  2e-12
I_IP7_34|I_1|B 0 _IP7_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_IP7_34|I_3|B _IP7_34|A3 _IP7_34|I_3|MID  2e-12
I_IP7_34|I_3|B 0 _IP7_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_IP7_34|I_T|B _IP7_34|T1 _IP7_34|I_T|MID  2e-12
I_IP7_34|I_T|B 0 _IP7_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_IP7_34|I_6|B _IP7_34|Q1 _IP7_34|I_6|MID  2e-12
I_IP7_34|I_6|B 0 _IP7_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_IP7_34|1|1 _IP7_34|A1 _IP7_34|1|MID_SERIES JJMIT AREA=2.5
L_IP7_34|1|P _IP7_34|1|MID_SERIES 0  2e-13
R_IP7_34|1|B _IP7_34|A1 _IP7_34|1|MID_SHUNT  2.7439617672
L_IP7_34|1|RB _IP7_34|1|MID_SHUNT 0  1.550338398468e-12
B_IP7_34|23|1 _IP7_34|A2 _IP7_34|A3 JJMIT AREA=1.7857142857142858
R_IP7_34|23|B _IP7_34|A2 _IP7_34|23|MID_SHUNT  3.84154647408
L_IP7_34|23|RB _IP7_34|23|MID_SHUNT _IP7_34|A3  2.1704737578552e-12
B_IP7_34|3|1 _IP7_34|A3 _IP7_34|3|MID_SERIES JJMIT AREA=2.5
L_IP7_34|3|P _IP7_34|3|MID_SERIES 0  2e-13
R_IP7_34|3|B _IP7_34|A3 _IP7_34|3|MID_SHUNT  2.7439617672
L_IP7_34|3|RB _IP7_34|3|MID_SHUNT 0  1.550338398468e-12
B_IP7_34|4|1 _IP7_34|A4 _IP7_34|4|MID_SERIES JJMIT AREA=2.5
L_IP7_34|4|P _IP7_34|4|MID_SERIES 0  2e-13
R_IP7_34|4|B _IP7_34|A4 _IP7_34|4|MID_SHUNT  2.7439617672
L_IP7_34|4|RB _IP7_34|4|MID_SHUNT 0  1.550338398468e-12
B_IP7_34|T|1 _IP7_34|T1 _IP7_34|T|MID_SERIES JJMIT AREA=2.5
L_IP7_34|T|P _IP7_34|T|MID_SERIES 0  2e-13
R_IP7_34|T|B _IP7_34|T1 _IP7_34|T|MID_SHUNT  2.7439617672
L_IP7_34|T|RB _IP7_34|T|MID_SHUNT 0  1.550338398468e-12
B_IP7_34|45|1 _IP7_34|T2 _IP7_34|A4 JJMIT AREA=1.7857142857142858
R_IP7_34|45|B _IP7_34|T2 _IP7_34|45|MID_SHUNT  3.84154647408
L_IP7_34|45|RB _IP7_34|45|MID_SHUNT _IP7_34|A4  2.1704737578552e-12
B_IP7_34|6|1 _IP7_34|Q1 _IP7_34|6|MID_SERIES JJMIT AREA=2.5
L_IP7_34|6|P _IP7_34|6|MID_SERIES 0  2e-13
R_IP7_34|6|B _IP7_34|Q1 _IP7_34|6|MID_SHUNT  2.7439617672
L_IP7_34|6|RB _IP7_34|6|MID_SHUNT 0  1.550338398468e-12
L_S8_34|I_1|B _S8_34|A1 _S8_34|I_1|MID  2e-12
I_S8_34|I_1|B 0 _S8_34|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S8_34|I_3|B _S8_34|A3 _S8_34|I_3|MID  2e-12
I_S8_34|I_3|B 0 _S8_34|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S8_34|I_T|B _S8_34|T1 _S8_34|I_T|MID  2e-12
I_S8_34|I_T|B 0 _S8_34|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S8_34|I_6|B _S8_34|Q1 _S8_34|I_6|MID  2e-12
I_S8_34|I_6|B 0 _S8_34|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S8_34|1|1 _S8_34|A1 _S8_34|1|MID_SERIES JJMIT AREA=2.5
L_S8_34|1|P _S8_34|1|MID_SERIES 0  2e-13
R_S8_34|1|B _S8_34|A1 _S8_34|1|MID_SHUNT  2.7439617672
L_S8_34|1|RB _S8_34|1|MID_SHUNT 0  1.550338398468e-12
B_S8_34|23|1 _S8_34|A2 _S8_34|A3 JJMIT AREA=1.7857142857142858
R_S8_34|23|B _S8_34|A2 _S8_34|23|MID_SHUNT  3.84154647408
L_S8_34|23|RB _S8_34|23|MID_SHUNT _S8_34|A3  2.1704737578552e-12
B_S8_34|3|1 _S8_34|A3 _S8_34|3|MID_SERIES JJMIT AREA=2.5
L_S8_34|3|P _S8_34|3|MID_SERIES 0  2e-13
R_S8_34|3|B _S8_34|A3 _S8_34|3|MID_SHUNT  2.7439617672
L_S8_34|3|RB _S8_34|3|MID_SHUNT 0  1.550338398468e-12
B_S8_34|4|1 _S8_34|A4 _S8_34|4|MID_SERIES JJMIT AREA=2.5
L_S8_34|4|P _S8_34|4|MID_SERIES 0  2e-13
R_S8_34|4|B _S8_34|A4 _S8_34|4|MID_SHUNT  2.7439617672
L_S8_34|4|RB _S8_34|4|MID_SHUNT 0  1.550338398468e-12
B_S8_34|T|1 _S8_34|T1 _S8_34|T|MID_SERIES JJMIT AREA=2.5
L_S8_34|T|P _S8_34|T|MID_SERIES 0  2e-13
R_S8_34|T|B _S8_34|T1 _S8_34|T|MID_SHUNT  2.7439617672
L_S8_34|T|RB _S8_34|T|MID_SHUNT 0  1.550338398468e-12
B_S8_34|45|1 _S8_34|T2 _S8_34|A4 JJMIT AREA=1.7857142857142858
R_S8_34|45|B _S8_34|T2 _S8_34|45|MID_SHUNT  3.84154647408
L_S8_34|45|RB _S8_34|45|MID_SHUNT _S8_34|A4  2.1704737578552e-12
B_S8_34|6|1 _S8_34|Q1 _S8_34|6|MID_SERIES JJMIT AREA=2.5
L_S8_34|6|P _S8_34|6|MID_SERIES 0  2e-13
R_S8_34|6|B _S8_34|Q1 _S8_34|6|MID_SHUNT  2.7439617672
L_S8_34|6|RB _S8_34|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_S0_4|_TX|1 _PTL_S0_4|_TX|1 _PTL_S0_4|_TX|2 JJMIT AREA=2.5
B_PTL_S0_4|_TX|2 _PTL_S0_4|_TX|4 _PTL_S0_4|_TX|5 JJMIT AREA=2.5
I_PTL_S0_4|_TX|B1 0 _PTL_S0_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S0_4|_TX|B2 0 _PTL_S0_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S0_4|_TX|B1 _PTL_S0_4|_TX|1 _PTL_S0_4|_TX|3  1.684e-12
L_PTL_S0_4|_TX|B2 _PTL_S0_4|_TX|4 _PTL_S0_4|_TX|6  3.596e-12
L_PTL_S0_4|_TX|1 S0_4_TX _PTL_S0_4|_TX|1  2.063e-12
L_PTL_S0_4|_TX|2 _PTL_S0_4|_TX|1 _PTL_S0_4|_TX|4  4.123e-12
L_PTL_S0_4|_TX|3 _PTL_S0_4|_TX|4 _PTL_S0_4|_TX|7  2.193e-12
R_PTL_S0_4|_TX|D _PTL_S0_4|_TX|7 _PTL_S0_4|A_PTL  1.36
L_PTL_S0_4|_TX|P1 _PTL_S0_4|_TX|2 0  5.254e-13
L_PTL_S0_4|_TX|P2 _PTL_S0_4|_TX|5 0  5.141e-13
R_PTL_S0_4|_TX|B1 _PTL_S0_4|_TX|1 _PTL_S0_4|_TX|101  2.7439617672
R_PTL_S0_4|_TX|B2 _PTL_S0_4|_TX|4 _PTL_S0_4|_TX|104  2.7439617672
L_PTL_S0_4|_TX|RB1 _PTL_S0_4|_TX|101 0  1.550338398468e-12
L_PTL_S0_4|_TX|RB2 _PTL_S0_4|_TX|104 0  1.550338398468e-12
B_PTL_S0_4|_RX|1 _PTL_S0_4|_RX|1 _PTL_S0_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S0_4|_RX|2 _PTL_S0_4|_RX|4 _PTL_S0_4|_RX|5 JJMIT AREA=2.0
B_PTL_S0_4|_RX|3 _PTL_S0_4|_RX|7 _PTL_S0_4|_RX|8 JJMIT AREA=2.5
I_PTL_S0_4|_RX|B1 0 _PTL_S0_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S0_4|_RX|B1 _PTL_S0_4|_RX|1 _PTL_S0_4|_RX|3  2.777e-12
I_PTL_S0_4|_RX|B2 0 _PTL_S0_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S0_4|_RX|B2 _PTL_S0_4|_RX|4 _PTL_S0_4|_RX|6  2.685e-12
I_PTL_S0_4|_RX|B3 0 _PTL_S0_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S0_4|_RX|B3 _PTL_S0_4|_RX|7 _PTL_S0_4|_RX|9  2.764e-12
L_PTL_S0_4|_RX|1 _PTL_S0_4|A_PTL _PTL_S0_4|_RX|1  1.346e-12
L_PTL_S0_4|_RX|2 _PTL_S0_4|_RX|1 _PTL_S0_4|_RX|4  6.348e-12
L_PTL_S0_4|_RX|3 _PTL_S0_4|_RX|4 _PTL_S0_4|_RX|7  5.197e-12
L_PTL_S0_4|_RX|4 _PTL_S0_4|_RX|7 S0_4  2.058e-12
L_PTL_S0_4|_RX|P1 _PTL_S0_4|_RX|2 0  4.795e-13
L_PTL_S0_4|_RX|P2 _PTL_S0_4|_RX|5 0  5.431e-13
L_PTL_S0_4|_RX|P3 _PTL_S0_4|_RX|8 0  5.339e-13
R_PTL_S0_4|_RX|B1 _PTL_S0_4|_RX|1 _PTL_S0_4|_RX|101  4.225701121488
R_PTL_S0_4|_RX|B2 _PTL_S0_4|_RX|4 _PTL_S0_4|_RX|104  3.429952209
R_PTL_S0_4|_RX|B3 _PTL_S0_4|_RX|7 _PTL_S0_4|_RX|107  2.7439617672
L_PTL_S0_4|_RX|RB1 _PTL_S0_4|_RX|101 0  2.38752113364072e-12
L_PTL_S0_4|_RX|RB2 _PTL_S0_4|_RX|104 0  1.937922998085e-12
L_PTL_S0_4|_RX|RB3 _PTL_S0_4|_RX|107 0  1.550338398468e-12
B_PTL_S1_4|_TX|1 _PTL_S1_4|_TX|1 _PTL_S1_4|_TX|2 JJMIT AREA=2.5
B_PTL_S1_4|_TX|2 _PTL_S1_4|_TX|4 _PTL_S1_4|_TX|5 JJMIT AREA=2.5
I_PTL_S1_4|_TX|B1 0 _PTL_S1_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S1_4|_TX|B2 0 _PTL_S1_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S1_4|_TX|B1 _PTL_S1_4|_TX|1 _PTL_S1_4|_TX|3  1.684e-12
L_PTL_S1_4|_TX|B2 _PTL_S1_4|_TX|4 _PTL_S1_4|_TX|6  3.596e-12
L_PTL_S1_4|_TX|1 S1_4_TX _PTL_S1_4|_TX|1  2.063e-12
L_PTL_S1_4|_TX|2 _PTL_S1_4|_TX|1 _PTL_S1_4|_TX|4  4.123e-12
L_PTL_S1_4|_TX|3 _PTL_S1_4|_TX|4 _PTL_S1_4|_TX|7  2.193e-12
R_PTL_S1_4|_TX|D _PTL_S1_4|_TX|7 _PTL_S1_4|A_PTL  1.36
L_PTL_S1_4|_TX|P1 _PTL_S1_4|_TX|2 0  5.254e-13
L_PTL_S1_4|_TX|P2 _PTL_S1_4|_TX|5 0  5.141e-13
R_PTL_S1_4|_TX|B1 _PTL_S1_4|_TX|1 _PTL_S1_4|_TX|101  2.7439617672
R_PTL_S1_4|_TX|B2 _PTL_S1_4|_TX|4 _PTL_S1_4|_TX|104  2.7439617672
L_PTL_S1_4|_TX|RB1 _PTL_S1_4|_TX|101 0  1.550338398468e-12
L_PTL_S1_4|_TX|RB2 _PTL_S1_4|_TX|104 0  1.550338398468e-12
B_PTL_S1_4|_RX|1 _PTL_S1_4|_RX|1 _PTL_S1_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S1_4|_RX|2 _PTL_S1_4|_RX|4 _PTL_S1_4|_RX|5 JJMIT AREA=2.0
B_PTL_S1_4|_RX|3 _PTL_S1_4|_RX|7 _PTL_S1_4|_RX|8 JJMIT AREA=2.5
I_PTL_S1_4|_RX|B1 0 _PTL_S1_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S1_4|_RX|B1 _PTL_S1_4|_RX|1 _PTL_S1_4|_RX|3  2.777e-12
I_PTL_S1_4|_RX|B2 0 _PTL_S1_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S1_4|_RX|B2 _PTL_S1_4|_RX|4 _PTL_S1_4|_RX|6  2.685e-12
I_PTL_S1_4|_RX|B3 0 _PTL_S1_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S1_4|_RX|B3 _PTL_S1_4|_RX|7 _PTL_S1_4|_RX|9  2.764e-12
L_PTL_S1_4|_RX|1 _PTL_S1_4|A_PTL _PTL_S1_4|_RX|1  1.346e-12
L_PTL_S1_4|_RX|2 _PTL_S1_4|_RX|1 _PTL_S1_4|_RX|4  6.348e-12
L_PTL_S1_4|_RX|3 _PTL_S1_4|_RX|4 _PTL_S1_4|_RX|7  5.197e-12
L_PTL_S1_4|_RX|4 _PTL_S1_4|_RX|7 S1_4  2.058e-12
L_PTL_S1_4|_RX|P1 _PTL_S1_4|_RX|2 0  4.795e-13
L_PTL_S1_4|_RX|P2 _PTL_S1_4|_RX|5 0  5.431e-13
L_PTL_S1_4|_RX|P3 _PTL_S1_4|_RX|8 0  5.339e-13
R_PTL_S1_4|_RX|B1 _PTL_S1_4|_RX|1 _PTL_S1_4|_RX|101  4.225701121488
R_PTL_S1_4|_RX|B2 _PTL_S1_4|_RX|4 _PTL_S1_4|_RX|104  3.429952209
R_PTL_S1_4|_RX|B3 _PTL_S1_4|_RX|7 _PTL_S1_4|_RX|107  2.7439617672
L_PTL_S1_4|_RX|RB1 _PTL_S1_4|_RX|101 0  2.38752113364072e-12
L_PTL_S1_4|_RX|RB2 _PTL_S1_4|_RX|104 0  1.937922998085e-12
L_PTL_S1_4|_RX|RB3 _PTL_S1_4|_RX|107 0  1.550338398468e-12
B_PTL_S2_4|_TX|1 _PTL_S2_4|_TX|1 _PTL_S2_4|_TX|2 JJMIT AREA=2.5
B_PTL_S2_4|_TX|2 _PTL_S2_4|_TX|4 _PTL_S2_4|_TX|5 JJMIT AREA=2.5
I_PTL_S2_4|_TX|B1 0 _PTL_S2_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S2_4|_TX|B2 0 _PTL_S2_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S2_4|_TX|B1 _PTL_S2_4|_TX|1 _PTL_S2_4|_TX|3  1.684e-12
L_PTL_S2_4|_TX|B2 _PTL_S2_4|_TX|4 _PTL_S2_4|_TX|6  3.596e-12
L_PTL_S2_4|_TX|1 S2_4_TX _PTL_S2_4|_TX|1  2.063e-12
L_PTL_S2_4|_TX|2 _PTL_S2_4|_TX|1 _PTL_S2_4|_TX|4  4.123e-12
L_PTL_S2_4|_TX|3 _PTL_S2_4|_TX|4 _PTL_S2_4|_TX|7  2.193e-12
R_PTL_S2_4|_TX|D _PTL_S2_4|_TX|7 _PTL_S2_4|A_PTL  1.36
L_PTL_S2_4|_TX|P1 _PTL_S2_4|_TX|2 0  5.254e-13
L_PTL_S2_4|_TX|P2 _PTL_S2_4|_TX|5 0  5.141e-13
R_PTL_S2_4|_TX|B1 _PTL_S2_4|_TX|1 _PTL_S2_4|_TX|101  2.7439617672
R_PTL_S2_4|_TX|B2 _PTL_S2_4|_TX|4 _PTL_S2_4|_TX|104  2.7439617672
L_PTL_S2_4|_TX|RB1 _PTL_S2_4|_TX|101 0  1.550338398468e-12
L_PTL_S2_4|_TX|RB2 _PTL_S2_4|_TX|104 0  1.550338398468e-12
B_PTL_S2_4|_RX|1 _PTL_S2_4|_RX|1 _PTL_S2_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S2_4|_RX|2 _PTL_S2_4|_RX|4 _PTL_S2_4|_RX|5 JJMIT AREA=2.0
B_PTL_S2_4|_RX|3 _PTL_S2_4|_RX|7 _PTL_S2_4|_RX|8 JJMIT AREA=2.5
I_PTL_S2_4|_RX|B1 0 _PTL_S2_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S2_4|_RX|B1 _PTL_S2_4|_RX|1 _PTL_S2_4|_RX|3  2.777e-12
I_PTL_S2_4|_RX|B2 0 _PTL_S2_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S2_4|_RX|B2 _PTL_S2_4|_RX|4 _PTL_S2_4|_RX|6  2.685e-12
I_PTL_S2_4|_RX|B3 0 _PTL_S2_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S2_4|_RX|B3 _PTL_S2_4|_RX|7 _PTL_S2_4|_RX|9  2.764e-12
L_PTL_S2_4|_RX|1 _PTL_S2_4|A_PTL _PTL_S2_4|_RX|1  1.346e-12
L_PTL_S2_4|_RX|2 _PTL_S2_4|_RX|1 _PTL_S2_4|_RX|4  6.348e-12
L_PTL_S2_4|_RX|3 _PTL_S2_4|_RX|4 _PTL_S2_4|_RX|7  5.197e-12
L_PTL_S2_4|_RX|4 _PTL_S2_4|_RX|7 S2_4  2.058e-12
L_PTL_S2_4|_RX|P1 _PTL_S2_4|_RX|2 0  4.795e-13
L_PTL_S2_4|_RX|P2 _PTL_S2_4|_RX|5 0  5.431e-13
L_PTL_S2_4|_RX|P3 _PTL_S2_4|_RX|8 0  5.339e-13
R_PTL_S2_4|_RX|B1 _PTL_S2_4|_RX|1 _PTL_S2_4|_RX|101  4.225701121488
R_PTL_S2_4|_RX|B2 _PTL_S2_4|_RX|4 _PTL_S2_4|_RX|104  3.429952209
R_PTL_S2_4|_RX|B3 _PTL_S2_4|_RX|7 _PTL_S2_4|_RX|107  2.7439617672
L_PTL_S2_4|_RX|RB1 _PTL_S2_4|_RX|101 0  2.38752113364072e-12
L_PTL_S2_4|_RX|RB2 _PTL_S2_4|_RX|104 0  1.937922998085e-12
L_PTL_S2_4|_RX|RB3 _PTL_S2_4|_RX|107 0  1.550338398468e-12
B_PTL_S3_4|_TX|1 _PTL_S3_4|_TX|1 _PTL_S3_4|_TX|2 JJMIT AREA=2.5
B_PTL_S3_4|_TX|2 _PTL_S3_4|_TX|4 _PTL_S3_4|_TX|5 JJMIT AREA=2.5
I_PTL_S3_4|_TX|B1 0 _PTL_S3_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S3_4|_TX|B2 0 _PTL_S3_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S3_4|_TX|B1 _PTL_S3_4|_TX|1 _PTL_S3_4|_TX|3  1.684e-12
L_PTL_S3_4|_TX|B2 _PTL_S3_4|_TX|4 _PTL_S3_4|_TX|6  3.596e-12
L_PTL_S3_4|_TX|1 S3_4_TX _PTL_S3_4|_TX|1  2.063e-12
L_PTL_S3_4|_TX|2 _PTL_S3_4|_TX|1 _PTL_S3_4|_TX|4  4.123e-12
L_PTL_S3_4|_TX|3 _PTL_S3_4|_TX|4 _PTL_S3_4|_TX|7  2.193e-12
R_PTL_S3_4|_TX|D _PTL_S3_4|_TX|7 _PTL_S3_4|A_PTL  1.36
L_PTL_S3_4|_TX|P1 _PTL_S3_4|_TX|2 0  5.254e-13
L_PTL_S3_4|_TX|P2 _PTL_S3_4|_TX|5 0  5.141e-13
R_PTL_S3_4|_TX|B1 _PTL_S3_4|_TX|1 _PTL_S3_4|_TX|101  2.7439617672
R_PTL_S3_4|_TX|B2 _PTL_S3_4|_TX|4 _PTL_S3_4|_TX|104  2.7439617672
L_PTL_S3_4|_TX|RB1 _PTL_S3_4|_TX|101 0  1.550338398468e-12
L_PTL_S3_4|_TX|RB2 _PTL_S3_4|_TX|104 0  1.550338398468e-12
B_PTL_S3_4|_RX|1 _PTL_S3_4|_RX|1 _PTL_S3_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S3_4|_RX|2 _PTL_S3_4|_RX|4 _PTL_S3_4|_RX|5 JJMIT AREA=2.0
B_PTL_S3_4|_RX|3 _PTL_S3_4|_RX|7 _PTL_S3_4|_RX|8 JJMIT AREA=2.5
I_PTL_S3_4|_RX|B1 0 _PTL_S3_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S3_4|_RX|B1 _PTL_S3_4|_RX|1 _PTL_S3_4|_RX|3  2.777e-12
I_PTL_S3_4|_RX|B2 0 _PTL_S3_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S3_4|_RX|B2 _PTL_S3_4|_RX|4 _PTL_S3_4|_RX|6  2.685e-12
I_PTL_S3_4|_RX|B3 0 _PTL_S3_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S3_4|_RX|B3 _PTL_S3_4|_RX|7 _PTL_S3_4|_RX|9  2.764e-12
L_PTL_S3_4|_RX|1 _PTL_S3_4|A_PTL _PTL_S3_4|_RX|1  1.346e-12
L_PTL_S3_4|_RX|2 _PTL_S3_4|_RX|1 _PTL_S3_4|_RX|4  6.348e-12
L_PTL_S3_4|_RX|3 _PTL_S3_4|_RX|4 _PTL_S3_4|_RX|7  5.197e-12
L_PTL_S3_4|_RX|4 _PTL_S3_4|_RX|7 S3_4  2.058e-12
L_PTL_S3_4|_RX|P1 _PTL_S3_4|_RX|2 0  4.795e-13
L_PTL_S3_4|_RX|P2 _PTL_S3_4|_RX|5 0  5.431e-13
L_PTL_S3_4|_RX|P3 _PTL_S3_4|_RX|8 0  5.339e-13
R_PTL_S3_4|_RX|B1 _PTL_S3_4|_RX|1 _PTL_S3_4|_RX|101  4.225701121488
R_PTL_S3_4|_RX|B2 _PTL_S3_4|_RX|4 _PTL_S3_4|_RX|104  3.429952209
R_PTL_S3_4|_RX|B3 _PTL_S3_4|_RX|7 _PTL_S3_4|_RX|107  2.7439617672
L_PTL_S3_4|_RX|RB1 _PTL_S3_4|_RX|101 0  2.38752113364072e-12
L_PTL_S3_4|_RX|RB2 _PTL_S3_4|_RX|104 0  1.937922998085e-12
L_PTL_S3_4|_RX|RB3 _PTL_S3_4|_RX|107 0  1.550338398468e-12
B_PTL_S4_4|_TX|1 _PTL_S4_4|_TX|1 _PTL_S4_4|_TX|2 JJMIT AREA=2.5
B_PTL_S4_4|_TX|2 _PTL_S4_4|_TX|4 _PTL_S4_4|_TX|5 JJMIT AREA=2.5
I_PTL_S4_4|_TX|B1 0 _PTL_S4_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S4_4|_TX|B2 0 _PTL_S4_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S4_4|_TX|B1 _PTL_S4_4|_TX|1 _PTL_S4_4|_TX|3  1.684e-12
L_PTL_S4_4|_TX|B2 _PTL_S4_4|_TX|4 _PTL_S4_4|_TX|6  3.596e-12
L_PTL_S4_4|_TX|1 S4_4_TX _PTL_S4_4|_TX|1  2.063e-12
L_PTL_S4_4|_TX|2 _PTL_S4_4|_TX|1 _PTL_S4_4|_TX|4  4.123e-12
L_PTL_S4_4|_TX|3 _PTL_S4_4|_TX|4 _PTL_S4_4|_TX|7  2.193e-12
R_PTL_S4_4|_TX|D _PTL_S4_4|_TX|7 _PTL_S4_4|A_PTL  1.36
L_PTL_S4_4|_TX|P1 _PTL_S4_4|_TX|2 0  5.254e-13
L_PTL_S4_4|_TX|P2 _PTL_S4_4|_TX|5 0  5.141e-13
R_PTL_S4_4|_TX|B1 _PTL_S4_4|_TX|1 _PTL_S4_4|_TX|101  2.7439617672
R_PTL_S4_4|_TX|B2 _PTL_S4_4|_TX|4 _PTL_S4_4|_TX|104  2.7439617672
L_PTL_S4_4|_TX|RB1 _PTL_S4_4|_TX|101 0  1.550338398468e-12
L_PTL_S4_4|_TX|RB2 _PTL_S4_4|_TX|104 0  1.550338398468e-12
B_PTL_S4_4|_RX|1 _PTL_S4_4|_RX|1 _PTL_S4_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S4_4|_RX|2 _PTL_S4_4|_RX|4 _PTL_S4_4|_RX|5 JJMIT AREA=2.0
B_PTL_S4_4|_RX|3 _PTL_S4_4|_RX|7 _PTL_S4_4|_RX|8 JJMIT AREA=2.5
I_PTL_S4_4|_RX|B1 0 _PTL_S4_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S4_4|_RX|B1 _PTL_S4_4|_RX|1 _PTL_S4_4|_RX|3  2.777e-12
I_PTL_S4_4|_RX|B2 0 _PTL_S4_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S4_4|_RX|B2 _PTL_S4_4|_RX|4 _PTL_S4_4|_RX|6  2.685e-12
I_PTL_S4_4|_RX|B3 0 _PTL_S4_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S4_4|_RX|B3 _PTL_S4_4|_RX|7 _PTL_S4_4|_RX|9  2.764e-12
L_PTL_S4_4|_RX|1 _PTL_S4_4|A_PTL _PTL_S4_4|_RX|1  1.346e-12
L_PTL_S4_4|_RX|2 _PTL_S4_4|_RX|1 _PTL_S4_4|_RX|4  6.348e-12
L_PTL_S4_4|_RX|3 _PTL_S4_4|_RX|4 _PTL_S4_4|_RX|7  5.197e-12
L_PTL_S4_4|_RX|4 _PTL_S4_4|_RX|7 S4_4  2.058e-12
L_PTL_S4_4|_RX|P1 _PTL_S4_4|_RX|2 0  4.795e-13
L_PTL_S4_4|_RX|P2 _PTL_S4_4|_RX|5 0  5.431e-13
L_PTL_S4_4|_RX|P3 _PTL_S4_4|_RX|8 0  5.339e-13
R_PTL_S4_4|_RX|B1 _PTL_S4_4|_RX|1 _PTL_S4_4|_RX|101  4.225701121488
R_PTL_S4_4|_RX|B2 _PTL_S4_4|_RX|4 _PTL_S4_4|_RX|104  3.429952209
R_PTL_S4_4|_RX|B3 _PTL_S4_4|_RX|7 _PTL_S4_4|_RX|107  2.7439617672
L_PTL_S4_4|_RX|RB1 _PTL_S4_4|_RX|101 0  2.38752113364072e-12
L_PTL_S4_4|_RX|RB2 _PTL_S4_4|_RX|104 0  1.937922998085e-12
L_PTL_S4_4|_RX|RB3 _PTL_S4_4|_RX|107 0  1.550338398468e-12
B_PTL_S5_4|_TX|1 _PTL_S5_4|_TX|1 _PTL_S5_4|_TX|2 JJMIT AREA=2.5
B_PTL_S5_4|_TX|2 _PTL_S5_4|_TX|4 _PTL_S5_4|_TX|5 JJMIT AREA=2.5
I_PTL_S5_4|_TX|B1 0 _PTL_S5_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S5_4|_TX|B2 0 _PTL_S5_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S5_4|_TX|B1 _PTL_S5_4|_TX|1 _PTL_S5_4|_TX|3  1.684e-12
L_PTL_S5_4|_TX|B2 _PTL_S5_4|_TX|4 _PTL_S5_4|_TX|6  3.596e-12
L_PTL_S5_4|_TX|1 S5_4_TX _PTL_S5_4|_TX|1  2.063e-12
L_PTL_S5_4|_TX|2 _PTL_S5_4|_TX|1 _PTL_S5_4|_TX|4  4.123e-12
L_PTL_S5_4|_TX|3 _PTL_S5_4|_TX|4 _PTL_S5_4|_TX|7  2.193e-12
R_PTL_S5_4|_TX|D _PTL_S5_4|_TX|7 _PTL_S5_4|A_PTL  1.36
L_PTL_S5_4|_TX|P1 _PTL_S5_4|_TX|2 0  5.254e-13
L_PTL_S5_4|_TX|P2 _PTL_S5_4|_TX|5 0  5.141e-13
R_PTL_S5_4|_TX|B1 _PTL_S5_4|_TX|1 _PTL_S5_4|_TX|101  2.7439617672
R_PTL_S5_4|_TX|B2 _PTL_S5_4|_TX|4 _PTL_S5_4|_TX|104  2.7439617672
L_PTL_S5_4|_TX|RB1 _PTL_S5_4|_TX|101 0  1.550338398468e-12
L_PTL_S5_4|_TX|RB2 _PTL_S5_4|_TX|104 0  1.550338398468e-12
B_PTL_S5_4|_RX|1 _PTL_S5_4|_RX|1 _PTL_S5_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S5_4|_RX|2 _PTL_S5_4|_RX|4 _PTL_S5_4|_RX|5 JJMIT AREA=2.0
B_PTL_S5_4|_RX|3 _PTL_S5_4|_RX|7 _PTL_S5_4|_RX|8 JJMIT AREA=2.5
I_PTL_S5_4|_RX|B1 0 _PTL_S5_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S5_4|_RX|B1 _PTL_S5_4|_RX|1 _PTL_S5_4|_RX|3  2.777e-12
I_PTL_S5_4|_RX|B2 0 _PTL_S5_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S5_4|_RX|B2 _PTL_S5_4|_RX|4 _PTL_S5_4|_RX|6  2.685e-12
I_PTL_S5_4|_RX|B3 0 _PTL_S5_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S5_4|_RX|B3 _PTL_S5_4|_RX|7 _PTL_S5_4|_RX|9  2.764e-12
L_PTL_S5_4|_RX|1 _PTL_S5_4|A_PTL _PTL_S5_4|_RX|1  1.346e-12
L_PTL_S5_4|_RX|2 _PTL_S5_4|_RX|1 _PTL_S5_4|_RX|4  6.348e-12
L_PTL_S5_4|_RX|3 _PTL_S5_4|_RX|4 _PTL_S5_4|_RX|7  5.197e-12
L_PTL_S5_4|_RX|4 _PTL_S5_4|_RX|7 S5_4  2.058e-12
L_PTL_S5_4|_RX|P1 _PTL_S5_4|_RX|2 0  4.795e-13
L_PTL_S5_4|_RX|P2 _PTL_S5_4|_RX|5 0  5.431e-13
L_PTL_S5_4|_RX|P3 _PTL_S5_4|_RX|8 0  5.339e-13
R_PTL_S5_4|_RX|B1 _PTL_S5_4|_RX|1 _PTL_S5_4|_RX|101  4.225701121488
R_PTL_S5_4|_RX|B2 _PTL_S5_4|_RX|4 _PTL_S5_4|_RX|104  3.429952209
R_PTL_S5_4|_RX|B3 _PTL_S5_4|_RX|7 _PTL_S5_4|_RX|107  2.7439617672
L_PTL_S5_4|_RX|RB1 _PTL_S5_4|_RX|101 0  2.38752113364072e-12
L_PTL_S5_4|_RX|RB2 _PTL_S5_4|_RX|104 0  1.937922998085e-12
L_PTL_S5_4|_RX|RB3 _PTL_S5_4|_RX|107 0  1.550338398468e-12
B_PTL_S6_4|_TX|1 _PTL_S6_4|_TX|1 _PTL_S6_4|_TX|2 JJMIT AREA=2.5
B_PTL_S6_4|_TX|2 _PTL_S6_4|_TX|4 _PTL_S6_4|_TX|5 JJMIT AREA=2.5
I_PTL_S6_4|_TX|B1 0 _PTL_S6_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S6_4|_TX|B2 0 _PTL_S6_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S6_4|_TX|B1 _PTL_S6_4|_TX|1 _PTL_S6_4|_TX|3  1.684e-12
L_PTL_S6_4|_TX|B2 _PTL_S6_4|_TX|4 _PTL_S6_4|_TX|6  3.596e-12
L_PTL_S6_4|_TX|1 S6_4_TX _PTL_S6_4|_TX|1  2.063e-12
L_PTL_S6_4|_TX|2 _PTL_S6_4|_TX|1 _PTL_S6_4|_TX|4  4.123e-12
L_PTL_S6_4|_TX|3 _PTL_S6_4|_TX|4 _PTL_S6_4|_TX|7  2.193e-12
R_PTL_S6_4|_TX|D _PTL_S6_4|_TX|7 _PTL_S6_4|A_PTL  1.36
L_PTL_S6_4|_TX|P1 _PTL_S6_4|_TX|2 0  5.254e-13
L_PTL_S6_4|_TX|P2 _PTL_S6_4|_TX|5 0  5.141e-13
R_PTL_S6_4|_TX|B1 _PTL_S6_4|_TX|1 _PTL_S6_4|_TX|101  2.7439617672
R_PTL_S6_4|_TX|B2 _PTL_S6_4|_TX|4 _PTL_S6_4|_TX|104  2.7439617672
L_PTL_S6_4|_TX|RB1 _PTL_S6_4|_TX|101 0  1.550338398468e-12
L_PTL_S6_4|_TX|RB2 _PTL_S6_4|_TX|104 0  1.550338398468e-12
B_PTL_S6_4|_RX|1 _PTL_S6_4|_RX|1 _PTL_S6_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S6_4|_RX|2 _PTL_S6_4|_RX|4 _PTL_S6_4|_RX|5 JJMIT AREA=2.0
B_PTL_S6_4|_RX|3 _PTL_S6_4|_RX|7 _PTL_S6_4|_RX|8 JJMIT AREA=2.5
I_PTL_S6_4|_RX|B1 0 _PTL_S6_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S6_4|_RX|B1 _PTL_S6_4|_RX|1 _PTL_S6_4|_RX|3  2.777e-12
I_PTL_S6_4|_RX|B2 0 _PTL_S6_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S6_4|_RX|B2 _PTL_S6_4|_RX|4 _PTL_S6_4|_RX|6  2.685e-12
I_PTL_S6_4|_RX|B3 0 _PTL_S6_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S6_4|_RX|B3 _PTL_S6_4|_RX|7 _PTL_S6_4|_RX|9  2.764e-12
L_PTL_S6_4|_RX|1 _PTL_S6_4|A_PTL _PTL_S6_4|_RX|1  1.346e-12
L_PTL_S6_4|_RX|2 _PTL_S6_4|_RX|1 _PTL_S6_4|_RX|4  6.348e-12
L_PTL_S6_4|_RX|3 _PTL_S6_4|_RX|4 _PTL_S6_4|_RX|7  5.197e-12
L_PTL_S6_4|_RX|4 _PTL_S6_4|_RX|7 S6_4  2.058e-12
L_PTL_S6_4|_RX|P1 _PTL_S6_4|_RX|2 0  4.795e-13
L_PTL_S6_4|_RX|P2 _PTL_S6_4|_RX|5 0  5.431e-13
L_PTL_S6_4|_RX|P3 _PTL_S6_4|_RX|8 0  5.339e-13
R_PTL_S6_4|_RX|B1 _PTL_S6_4|_RX|1 _PTL_S6_4|_RX|101  4.225701121488
R_PTL_S6_4|_RX|B2 _PTL_S6_4|_RX|4 _PTL_S6_4|_RX|104  3.429952209
R_PTL_S6_4|_RX|B3 _PTL_S6_4|_RX|7 _PTL_S6_4|_RX|107  2.7439617672
L_PTL_S6_4|_RX|RB1 _PTL_S6_4|_RX|101 0  2.38752113364072e-12
L_PTL_S6_4|_RX|RB2 _PTL_S6_4|_RX|104 0  1.937922998085e-12
L_PTL_S6_4|_RX|RB3 _PTL_S6_4|_RX|107 0  1.550338398468e-12
B_PTL_G6_4|_TX|1 _PTL_G6_4|_TX|1 _PTL_G6_4|_TX|2 JJMIT AREA=2.5
B_PTL_G6_4|_TX|2 _PTL_G6_4|_TX|4 _PTL_G6_4|_TX|5 JJMIT AREA=2.5
I_PTL_G6_4|_TX|B1 0 _PTL_G6_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_G6_4|_TX|B2 0 _PTL_G6_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_G6_4|_TX|B1 _PTL_G6_4|_TX|1 _PTL_G6_4|_TX|3  1.684e-12
L_PTL_G6_4|_TX|B2 _PTL_G6_4|_TX|4 _PTL_G6_4|_TX|6  3.596e-12
L_PTL_G6_4|_TX|1 G6_4_TX _PTL_G6_4|_TX|1  2.063e-12
L_PTL_G6_4|_TX|2 _PTL_G6_4|_TX|1 _PTL_G6_4|_TX|4  4.123e-12
L_PTL_G6_4|_TX|3 _PTL_G6_4|_TX|4 _PTL_G6_4|_TX|7  2.193e-12
R_PTL_G6_4|_TX|D _PTL_G6_4|_TX|7 _PTL_G6_4|A_PTL  1.36
L_PTL_G6_4|_TX|P1 _PTL_G6_4|_TX|2 0  5.254e-13
L_PTL_G6_4|_TX|P2 _PTL_G6_4|_TX|5 0  5.141e-13
R_PTL_G6_4|_TX|B1 _PTL_G6_4|_TX|1 _PTL_G6_4|_TX|101  2.7439617672
R_PTL_G6_4|_TX|B2 _PTL_G6_4|_TX|4 _PTL_G6_4|_TX|104  2.7439617672
L_PTL_G6_4|_TX|RB1 _PTL_G6_4|_TX|101 0  1.550338398468e-12
L_PTL_G6_4|_TX|RB2 _PTL_G6_4|_TX|104 0  1.550338398468e-12
B_PTL_G6_4|_RX|1 _PTL_G6_4|_RX|1 _PTL_G6_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_G6_4|_RX|2 _PTL_G6_4|_RX|4 _PTL_G6_4|_RX|5 JJMIT AREA=2.0
B_PTL_G6_4|_RX|3 _PTL_G6_4|_RX|7 _PTL_G6_4|_RX|8 JJMIT AREA=2.5
I_PTL_G6_4|_RX|B1 0 _PTL_G6_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_G6_4|_RX|B1 _PTL_G6_4|_RX|1 _PTL_G6_4|_RX|3  2.777e-12
I_PTL_G6_4|_RX|B2 0 _PTL_G6_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_G6_4|_RX|B2 _PTL_G6_4|_RX|4 _PTL_G6_4|_RX|6  2.685e-12
I_PTL_G6_4|_RX|B3 0 _PTL_G6_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_G6_4|_RX|B3 _PTL_G6_4|_RX|7 _PTL_G6_4|_RX|9  2.764e-12
L_PTL_G6_4|_RX|1 _PTL_G6_4|A_PTL _PTL_G6_4|_RX|1  1.346e-12
L_PTL_G6_4|_RX|2 _PTL_G6_4|_RX|1 _PTL_G6_4|_RX|4  6.348e-12
L_PTL_G6_4|_RX|3 _PTL_G6_4|_RX|4 _PTL_G6_4|_RX|7  5.197e-12
L_PTL_G6_4|_RX|4 _PTL_G6_4|_RX|7 G6_4_OUT  2.058e-12
L_PTL_G6_4|_RX|P1 _PTL_G6_4|_RX|2 0  4.795e-13
L_PTL_G6_4|_RX|P2 _PTL_G6_4|_RX|5 0  5.431e-13
L_PTL_G6_4|_RX|P3 _PTL_G6_4|_RX|8 0  5.339e-13
R_PTL_G6_4|_RX|B1 _PTL_G6_4|_RX|1 _PTL_G6_4|_RX|101  4.225701121488
R_PTL_G6_4|_RX|B2 _PTL_G6_4|_RX|4 _PTL_G6_4|_RX|104  3.429952209
R_PTL_G6_4|_RX|B3 _PTL_G6_4|_RX|7 _PTL_G6_4|_RX|107  2.7439617672
L_PTL_G6_4|_RX|RB1 _PTL_G6_4|_RX|101 0  2.38752113364072e-12
L_PTL_G6_4|_RX|RB2 _PTL_G6_4|_RX|104 0  1.937922998085e-12
L_PTL_G6_4|_RX|RB3 _PTL_G6_4|_RX|107 0  1.550338398468e-12
B_PTL_IP7_4|_TX|1 _PTL_IP7_4|_TX|1 _PTL_IP7_4|_TX|2 JJMIT AREA=2.5
B_PTL_IP7_4|_TX|2 _PTL_IP7_4|_TX|4 _PTL_IP7_4|_TX|5 JJMIT AREA=2.5
I_PTL_IP7_4|_TX|B1 0 _PTL_IP7_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_IP7_4|_TX|B2 0 _PTL_IP7_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_4|_TX|B1 _PTL_IP7_4|_TX|1 _PTL_IP7_4|_TX|3  1.684e-12
L_PTL_IP7_4|_TX|B2 _PTL_IP7_4|_TX|4 _PTL_IP7_4|_TX|6  3.596e-12
L_PTL_IP7_4|_TX|1 IP7_4_OUT_TX _PTL_IP7_4|_TX|1  2.063e-12
L_PTL_IP7_4|_TX|2 _PTL_IP7_4|_TX|1 _PTL_IP7_4|_TX|4  4.123e-12
L_PTL_IP7_4|_TX|3 _PTL_IP7_4|_TX|4 _PTL_IP7_4|_TX|7  2.193e-12
R_PTL_IP7_4|_TX|D _PTL_IP7_4|_TX|7 _PTL_IP7_4|A_PTL  1.36
L_PTL_IP7_4|_TX|P1 _PTL_IP7_4|_TX|2 0  5.254e-13
L_PTL_IP7_4|_TX|P2 _PTL_IP7_4|_TX|5 0  5.141e-13
R_PTL_IP7_4|_TX|B1 _PTL_IP7_4|_TX|1 _PTL_IP7_4|_TX|101  2.7439617672
R_PTL_IP7_4|_TX|B2 _PTL_IP7_4|_TX|4 _PTL_IP7_4|_TX|104  2.7439617672
L_PTL_IP7_4|_TX|RB1 _PTL_IP7_4|_TX|101 0  1.550338398468e-12
L_PTL_IP7_4|_TX|RB2 _PTL_IP7_4|_TX|104 0  1.550338398468e-12
B_PTL_IP7_4|_RX|1 _PTL_IP7_4|_RX|1 _PTL_IP7_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_IP7_4|_RX|2 _PTL_IP7_4|_RX|4 _PTL_IP7_4|_RX|5 JJMIT AREA=2.0
B_PTL_IP7_4|_RX|3 _PTL_IP7_4|_RX|7 _PTL_IP7_4|_RX|8 JJMIT AREA=2.5
I_PTL_IP7_4|_RX|B1 0 _PTL_IP7_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_IP7_4|_RX|B1 _PTL_IP7_4|_RX|1 _PTL_IP7_4|_RX|3  2.777e-12
I_PTL_IP7_4|_RX|B2 0 _PTL_IP7_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_IP7_4|_RX|B2 _PTL_IP7_4|_RX|4 _PTL_IP7_4|_RX|6  2.685e-12
I_PTL_IP7_4|_RX|B3 0 _PTL_IP7_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_4|_RX|B3 _PTL_IP7_4|_RX|7 _PTL_IP7_4|_RX|9  2.764e-12
L_PTL_IP7_4|_RX|1 _PTL_IP7_4|A_PTL _PTL_IP7_4|_RX|1  1.346e-12
L_PTL_IP7_4|_RX|2 _PTL_IP7_4|_RX|1 _PTL_IP7_4|_RX|4  6.348e-12
L_PTL_IP7_4|_RX|3 _PTL_IP7_4|_RX|4 _PTL_IP7_4|_RX|7  5.197e-12
L_PTL_IP7_4|_RX|4 _PTL_IP7_4|_RX|7 IP7_4_OUT  2.058e-12
L_PTL_IP7_4|_RX|P1 _PTL_IP7_4|_RX|2 0  4.795e-13
L_PTL_IP7_4|_RX|P2 _PTL_IP7_4|_RX|5 0  5.431e-13
L_PTL_IP7_4|_RX|P3 _PTL_IP7_4|_RX|8 0  5.339e-13
R_PTL_IP7_4|_RX|B1 _PTL_IP7_4|_RX|1 _PTL_IP7_4|_RX|101  4.225701121488
R_PTL_IP7_4|_RX|B2 _PTL_IP7_4|_RX|4 _PTL_IP7_4|_RX|104  3.429952209
R_PTL_IP7_4|_RX|B3 _PTL_IP7_4|_RX|7 _PTL_IP7_4|_RX|107  2.7439617672
L_PTL_IP7_4|_RX|RB1 _PTL_IP7_4|_RX|101 0  2.38752113364072e-12
L_PTL_IP7_4|_RX|RB2 _PTL_IP7_4|_RX|104 0  1.937922998085e-12
L_PTL_IP7_4|_RX|RB3 _PTL_IP7_4|_RX|107 0  1.550338398468e-12
B_PTL_S8_4|_TX|1 _PTL_S8_4|_TX|1 _PTL_S8_4|_TX|2 JJMIT AREA=2.5
B_PTL_S8_4|_TX|2 _PTL_S8_4|_TX|4 _PTL_S8_4|_TX|5 JJMIT AREA=2.5
I_PTL_S8_4|_TX|B1 0 _PTL_S8_4|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S8_4|_TX|B2 0 _PTL_S8_4|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S8_4|_TX|B1 _PTL_S8_4|_TX|1 _PTL_S8_4|_TX|3  1.684e-12
L_PTL_S8_4|_TX|B2 _PTL_S8_4|_TX|4 _PTL_S8_4|_TX|6  3.596e-12
L_PTL_S8_4|_TX|1 S8_4_TX _PTL_S8_4|_TX|1  2.063e-12
L_PTL_S8_4|_TX|2 _PTL_S8_4|_TX|1 _PTL_S8_4|_TX|4  4.123e-12
L_PTL_S8_4|_TX|3 _PTL_S8_4|_TX|4 _PTL_S8_4|_TX|7  2.193e-12
R_PTL_S8_4|_TX|D _PTL_S8_4|_TX|7 _PTL_S8_4|A_PTL  1.36
L_PTL_S8_4|_TX|P1 _PTL_S8_4|_TX|2 0  5.254e-13
L_PTL_S8_4|_TX|P2 _PTL_S8_4|_TX|5 0  5.141e-13
R_PTL_S8_4|_TX|B1 _PTL_S8_4|_TX|1 _PTL_S8_4|_TX|101  2.7439617672
R_PTL_S8_4|_TX|B2 _PTL_S8_4|_TX|4 _PTL_S8_4|_TX|104  2.7439617672
L_PTL_S8_4|_TX|RB1 _PTL_S8_4|_TX|101 0  1.550338398468e-12
L_PTL_S8_4|_TX|RB2 _PTL_S8_4|_TX|104 0  1.550338398468e-12
B_PTL_S8_4|_RX|1 _PTL_S8_4|_RX|1 _PTL_S8_4|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S8_4|_RX|2 _PTL_S8_4|_RX|4 _PTL_S8_4|_RX|5 JJMIT AREA=2.0
B_PTL_S8_4|_RX|3 _PTL_S8_4|_RX|7 _PTL_S8_4|_RX|8 JJMIT AREA=2.5
I_PTL_S8_4|_RX|B1 0 _PTL_S8_4|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S8_4|_RX|B1 _PTL_S8_4|_RX|1 _PTL_S8_4|_RX|3  2.777e-12
I_PTL_S8_4|_RX|B2 0 _PTL_S8_4|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S8_4|_RX|B2 _PTL_S8_4|_RX|4 _PTL_S8_4|_RX|6  2.685e-12
I_PTL_S8_4|_RX|B3 0 _PTL_S8_4|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S8_4|_RX|B3 _PTL_S8_4|_RX|7 _PTL_S8_4|_RX|9  2.764e-12
L_PTL_S8_4|_RX|1 _PTL_S8_4|A_PTL _PTL_S8_4|_RX|1  1.346e-12
L_PTL_S8_4|_RX|2 _PTL_S8_4|_RX|1 _PTL_S8_4|_RX|4  6.348e-12
L_PTL_S8_4|_RX|3 _PTL_S8_4|_RX|4 _PTL_S8_4|_RX|7  5.197e-12
L_PTL_S8_4|_RX|4 _PTL_S8_4|_RX|7 S8_4  2.058e-12
L_PTL_S8_4|_RX|P1 _PTL_S8_4|_RX|2 0  4.795e-13
L_PTL_S8_4|_RX|P2 _PTL_S8_4|_RX|5 0  5.431e-13
L_PTL_S8_4|_RX|P3 _PTL_S8_4|_RX|8 0  5.339e-13
R_PTL_S8_4|_RX|B1 _PTL_S8_4|_RX|1 _PTL_S8_4|_RX|101  4.225701121488
R_PTL_S8_4|_RX|B2 _PTL_S8_4|_RX|4 _PTL_S8_4|_RX|104  3.429952209
R_PTL_S8_4|_RX|B3 _PTL_S8_4|_RX|7 _PTL_S8_4|_RX|107  2.7439617672
L_PTL_S8_4|_RX|RB1 _PTL_S8_4|_RX|101 0  2.38752113364072e-12
L_PTL_S8_4|_RX|RB2 _PTL_S8_4|_RX|104 0  1.937922998085e-12
L_PTL_S8_4|_RX|RB3 _PTL_S8_4|_RX|107 0  1.550338398468e-12
L_S0_45|I_1|B _S0_45|A1 _S0_45|I_1|MID  2e-12
I_S0_45|I_1|B 0 _S0_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0_45|I_3|B _S0_45|A3 _S0_45|I_3|MID  2e-12
I_S0_45|I_3|B 0 _S0_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0_45|I_T|B _S0_45|T1 _S0_45|I_T|MID  2e-12
I_S0_45|I_T|B 0 _S0_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0_45|I_6|B _S0_45|Q1 _S0_45|I_6|MID  2e-12
I_S0_45|I_6|B 0 _S0_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0_45|1|1 _S0_45|A1 _S0_45|1|MID_SERIES JJMIT AREA=2.5
L_S0_45|1|P _S0_45|1|MID_SERIES 0  2e-13
R_S0_45|1|B _S0_45|A1 _S0_45|1|MID_SHUNT  2.7439617672
L_S0_45|1|RB _S0_45|1|MID_SHUNT 0  1.550338398468e-12
B_S0_45|23|1 _S0_45|A2 _S0_45|A3 JJMIT AREA=1.7857142857142858
R_S0_45|23|B _S0_45|A2 _S0_45|23|MID_SHUNT  3.84154647408
L_S0_45|23|RB _S0_45|23|MID_SHUNT _S0_45|A3  2.1704737578552e-12
B_S0_45|3|1 _S0_45|A3 _S0_45|3|MID_SERIES JJMIT AREA=2.5
L_S0_45|3|P _S0_45|3|MID_SERIES 0  2e-13
R_S0_45|3|B _S0_45|A3 _S0_45|3|MID_SHUNT  2.7439617672
L_S0_45|3|RB _S0_45|3|MID_SHUNT 0  1.550338398468e-12
B_S0_45|4|1 _S0_45|A4 _S0_45|4|MID_SERIES JJMIT AREA=2.5
L_S0_45|4|P _S0_45|4|MID_SERIES 0  2e-13
R_S0_45|4|B _S0_45|A4 _S0_45|4|MID_SHUNT  2.7439617672
L_S0_45|4|RB _S0_45|4|MID_SHUNT 0  1.550338398468e-12
B_S0_45|T|1 _S0_45|T1 _S0_45|T|MID_SERIES JJMIT AREA=2.5
L_S0_45|T|P _S0_45|T|MID_SERIES 0  2e-13
R_S0_45|T|B _S0_45|T1 _S0_45|T|MID_SHUNT  2.7439617672
L_S0_45|T|RB _S0_45|T|MID_SHUNT 0  1.550338398468e-12
B_S0_45|45|1 _S0_45|T2 _S0_45|A4 JJMIT AREA=1.7857142857142858
R_S0_45|45|B _S0_45|T2 _S0_45|45|MID_SHUNT  3.84154647408
L_S0_45|45|RB _S0_45|45|MID_SHUNT _S0_45|A4  2.1704737578552e-12
B_S0_45|6|1 _S0_45|Q1 _S0_45|6|MID_SERIES JJMIT AREA=2.5
L_S0_45|6|P _S0_45|6|MID_SERIES 0  2e-13
R_S0_45|6|B _S0_45|Q1 _S0_45|6|MID_SHUNT  2.7439617672
L_S0_45|6|RB _S0_45|6|MID_SHUNT 0  1.550338398468e-12
L_S1_45|I_1|B _S1_45|A1 _S1_45|I_1|MID  2e-12
I_S1_45|I_1|B 0 _S1_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S1_45|I_3|B _S1_45|A3 _S1_45|I_3|MID  2e-12
I_S1_45|I_3|B 0 _S1_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S1_45|I_T|B _S1_45|T1 _S1_45|I_T|MID  2e-12
I_S1_45|I_T|B 0 _S1_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S1_45|I_6|B _S1_45|Q1 _S1_45|I_6|MID  2e-12
I_S1_45|I_6|B 0 _S1_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S1_45|1|1 _S1_45|A1 _S1_45|1|MID_SERIES JJMIT AREA=2.5
L_S1_45|1|P _S1_45|1|MID_SERIES 0  2e-13
R_S1_45|1|B _S1_45|A1 _S1_45|1|MID_SHUNT  2.7439617672
L_S1_45|1|RB _S1_45|1|MID_SHUNT 0  1.550338398468e-12
B_S1_45|23|1 _S1_45|A2 _S1_45|A3 JJMIT AREA=1.7857142857142858
R_S1_45|23|B _S1_45|A2 _S1_45|23|MID_SHUNT  3.84154647408
L_S1_45|23|RB _S1_45|23|MID_SHUNT _S1_45|A3  2.1704737578552e-12
B_S1_45|3|1 _S1_45|A3 _S1_45|3|MID_SERIES JJMIT AREA=2.5
L_S1_45|3|P _S1_45|3|MID_SERIES 0  2e-13
R_S1_45|3|B _S1_45|A3 _S1_45|3|MID_SHUNT  2.7439617672
L_S1_45|3|RB _S1_45|3|MID_SHUNT 0  1.550338398468e-12
B_S1_45|4|1 _S1_45|A4 _S1_45|4|MID_SERIES JJMIT AREA=2.5
L_S1_45|4|P _S1_45|4|MID_SERIES 0  2e-13
R_S1_45|4|B _S1_45|A4 _S1_45|4|MID_SHUNT  2.7439617672
L_S1_45|4|RB _S1_45|4|MID_SHUNT 0  1.550338398468e-12
B_S1_45|T|1 _S1_45|T1 _S1_45|T|MID_SERIES JJMIT AREA=2.5
L_S1_45|T|P _S1_45|T|MID_SERIES 0  2e-13
R_S1_45|T|B _S1_45|T1 _S1_45|T|MID_SHUNT  2.7439617672
L_S1_45|T|RB _S1_45|T|MID_SHUNT 0  1.550338398468e-12
B_S1_45|45|1 _S1_45|T2 _S1_45|A4 JJMIT AREA=1.7857142857142858
R_S1_45|45|B _S1_45|T2 _S1_45|45|MID_SHUNT  3.84154647408
L_S1_45|45|RB _S1_45|45|MID_SHUNT _S1_45|A4  2.1704737578552e-12
B_S1_45|6|1 _S1_45|Q1 _S1_45|6|MID_SERIES JJMIT AREA=2.5
L_S1_45|6|P _S1_45|6|MID_SERIES 0  2e-13
R_S1_45|6|B _S1_45|Q1 _S1_45|6|MID_SHUNT  2.7439617672
L_S1_45|6|RB _S1_45|6|MID_SHUNT 0  1.550338398468e-12
L_S2_45|I_1|B _S2_45|A1 _S2_45|I_1|MID  2e-12
I_S2_45|I_1|B 0 _S2_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S2_45|I_3|B _S2_45|A3 _S2_45|I_3|MID  2e-12
I_S2_45|I_3|B 0 _S2_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S2_45|I_T|B _S2_45|T1 _S2_45|I_T|MID  2e-12
I_S2_45|I_T|B 0 _S2_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S2_45|I_6|B _S2_45|Q1 _S2_45|I_6|MID  2e-12
I_S2_45|I_6|B 0 _S2_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S2_45|1|1 _S2_45|A1 _S2_45|1|MID_SERIES JJMIT AREA=2.5
L_S2_45|1|P _S2_45|1|MID_SERIES 0  2e-13
R_S2_45|1|B _S2_45|A1 _S2_45|1|MID_SHUNT  2.7439617672
L_S2_45|1|RB _S2_45|1|MID_SHUNT 0  1.550338398468e-12
B_S2_45|23|1 _S2_45|A2 _S2_45|A3 JJMIT AREA=1.7857142857142858
R_S2_45|23|B _S2_45|A2 _S2_45|23|MID_SHUNT  3.84154647408
L_S2_45|23|RB _S2_45|23|MID_SHUNT _S2_45|A3  2.1704737578552e-12
B_S2_45|3|1 _S2_45|A3 _S2_45|3|MID_SERIES JJMIT AREA=2.5
L_S2_45|3|P _S2_45|3|MID_SERIES 0  2e-13
R_S2_45|3|B _S2_45|A3 _S2_45|3|MID_SHUNT  2.7439617672
L_S2_45|3|RB _S2_45|3|MID_SHUNT 0  1.550338398468e-12
B_S2_45|4|1 _S2_45|A4 _S2_45|4|MID_SERIES JJMIT AREA=2.5
L_S2_45|4|P _S2_45|4|MID_SERIES 0  2e-13
R_S2_45|4|B _S2_45|A4 _S2_45|4|MID_SHUNT  2.7439617672
L_S2_45|4|RB _S2_45|4|MID_SHUNT 0  1.550338398468e-12
B_S2_45|T|1 _S2_45|T1 _S2_45|T|MID_SERIES JJMIT AREA=2.5
L_S2_45|T|P _S2_45|T|MID_SERIES 0  2e-13
R_S2_45|T|B _S2_45|T1 _S2_45|T|MID_SHUNT  2.7439617672
L_S2_45|T|RB _S2_45|T|MID_SHUNT 0  1.550338398468e-12
B_S2_45|45|1 _S2_45|T2 _S2_45|A4 JJMIT AREA=1.7857142857142858
R_S2_45|45|B _S2_45|T2 _S2_45|45|MID_SHUNT  3.84154647408
L_S2_45|45|RB _S2_45|45|MID_SHUNT _S2_45|A4  2.1704737578552e-12
B_S2_45|6|1 _S2_45|Q1 _S2_45|6|MID_SERIES JJMIT AREA=2.5
L_S2_45|6|P _S2_45|6|MID_SERIES 0  2e-13
R_S2_45|6|B _S2_45|Q1 _S2_45|6|MID_SHUNT  2.7439617672
L_S2_45|6|RB _S2_45|6|MID_SHUNT 0  1.550338398468e-12
L_S3_45|I_1|B _S3_45|A1 _S3_45|I_1|MID  2e-12
I_S3_45|I_1|B 0 _S3_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S3_45|I_3|B _S3_45|A3 _S3_45|I_3|MID  2e-12
I_S3_45|I_3|B 0 _S3_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S3_45|I_T|B _S3_45|T1 _S3_45|I_T|MID  2e-12
I_S3_45|I_T|B 0 _S3_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S3_45|I_6|B _S3_45|Q1 _S3_45|I_6|MID  2e-12
I_S3_45|I_6|B 0 _S3_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S3_45|1|1 _S3_45|A1 _S3_45|1|MID_SERIES JJMIT AREA=2.5
L_S3_45|1|P _S3_45|1|MID_SERIES 0  2e-13
R_S3_45|1|B _S3_45|A1 _S3_45|1|MID_SHUNT  2.7439617672
L_S3_45|1|RB _S3_45|1|MID_SHUNT 0  1.550338398468e-12
B_S3_45|23|1 _S3_45|A2 _S3_45|A3 JJMIT AREA=1.7857142857142858
R_S3_45|23|B _S3_45|A2 _S3_45|23|MID_SHUNT  3.84154647408
L_S3_45|23|RB _S3_45|23|MID_SHUNT _S3_45|A3  2.1704737578552e-12
B_S3_45|3|1 _S3_45|A3 _S3_45|3|MID_SERIES JJMIT AREA=2.5
L_S3_45|3|P _S3_45|3|MID_SERIES 0  2e-13
R_S3_45|3|B _S3_45|A3 _S3_45|3|MID_SHUNT  2.7439617672
L_S3_45|3|RB _S3_45|3|MID_SHUNT 0  1.550338398468e-12
B_S3_45|4|1 _S3_45|A4 _S3_45|4|MID_SERIES JJMIT AREA=2.5
L_S3_45|4|P _S3_45|4|MID_SERIES 0  2e-13
R_S3_45|4|B _S3_45|A4 _S3_45|4|MID_SHUNT  2.7439617672
L_S3_45|4|RB _S3_45|4|MID_SHUNT 0  1.550338398468e-12
B_S3_45|T|1 _S3_45|T1 _S3_45|T|MID_SERIES JJMIT AREA=2.5
L_S3_45|T|P _S3_45|T|MID_SERIES 0  2e-13
R_S3_45|T|B _S3_45|T1 _S3_45|T|MID_SHUNT  2.7439617672
L_S3_45|T|RB _S3_45|T|MID_SHUNT 0  1.550338398468e-12
B_S3_45|45|1 _S3_45|T2 _S3_45|A4 JJMIT AREA=1.7857142857142858
R_S3_45|45|B _S3_45|T2 _S3_45|45|MID_SHUNT  3.84154647408
L_S3_45|45|RB _S3_45|45|MID_SHUNT _S3_45|A4  2.1704737578552e-12
B_S3_45|6|1 _S3_45|Q1 _S3_45|6|MID_SERIES JJMIT AREA=2.5
L_S3_45|6|P _S3_45|6|MID_SERIES 0  2e-13
R_S3_45|6|B _S3_45|Q1 _S3_45|6|MID_SHUNT  2.7439617672
L_S3_45|6|RB _S3_45|6|MID_SHUNT 0  1.550338398468e-12
L_S4_45|I_1|B _S4_45|A1 _S4_45|I_1|MID  2e-12
I_S4_45|I_1|B 0 _S4_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S4_45|I_3|B _S4_45|A3 _S4_45|I_3|MID  2e-12
I_S4_45|I_3|B 0 _S4_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S4_45|I_T|B _S4_45|T1 _S4_45|I_T|MID  2e-12
I_S4_45|I_T|B 0 _S4_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S4_45|I_6|B _S4_45|Q1 _S4_45|I_6|MID  2e-12
I_S4_45|I_6|B 0 _S4_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S4_45|1|1 _S4_45|A1 _S4_45|1|MID_SERIES JJMIT AREA=2.5
L_S4_45|1|P _S4_45|1|MID_SERIES 0  2e-13
R_S4_45|1|B _S4_45|A1 _S4_45|1|MID_SHUNT  2.7439617672
L_S4_45|1|RB _S4_45|1|MID_SHUNT 0  1.550338398468e-12
B_S4_45|23|1 _S4_45|A2 _S4_45|A3 JJMIT AREA=1.7857142857142858
R_S4_45|23|B _S4_45|A2 _S4_45|23|MID_SHUNT  3.84154647408
L_S4_45|23|RB _S4_45|23|MID_SHUNT _S4_45|A3  2.1704737578552e-12
B_S4_45|3|1 _S4_45|A3 _S4_45|3|MID_SERIES JJMIT AREA=2.5
L_S4_45|3|P _S4_45|3|MID_SERIES 0  2e-13
R_S4_45|3|B _S4_45|A3 _S4_45|3|MID_SHUNT  2.7439617672
L_S4_45|3|RB _S4_45|3|MID_SHUNT 0  1.550338398468e-12
B_S4_45|4|1 _S4_45|A4 _S4_45|4|MID_SERIES JJMIT AREA=2.5
L_S4_45|4|P _S4_45|4|MID_SERIES 0  2e-13
R_S4_45|4|B _S4_45|A4 _S4_45|4|MID_SHUNT  2.7439617672
L_S4_45|4|RB _S4_45|4|MID_SHUNT 0  1.550338398468e-12
B_S4_45|T|1 _S4_45|T1 _S4_45|T|MID_SERIES JJMIT AREA=2.5
L_S4_45|T|P _S4_45|T|MID_SERIES 0  2e-13
R_S4_45|T|B _S4_45|T1 _S4_45|T|MID_SHUNT  2.7439617672
L_S4_45|T|RB _S4_45|T|MID_SHUNT 0  1.550338398468e-12
B_S4_45|45|1 _S4_45|T2 _S4_45|A4 JJMIT AREA=1.7857142857142858
R_S4_45|45|B _S4_45|T2 _S4_45|45|MID_SHUNT  3.84154647408
L_S4_45|45|RB _S4_45|45|MID_SHUNT _S4_45|A4  2.1704737578552e-12
B_S4_45|6|1 _S4_45|Q1 _S4_45|6|MID_SERIES JJMIT AREA=2.5
L_S4_45|6|P _S4_45|6|MID_SERIES 0  2e-13
R_S4_45|6|B _S4_45|Q1 _S4_45|6|MID_SHUNT  2.7439617672
L_S4_45|6|RB _S4_45|6|MID_SHUNT 0  1.550338398468e-12
L_S5_45|I_1|B _S5_45|A1 _S5_45|I_1|MID  2e-12
I_S5_45|I_1|B 0 _S5_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S5_45|I_3|B _S5_45|A3 _S5_45|I_3|MID  2e-12
I_S5_45|I_3|B 0 _S5_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S5_45|I_T|B _S5_45|T1 _S5_45|I_T|MID  2e-12
I_S5_45|I_T|B 0 _S5_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S5_45|I_6|B _S5_45|Q1 _S5_45|I_6|MID  2e-12
I_S5_45|I_6|B 0 _S5_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S5_45|1|1 _S5_45|A1 _S5_45|1|MID_SERIES JJMIT AREA=2.5
L_S5_45|1|P _S5_45|1|MID_SERIES 0  2e-13
R_S5_45|1|B _S5_45|A1 _S5_45|1|MID_SHUNT  2.7439617672
L_S5_45|1|RB _S5_45|1|MID_SHUNT 0  1.550338398468e-12
B_S5_45|23|1 _S5_45|A2 _S5_45|A3 JJMIT AREA=1.7857142857142858
R_S5_45|23|B _S5_45|A2 _S5_45|23|MID_SHUNT  3.84154647408
L_S5_45|23|RB _S5_45|23|MID_SHUNT _S5_45|A3  2.1704737578552e-12
B_S5_45|3|1 _S5_45|A3 _S5_45|3|MID_SERIES JJMIT AREA=2.5
L_S5_45|3|P _S5_45|3|MID_SERIES 0  2e-13
R_S5_45|3|B _S5_45|A3 _S5_45|3|MID_SHUNT  2.7439617672
L_S5_45|3|RB _S5_45|3|MID_SHUNT 0  1.550338398468e-12
B_S5_45|4|1 _S5_45|A4 _S5_45|4|MID_SERIES JJMIT AREA=2.5
L_S5_45|4|P _S5_45|4|MID_SERIES 0  2e-13
R_S5_45|4|B _S5_45|A4 _S5_45|4|MID_SHUNT  2.7439617672
L_S5_45|4|RB _S5_45|4|MID_SHUNT 0  1.550338398468e-12
B_S5_45|T|1 _S5_45|T1 _S5_45|T|MID_SERIES JJMIT AREA=2.5
L_S5_45|T|P _S5_45|T|MID_SERIES 0  2e-13
R_S5_45|T|B _S5_45|T1 _S5_45|T|MID_SHUNT  2.7439617672
L_S5_45|T|RB _S5_45|T|MID_SHUNT 0  1.550338398468e-12
B_S5_45|45|1 _S5_45|T2 _S5_45|A4 JJMIT AREA=1.7857142857142858
R_S5_45|45|B _S5_45|T2 _S5_45|45|MID_SHUNT  3.84154647408
L_S5_45|45|RB _S5_45|45|MID_SHUNT _S5_45|A4  2.1704737578552e-12
B_S5_45|6|1 _S5_45|Q1 _S5_45|6|MID_SERIES JJMIT AREA=2.5
L_S5_45|6|P _S5_45|6|MID_SERIES 0  2e-13
R_S5_45|6|B _S5_45|Q1 _S5_45|6|MID_SHUNT  2.7439617672
L_S5_45|6|RB _S5_45|6|MID_SHUNT 0  1.550338398468e-12
L_S6_45|I_1|B _S6_45|A1 _S6_45|I_1|MID  2e-12
I_S6_45|I_1|B 0 _S6_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S6_45|I_3|B _S6_45|A3 _S6_45|I_3|MID  2e-12
I_S6_45|I_3|B 0 _S6_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S6_45|I_T|B _S6_45|T1 _S6_45|I_T|MID  2e-12
I_S6_45|I_T|B 0 _S6_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S6_45|I_6|B _S6_45|Q1 _S6_45|I_6|MID  2e-12
I_S6_45|I_6|B 0 _S6_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S6_45|1|1 _S6_45|A1 _S6_45|1|MID_SERIES JJMIT AREA=2.5
L_S6_45|1|P _S6_45|1|MID_SERIES 0  2e-13
R_S6_45|1|B _S6_45|A1 _S6_45|1|MID_SHUNT  2.7439617672
L_S6_45|1|RB _S6_45|1|MID_SHUNT 0  1.550338398468e-12
B_S6_45|23|1 _S6_45|A2 _S6_45|A3 JJMIT AREA=1.7857142857142858
R_S6_45|23|B _S6_45|A2 _S6_45|23|MID_SHUNT  3.84154647408
L_S6_45|23|RB _S6_45|23|MID_SHUNT _S6_45|A3  2.1704737578552e-12
B_S6_45|3|1 _S6_45|A3 _S6_45|3|MID_SERIES JJMIT AREA=2.5
L_S6_45|3|P _S6_45|3|MID_SERIES 0  2e-13
R_S6_45|3|B _S6_45|A3 _S6_45|3|MID_SHUNT  2.7439617672
L_S6_45|3|RB _S6_45|3|MID_SHUNT 0  1.550338398468e-12
B_S6_45|4|1 _S6_45|A4 _S6_45|4|MID_SERIES JJMIT AREA=2.5
L_S6_45|4|P _S6_45|4|MID_SERIES 0  2e-13
R_S6_45|4|B _S6_45|A4 _S6_45|4|MID_SHUNT  2.7439617672
L_S6_45|4|RB _S6_45|4|MID_SHUNT 0  1.550338398468e-12
B_S6_45|T|1 _S6_45|T1 _S6_45|T|MID_SERIES JJMIT AREA=2.5
L_S6_45|T|P _S6_45|T|MID_SERIES 0  2e-13
R_S6_45|T|B _S6_45|T1 _S6_45|T|MID_SHUNT  2.7439617672
L_S6_45|T|RB _S6_45|T|MID_SHUNT 0  1.550338398468e-12
B_S6_45|45|1 _S6_45|T2 _S6_45|A4 JJMIT AREA=1.7857142857142858
R_S6_45|45|B _S6_45|T2 _S6_45|45|MID_SHUNT  3.84154647408
L_S6_45|45|RB _S6_45|45|MID_SHUNT _S6_45|A4  2.1704737578552e-12
B_S6_45|6|1 _S6_45|Q1 _S6_45|6|MID_SERIES JJMIT AREA=2.5
L_S6_45|6|P _S6_45|6|MID_SERIES 0  2e-13
R_S6_45|6|B _S6_45|Q1 _S6_45|6|MID_SHUNT  2.7439617672
L_S6_45|6|RB _S6_45|6|MID_SHUNT 0  1.550338398468e-12
L_S7_45|I_A1|B _S7_45|A1 _S7_45|I_A1|MID  2e-12
I_S7_45|I_A1|B 0 _S7_45|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S7_45|I_A3|B _S7_45|A3 _S7_45|I_A3|MID  2e-12
I_S7_45|I_A3|B 0 _S7_45|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S7_45|I_B1|B _S7_45|B1 _S7_45|I_B1|MID  2e-12
I_S7_45|I_B1|B 0 _S7_45|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S7_45|I_B3|B _S7_45|B3 _S7_45|I_B3|MID  2e-12
I_S7_45|I_B3|B 0 _S7_45|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S7_45|I_Q1|B _S7_45|Q1 _S7_45|I_Q1|MID  2e-12
I_S7_45|I_Q1|B 0 _S7_45|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S7_45|A1|1 _S7_45|A1 _S7_45|A1|MID_SERIES JJMIT AREA=2.5
L_S7_45|A1|P _S7_45|A1|MID_SERIES 0  5e-13
R_S7_45|A1|B _S7_45|A1 _S7_45|A1|MID_SHUNT  2.7439617672
L_S7_45|A1|RB _S7_45|A1|MID_SHUNT 0  2.050338398468e-12
B_S7_45|A2|1 _S7_45|A2 _S7_45|A2|MID_SERIES JJMIT AREA=2.5
L_S7_45|A2|P _S7_45|A2|MID_SERIES 0  5e-13
R_S7_45|A2|B _S7_45|A2 _S7_45|A2|MID_SHUNT  2.7439617672
L_S7_45|A2|RB _S7_45|A2|MID_SHUNT 0  2.050338398468e-12
B_S7_45|A3|1 _S7_45|A2 _S7_45|A3|MID_SERIES JJMIT AREA=2.5
L_S7_45|A3|P _S7_45|A3|MID_SERIES _S7_45|A3  1.2e-12
R_S7_45|A3|B _S7_45|A2 _S7_45|A3|MID_SHUNT  2.7439617672
L_S7_45|A3|RB _S7_45|A3|MID_SHUNT _S7_45|A3  2.050338398468e-12
B_S7_45|B1|1 _S7_45|B1 _S7_45|B1|MID_SERIES JJMIT AREA=2.5
L_S7_45|B1|P _S7_45|B1|MID_SERIES 0  5e-13
R_S7_45|B1|B _S7_45|B1 _S7_45|B1|MID_SHUNT  2.7439617672
L_S7_45|B1|RB _S7_45|B1|MID_SHUNT 0  2.050338398468e-12
B_S7_45|B2|1 _S7_45|B2 _S7_45|B2|MID_SERIES JJMIT AREA=2.5
L_S7_45|B2|P _S7_45|B2|MID_SERIES 0  5e-13
R_S7_45|B2|B _S7_45|B2 _S7_45|B2|MID_SHUNT  2.7439617672
L_S7_45|B2|RB _S7_45|B2|MID_SHUNT 0  2.050338398468e-12
B_S7_45|B3|1 _S7_45|B2 _S7_45|B3|MID_SERIES JJMIT AREA=2.5
L_S7_45|B3|P _S7_45|B3|MID_SERIES _S7_45|B3  1.2e-12
R_S7_45|B3|B _S7_45|B2 _S7_45|B3|MID_SHUNT  2.7439617672
L_S7_45|B3|RB _S7_45|B3|MID_SHUNT _S7_45|B3  2.050338398468e-12
B_S7_45|T1|1 _S7_45|T1 _S7_45|T1|MID_SERIES JJMIT AREA=2.5
L_S7_45|T1|P _S7_45|T1|MID_SERIES 0  5e-13
R_S7_45|T1|B _S7_45|T1 _S7_45|T1|MID_SHUNT  2.7439617672
L_S7_45|T1|RB _S7_45|T1|MID_SHUNT 0  2.050338398468e-12
B_S7_45|T2|1 _S7_45|T2 _S7_45|ABTQ JJMIT AREA=2.0
R_S7_45|T2|B _S7_45|T2 _S7_45|T2|MID_SHUNT  3.429952209
L_S7_45|T2|RB _S7_45|T2|MID_SHUNT _S7_45|ABTQ  2.437922998085e-12
B_S7_45|AB|1 _S7_45|AB _S7_45|AB|MID_SERIES JJMIT AREA=1.5
L_S7_45|AB|P _S7_45|AB|MID_SERIES _S7_45|ABTQ  1.2e-12
R_S7_45|AB|B _S7_45|AB _S7_45|AB|MID_SHUNT  4.573269612
L_S7_45|AB|RB _S7_45|AB|MID_SHUNT _S7_45|ABTQ  3.08389733078e-12
B_S7_45|ABTQ|1 _S7_45|ABTQ _S7_45|ABTQ|MID_SERIES JJMIT AREA=1.875
L_S7_45|ABTQ|P _S7_45|ABTQ|MID_SERIES 0  5e-13
R_S7_45|ABTQ|B _S7_45|ABTQ _S7_45|ABTQ|MID_SHUNT  3.6586156896
L_S7_45|ABTQ|RB _S7_45|ABTQ|MID_SHUNT 0  2.567117864624e-12
B_S7_45|Q1|1 _S7_45|Q1 _S7_45|Q1|MID_SERIES JJMIT AREA=2.5
L_S7_45|Q1|P _S7_45|Q1|MID_SERIES 0  5e-13
R_S7_45|Q1|B _S7_45|Q1 _S7_45|Q1|MID_SHUNT  2.7439617672
L_S7_45|Q1|RB _S7_45|Q1|MID_SHUNT 0  2.050338398468e-12
L_S8_45|I_1|B _S8_45|A1 _S8_45|I_1|MID  2e-12
I_S8_45|I_1|B 0 _S8_45|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S8_45|I_3|B _S8_45|A3 _S8_45|I_3|MID  2e-12
I_S8_45|I_3|B 0 _S8_45|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S8_45|I_T|B _S8_45|T1 _S8_45|I_T|MID  2e-12
I_S8_45|I_T|B 0 _S8_45|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S8_45|I_6|B _S8_45|Q1 _S8_45|I_6|MID  2e-12
I_S8_45|I_6|B 0 _S8_45|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S8_45|1|1 _S8_45|A1 _S8_45|1|MID_SERIES JJMIT AREA=2.5
L_S8_45|1|P _S8_45|1|MID_SERIES 0  2e-13
R_S8_45|1|B _S8_45|A1 _S8_45|1|MID_SHUNT  2.7439617672
L_S8_45|1|RB _S8_45|1|MID_SHUNT 0  1.550338398468e-12
B_S8_45|23|1 _S8_45|A2 _S8_45|A3 JJMIT AREA=1.7857142857142858
R_S8_45|23|B _S8_45|A2 _S8_45|23|MID_SHUNT  3.84154647408
L_S8_45|23|RB _S8_45|23|MID_SHUNT _S8_45|A3  2.1704737578552e-12
B_S8_45|3|1 _S8_45|A3 _S8_45|3|MID_SERIES JJMIT AREA=2.5
L_S8_45|3|P _S8_45|3|MID_SERIES 0  2e-13
R_S8_45|3|B _S8_45|A3 _S8_45|3|MID_SHUNT  2.7439617672
L_S8_45|3|RB _S8_45|3|MID_SHUNT 0  1.550338398468e-12
B_S8_45|4|1 _S8_45|A4 _S8_45|4|MID_SERIES JJMIT AREA=2.5
L_S8_45|4|P _S8_45|4|MID_SERIES 0  2e-13
R_S8_45|4|B _S8_45|A4 _S8_45|4|MID_SHUNT  2.7439617672
L_S8_45|4|RB _S8_45|4|MID_SHUNT 0  1.550338398468e-12
B_S8_45|T|1 _S8_45|T1 _S8_45|T|MID_SERIES JJMIT AREA=2.5
L_S8_45|T|P _S8_45|T|MID_SERIES 0  2e-13
R_S8_45|T|B _S8_45|T1 _S8_45|T|MID_SHUNT  2.7439617672
L_S8_45|T|RB _S8_45|T|MID_SHUNT 0  1.550338398468e-12
B_S8_45|45|1 _S8_45|T2 _S8_45|A4 JJMIT AREA=1.7857142857142858
R_S8_45|45|B _S8_45|T2 _S8_45|45|MID_SHUNT  3.84154647408
L_S8_45|45|RB _S8_45|45|MID_SHUNT _S8_45|A4  2.1704737578552e-12
B_S8_45|6|1 _S8_45|Q1 _S8_45|6|MID_SERIES JJMIT AREA=2.5
L_S8_45|6|P _S8_45|6|MID_SERIES 0  2e-13
R_S8_45|6|B _S8_45|Q1 _S8_45|6|MID_SHUNT  2.7439617672
L_S8_45|6|RB _S8_45|6|MID_SHUNT 0  1.550338398468e-12
B_PTL_S0_5|_TX|1 _PTL_S0_5|_TX|1 _PTL_S0_5|_TX|2 JJMIT AREA=2.5
B_PTL_S0_5|_TX|2 _PTL_S0_5|_TX|4 _PTL_S0_5|_TX|5 JJMIT AREA=2.5
I_PTL_S0_5|_TX|B1 0 _PTL_S0_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S0_5|_TX|B2 0 _PTL_S0_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S0_5|_TX|B1 _PTL_S0_5|_TX|1 _PTL_S0_5|_TX|3  1.684e-12
L_PTL_S0_5|_TX|B2 _PTL_S0_5|_TX|4 _PTL_S0_5|_TX|6  3.596e-12
L_PTL_S0_5|_TX|1 S0_5_TX _PTL_S0_5|_TX|1  2.063e-12
L_PTL_S0_5|_TX|2 _PTL_S0_5|_TX|1 _PTL_S0_5|_TX|4  4.123e-12
L_PTL_S0_5|_TX|3 _PTL_S0_5|_TX|4 _PTL_S0_5|_TX|7  2.193e-12
R_PTL_S0_5|_TX|D _PTL_S0_5|_TX|7 _PTL_S0_5|A_PTL  1.36
L_PTL_S0_5|_TX|P1 _PTL_S0_5|_TX|2 0  5.254e-13
L_PTL_S0_5|_TX|P2 _PTL_S0_5|_TX|5 0  5.141e-13
R_PTL_S0_5|_TX|B1 _PTL_S0_5|_TX|1 _PTL_S0_5|_TX|101  2.7439617672
R_PTL_S0_5|_TX|B2 _PTL_S0_5|_TX|4 _PTL_S0_5|_TX|104  2.7439617672
L_PTL_S0_5|_TX|RB1 _PTL_S0_5|_TX|101 0  1.550338398468e-12
L_PTL_S0_5|_TX|RB2 _PTL_S0_5|_TX|104 0  1.550338398468e-12
B_PTL_S0_5|_RX|1 _PTL_S0_5|_RX|1 _PTL_S0_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S0_5|_RX|2 _PTL_S0_5|_RX|4 _PTL_S0_5|_RX|5 JJMIT AREA=2.0
B_PTL_S0_5|_RX|3 _PTL_S0_5|_RX|7 _PTL_S0_5|_RX|8 JJMIT AREA=2.5
I_PTL_S0_5|_RX|B1 0 _PTL_S0_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S0_5|_RX|B1 _PTL_S0_5|_RX|1 _PTL_S0_5|_RX|3  2.777e-12
I_PTL_S0_5|_RX|B2 0 _PTL_S0_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S0_5|_RX|B2 _PTL_S0_5|_RX|4 _PTL_S0_5|_RX|6  2.685e-12
I_PTL_S0_5|_RX|B3 0 _PTL_S0_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S0_5|_RX|B3 _PTL_S0_5|_RX|7 _PTL_S0_5|_RX|9  2.764e-12
L_PTL_S0_5|_RX|1 _PTL_S0_5|A_PTL _PTL_S0_5|_RX|1  1.346e-12
L_PTL_S0_5|_RX|2 _PTL_S0_5|_RX|1 _PTL_S0_5|_RX|4  6.348e-12
L_PTL_S0_5|_RX|3 _PTL_S0_5|_RX|4 _PTL_S0_5|_RX|7  5.197e-12
L_PTL_S0_5|_RX|4 _PTL_S0_5|_RX|7 S0_5  2.058e-12
L_PTL_S0_5|_RX|P1 _PTL_S0_5|_RX|2 0  4.795e-13
L_PTL_S0_5|_RX|P2 _PTL_S0_5|_RX|5 0  5.431e-13
L_PTL_S0_5|_RX|P3 _PTL_S0_5|_RX|8 0  5.339e-13
R_PTL_S0_5|_RX|B1 _PTL_S0_5|_RX|1 _PTL_S0_5|_RX|101  4.225701121488
R_PTL_S0_5|_RX|B2 _PTL_S0_5|_RX|4 _PTL_S0_5|_RX|104  3.429952209
R_PTL_S0_5|_RX|B3 _PTL_S0_5|_RX|7 _PTL_S0_5|_RX|107  2.7439617672
L_PTL_S0_5|_RX|RB1 _PTL_S0_5|_RX|101 0  2.38752113364072e-12
L_PTL_S0_5|_RX|RB2 _PTL_S0_5|_RX|104 0  1.937922998085e-12
L_PTL_S0_5|_RX|RB3 _PTL_S0_5|_RX|107 0  1.550338398468e-12
B_PTL_S1_5|_TX|1 _PTL_S1_5|_TX|1 _PTL_S1_5|_TX|2 JJMIT AREA=2.5
B_PTL_S1_5|_TX|2 _PTL_S1_5|_TX|4 _PTL_S1_5|_TX|5 JJMIT AREA=2.5
I_PTL_S1_5|_TX|B1 0 _PTL_S1_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S1_5|_TX|B2 0 _PTL_S1_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S1_5|_TX|B1 _PTL_S1_5|_TX|1 _PTL_S1_5|_TX|3  1.684e-12
L_PTL_S1_5|_TX|B2 _PTL_S1_5|_TX|4 _PTL_S1_5|_TX|6  3.596e-12
L_PTL_S1_5|_TX|1 S1_5_TX _PTL_S1_5|_TX|1  2.063e-12
L_PTL_S1_5|_TX|2 _PTL_S1_5|_TX|1 _PTL_S1_5|_TX|4  4.123e-12
L_PTL_S1_5|_TX|3 _PTL_S1_5|_TX|4 _PTL_S1_5|_TX|7  2.193e-12
R_PTL_S1_5|_TX|D _PTL_S1_5|_TX|7 _PTL_S1_5|A_PTL  1.36
L_PTL_S1_5|_TX|P1 _PTL_S1_5|_TX|2 0  5.254e-13
L_PTL_S1_5|_TX|P2 _PTL_S1_5|_TX|5 0  5.141e-13
R_PTL_S1_5|_TX|B1 _PTL_S1_5|_TX|1 _PTL_S1_5|_TX|101  2.7439617672
R_PTL_S1_5|_TX|B2 _PTL_S1_5|_TX|4 _PTL_S1_5|_TX|104  2.7439617672
L_PTL_S1_5|_TX|RB1 _PTL_S1_5|_TX|101 0  1.550338398468e-12
L_PTL_S1_5|_TX|RB2 _PTL_S1_5|_TX|104 0  1.550338398468e-12
B_PTL_S1_5|_RX|1 _PTL_S1_5|_RX|1 _PTL_S1_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S1_5|_RX|2 _PTL_S1_5|_RX|4 _PTL_S1_5|_RX|5 JJMIT AREA=2.0
B_PTL_S1_5|_RX|3 _PTL_S1_5|_RX|7 _PTL_S1_5|_RX|8 JJMIT AREA=2.5
I_PTL_S1_5|_RX|B1 0 _PTL_S1_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S1_5|_RX|B1 _PTL_S1_5|_RX|1 _PTL_S1_5|_RX|3  2.777e-12
I_PTL_S1_5|_RX|B2 0 _PTL_S1_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S1_5|_RX|B2 _PTL_S1_5|_RX|4 _PTL_S1_5|_RX|6  2.685e-12
I_PTL_S1_5|_RX|B3 0 _PTL_S1_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S1_5|_RX|B3 _PTL_S1_5|_RX|7 _PTL_S1_5|_RX|9  2.764e-12
L_PTL_S1_5|_RX|1 _PTL_S1_5|A_PTL _PTL_S1_5|_RX|1  1.346e-12
L_PTL_S1_5|_RX|2 _PTL_S1_5|_RX|1 _PTL_S1_5|_RX|4  6.348e-12
L_PTL_S1_5|_RX|3 _PTL_S1_5|_RX|4 _PTL_S1_5|_RX|7  5.197e-12
L_PTL_S1_5|_RX|4 _PTL_S1_5|_RX|7 S1_5  2.058e-12
L_PTL_S1_5|_RX|P1 _PTL_S1_5|_RX|2 0  4.795e-13
L_PTL_S1_5|_RX|P2 _PTL_S1_5|_RX|5 0  5.431e-13
L_PTL_S1_5|_RX|P3 _PTL_S1_5|_RX|8 0  5.339e-13
R_PTL_S1_5|_RX|B1 _PTL_S1_5|_RX|1 _PTL_S1_5|_RX|101  4.225701121488
R_PTL_S1_5|_RX|B2 _PTL_S1_5|_RX|4 _PTL_S1_5|_RX|104  3.429952209
R_PTL_S1_5|_RX|B3 _PTL_S1_5|_RX|7 _PTL_S1_5|_RX|107  2.7439617672
L_PTL_S1_5|_RX|RB1 _PTL_S1_5|_RX|101 0  2.38752113364072e-12
L_PTL_S1_5|_RX|RB2 _PTL_S1_5|_RX|104 0  1.937922998085e-12
L_PTL_S1_5|_RX|RB3 _PTL_S1_5|_RX|107 0  1.550338398468e-12
B_PTL_S2_5|_TX|1 _PTL_S2_5|_TX|1 _PTL_S2_5|_TX|2 JJMIT AREA=2.5
B_PTL_S2_5|_TX|2 _PTL_S2_5|_TX|4 _PTL_S2_5|_TX|5 JJMIT AREA=2.5
I_PTL_S2_5|_TX|B1 0 _PTL_S2_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S2_5|_TX|B2 0 _PTL_S2_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S2_5|_TX|B1 _PTL_S2_5|_TX|1 _PTL_S2_5|_TX|3  1.684e-12
L_PTL_S2_5|_TX|B2 _PTL_S2_5|_TX|4 _PTL_S2_5|_TX|6  3.596e-12
L_PTL_S2_5|_TX|1 S2_5_TX _PTL_S2_5|_TX|1  2.063e-12
L_PTL_S2_5|_TX|2 _PTL_S2_5|_TX|1 _PTL_S2_5|_TX|4  4.123e-12
L_PTL_S2_5|_TX|3 _PTL_S2_5|_TX|4 _PTL_S2_5|_TX|7  2.193e-12
R_PTL_S2_5|_TX|D _PTL_S2_5|_TX|7 _PTL_S2_5|A_PTL  1.36
L_PTL_S2_5|_TX|P1 _PTL_S2_5|_TX|2 0  5.254e-13
L_PTL_S2_5|_TX|P2 _PTL_S2_5|_TX|5 0  5.141e-13
R_PTL_S2_5|_TX|B1 _PTL_S2_5|_TX|1 _PTL_S2_5|_TX|101  2.7439617672
R_PTL_S2_5|_TX|B2 _PTL_S2_5|_TX|4 _PTL_S2_5|_TX|104  2.7439617672
L_PTL_S2_5|_TX|RB1 _PTL_S2_5|_TX|101 0  1.550338398468e-12
L_PTL_S2_5|_TX|RB2 _PTL_S2_5|_TX|104 0  1.550338398468e-12
B_PTL_S2_5|_RX|1 _PTL_S2_5|_RX|1 _PTL_S2_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S2_5|_RX|2 _PTL_S2_5|_RX|4 _PTL_S2_5|_RX|5 JJMIT AREA=2.0
B_PTL_S2_5|_RX|3 _PTL_S2_5|_RX|7 _PTL_S2_5|_RX|8 JJMIT AREA=2.5
I_PTL_S2_5|_RX|B1 0 _PTL_S2_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S2_5|_RX|B1 _PTL_S2_5|_RX|1 _PTL_S2_5|_RX|3  2.777e-12
I_PTL_S2_5|_RX|B2 0 _PTL_S2_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S2_5|_RX|B2 _PTL_S2_5|_RX|4 _PTL_S2_5|_RX|6  2.685e-12
I_PTL_S2_5|_RX|B3 0 _PTL_S2_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S2_5|_RX|B3 _PTL_S2_5|_RX|7 _PTL_S2_5|_RX|9  2.764e-12
L_PTL_S2_5|_RX|1 _PTL_S2_5|A_PTL _PTL_S2_5|_RX|1  1.346e-12
L_PTL_S2_5|_RX|2 _PTL_S2_5|_RX|1 _PTL_S2_5|_RX|4  6.348e-12
L_PTL_S2_5|_RX|3 _PTL_S2_5|_RX|4 _PTL_S2_5|_RX|7  5.197e-12
L_PTL_S2_5|_RX|4 _PTL_S2_5|_RX|7 S2_5  2.058e-12
L_PTL_S2_5|_RX|P1 _PTL_S2_5|_RX|2 0  4.795e-13
L_PTL_S2_5|_RX|P2 _PTL_S2_5|_RX|5 0  5.431e-13
L_PTL_S2_5|_RX|P3 _PTL_S2_5|_RX|8 0  5.339e-13
R_PTL_S2_5|_RX|B1 _PTL_S2_5|_RX|1 _PTL_S2_5|_RX|101  4.225701121488
R_PTL_S2_5|_RX|B2 _PTL_S2_5|_RX|4 _PTL_S2_5|_RX|104  3.429952209
R_PTL_S2_5|_RX|B3 _PTL_S2_5|_RX|7 _PTL_S2_5|_RX|107  2.7439617672
L_PTL_S2_5|_RX|RB1 _PTL_S2_5|_RX|101 0  2.38752113364072e-12
L_PTL_S2_5|_RX|RB2 _PTL_S2_5|_RX|104 0  1.937922998085e-12
L_PTL_S2_5|_RX|RB3 _PTL_S2_5|_RX|107 0  1.550338398468e-12
B_PTL_S3_5|_TX|1 _PTL_S3_5|_TX|1 _PTL_S3_5|_TX|2 JJMIT AREA=2.5
B_PTL_S3_5|_TX|2 _PTL_S3_5|_TX|4 _PTL_S3_5|_TX|5 JJMIT AREA=2.5
I_PTL_S3_5|_TX|B1 0 _PTL_S3_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S3_5|_TX|B2 0 _PTL_S3_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S3_5|_TX|B1 _PTL_S3_5|_TX|1 _PTL_S3_5|_TX|3  1.684e-12
L_PTL_S3_5|_TX|B2 _PTL_S3_5|_TX|4 _PTL_S3_5|_TX|6  3.596e-12
L_PTL_S3_5|_TX|1 S3_5_TX _PTL_S3_5|_TX|1  2.063e-12
L_PTL_S3_5|_TX|2 _PTL_S3_5|_TX|1 _PTL_S3_5|_TX|4  4.123e-12
L_PTL_S3_5|_TX|3 _PTL_S3_5|_TX|4 _PTL_S3_5|_TX|7  2.193e-12
R_PTL_S3_5|_TX|D _PTL_S3_5|_TX|7 _PTL_S3_5|A_PTL  1.36
L_PTL_S3_5|_TX|P1 _PTL_S3_5|_TX|2 0  5.254e-13
L_PTL_S3_5|_TX|P2 _PTL_S3_5|_TX|5 0  5.141e-13
R_PTL_S3_5|_TX|B1 _PTL_S3_5|_TX|1 _PTL_S3_5|_TX|101  2.7439617672
R_PTL_S3_5|_TX|B2 _PTL_S3_5|_TX|4 _PTL_S3_5|_TX|104  2.7439617672
L_PTL_S3_5|_TX|RB1 _PTL_S3_5|_TX|101 0  1.550338398468e-12
L_PTL_S3_5|_TX|RB2 _PTL_S3_5|_TX|104 0  1.550338398468e-12
B_PTL_S3_5|_RX|1 _PTL_S3_5|_RX|1 _PTL_S3_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S3_5|_RX|2 _PTL_S3_5|_RX|4 _PTL_S3_5|_RX|5 JJMIT AREA=2.0
B_PTL_S3_5|_RX|3 _PTL_S3_5|_RX|7 _PTL_S3_5|_RX|8 JJMIT AREA=2.5
I_PTL_S3_5|_RX|B1 0 _PTL_S3_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S3_5|_RX|B1 _PTL_S3_5|_RX|1 _PTL_S3_5|_RX|3  2.777e-12
I_PTL_S3_5|_RX|B2 0 _PTL_S3_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S3_5|_RX|B2 _PTL_S3_5|_RX|4 _PTL_S3_5|_RX|6  2.685e-12
I_PTL_S3_5|_RX|B3 0 _PTL_S3_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S3_5|_RX|B3 _PTL_S3_5|_RX|7 _PTL_S3_5|_RX|9  2.764e-12
L_PTL_S3_5|_RX|1 _PTL_S3_5|A_PTL _PTL_S3_5|_RX|1  1.346e-12
L_PTL_S3_5|_RX|2 _PTL_S3_5|_RX|1 _PTL_S3_5|_RX|4  6.348e-12
L_PTL_S3_5|_RX|3 _PTL_S3_5|_RX|4 _PTL_S3_5|_RX|7  5.197e-12
L_PTL_S3_5|_RX|4 _PTL_S3_5|_RX|7 S3_5  2.058e-12
L_PTL_S3_5|_RX|P1 _PTL_S3_5|_RX|2 0  4.795e-13
L_PTL_S3_5|_RX|P2 _PTL_S3_5|_RX|5 0  5.431e-13
L_PTL_S3_5|_RX|P3 _PTL_S3_5|_RX|8 0  5.339e-13
R_PTL_S3_5|_RX|B1 _PTL_S3_5|_RX|1 _PTL_S3_5|_RX|101  4.225701121488
R_PTL_S3_5|_RX|B2 _PTL_S3_5|_RX|4 _PTL_S3_5|_RX|104  3.429952209
R_PTL_S3_5|_RX|B3 _PTL_S3_5|_RX|7 _PTL_S3_5|_RX|107  2.7439617672
L_PTL_S3_5|_RX|RB1 _PTL_S3_5|_RX|101 0  2.38752113364072e-12
L_PTL_S3_5|_RX|RB2 _PTL_S3_5|_RX|104 0  1.937922998085e-12
L_PTL_S3_5|_RX|RB3 _PTL_S3_5|_RX|107 0  1.550338398468e-12
B_PTL_S4_5|_TX|1 _PTL_S4_5|_TX|1 _PTL_S4_5|_TX|2 JJMIT AREA=2.5
B_PTL_S4_5|_TX|2 _PTL_S4_5|_TX|4 _PTL_S4_5|_TX|5 JJMIT AREA=2.5
I_PTL_S4_5|_TX|B1 0 _PTL_S4_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S4_5|_TX|B2 0 _PTL_S4_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S4_5|_TX|B1 _PTL_S4_5|_TX|1 _PTL_S4_5|_TX|3  1.684e-12
L_PTL_S4_5|_TX|B2 _PTL_S4_5|_TX|4 _PTL_S4_5|_TX|6  3.596e-12
L_PTL_S4_5|_TX|1 S4_5_TX _PTL_S4_5|_TX|1  2.063e-12
L_PTL_S4_5|_TX|2 _PTL_S4_5|_TX|1 _PTL_S4_5|_TX|4  4.123e-12
L_PTL_S4_5|_TX|3 _PTL_S4_5|_TX|4 _PTL_S4_5|_TX|7  2.193e-12
R_PTL_S4_5|_TX|D _PTL_S4_5|_TX|7 _PTL_S4_5|A_PTL  1.36
L_PTL_S4_5|_TX|P1 _PTL_S4_5|_TX|2 0  5.254e-13
L_PTL_S4_5|_TX|P2 _PTL_S4_5|_TX|5 0  5.141e-13
R_PTL_S4_5|_TX|B1 _PTL_S4_5|_TX|1 _PTL_S4_5|_TX|101  2.7439617672
R_PTL_S4_5|_TX|B2 _PTL_S4_5|_TX|4 _PTL_S4_5|_TX|104  2.7439617672
L_PTL_S4_5|_TX|RB1 _PTL_S4_5|_TX|101 0  1.550338398468e-12
L_PTL_S4_5|_TX|RB2 _PTL_S4_5|_TX|104 0  1.550338398468e-12
B_PTL_S4_5|_RX|1 _PTL_S4_5|_RX|1 _PTL_S4_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S4_5|_RX|2 _PTL_S4_5|_RX|4 _PTL_S4_5|_RX|5 JJMIT AREA=2.0
B_PTL_S4_5|_RX|3 _PTL_S4_5|_RX|7 _PTL_S4_5|_RX|8 JJMIT AREA=2.5
I_PTL_S4_5|_RX|B1 0 _PTL_S4_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S4_5|_RX|B1 _PTL_S4_5|_RX|1 _PTL_S4_5|_RX|3  2.777e-12
I_PTL_S4_5|_RX|B2 0 _PTL_S4_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S4_5|_RX|B2 _PTL_S4_5|_RX|4 _PTL_S4_5|_RX|6  2.685e-12
I_PTL_S4_5|_RX|B3 0 _PTL_S4_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S4_5|_RX|B3 _PTL_S4_5|_RX|7 _PTL_S4_5|_RX|9  2.764e-12
L_PTL_S4_5|_RX|1 _PTL_S4_5|A_PTL _PTL_S4_5|_RX|1  1.346e-12
L_PTL_S4_5|_RX|2 _PTL_S4_5|_RX|1 _PTL_S4_5|_RX|4  6.348e-12
L_PTL_S4_5|_RX|3 _PTL_S4_5|_RX|4 _PTL_S4_5|_RX|7  5.197e-12
L_PTL_S4_5|_RX|4 _PTL_S4_5|_RX|7 S4_5  2.058e-12
L_PTL_S4_5|_RX|P1 _PTL_S4_5|_RX|2 0  4.795e-13
L_PTL_S4_5|_RX|P2 _PTL_S4_5|_RX|5 0  5.431e-13
L_PTL_S4_5|_RX|P3 _PTL_S4_5|_RX|8 0  5.339e-13
R_PTL_S4_5|_RX|B1 _PTL_S4_5|_RX|1 _PTL_S4_5|_RX|101  4.225701121488
R_PTL_S4_5|_RX|B2 _PTL_S4_5|_RX|4 _PTL_S4_5|_RX|104  3.429952209
R_PTL_S4_5|_RX|B3 _PTL_S4_5|_RX|7 _PTL_S4_5|_RX|107  2.7439617672
L_PTL_S4_5|_RX|RB1 _PTL_S4_5|_RX|101 0  2.38752113364072e-12
L_PTL_S4_5|_RX|RB2 _PTL_S4_5|_RX|104 0  1.937922998085e-12
L_PTL_S4_5|_RX|RB3 _PTL_S4_5|_RX|107 0  1.550338398468e-12
B_PTL_S5_5|_TX|1 _PTL_S5_5|_TX|1 _PTL_S5_5|_TX|2 JJMIT AREA=2.5
B_PTL_S5_5|_TX|2 _PTL_S5_5|_TX|4 _PTL_S5_5|_TX|5 JJMIT AREA=2.5
I_PTL_S5_5|_TX|B1 0 _PTL_S5_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S5_5|_TX|B2 0 _PTL_S5_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S5_5|_TX|B1 _PTL_S5_5|_TX|1 _PTL_S5_5|_TX|3  1.684e-12
L_PTL_S5_5|_TX|B2 _PTL_S5_5|_TX|4 _PTL_S5_5|_TX|6  3.596e-12
L_PTL_S5_5|_TX|1 S5_5_TX _PTL_S5_5|_TX|1  2.063e-12
L_PTL_S5_5|_TX|2 _PTL_S5_5|_TX|1 _PTL_S5_5|_TX|4  4.123e-12
L_PTL_S5_5|_TX|3 _PTL_S5_5|_TX|4 _PTL_S5_5|_TX|7  2.193e-12
R_PTL_S5_5|_TX|D _PTL_S5_5|_TX|7 _PTL_S5_5|A_PTL  1.36
L_PTL_S5_5|_TX|P1 _PTL_S5_5|_TX|2 0  5.254e-13
L_PTL_S5_5|_TX|P2 _PTL_S5_5|_TX|5 0  5.141e-13
R_PTL_S5_5|_TX|B1 _PTL_S5_5|_TX|1 _PTL_S5_5|_TX|101  2.7439617672
R_PTL_S5_5|_TX|B2 _PTL_S5_5|_TX|4 _PTL_S5_5|_TX|104  2.7439617672
L_PTL_S5_5|_TX|RB1 _PTL_S5_5|_TX|101 0  1.550338398468e-12
L_PTL_S5_5|_TX|RB2 _PTL_S5_5|_TX|104 0  1.550338398468e-12
B_PTL_S5_5|_RX|1 _PTL_S5_5|_RX|1 _PTL_S5_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S5_5|_RX|2 _PTL_S5_5|_RX|4 _PTL_S5_5|_RX|5 JJMIT AREA=2.0
B_PTL_S5_5|_RX|3 _PTL_S5_5|_RX|7 _PTL_S5_5|_RX|8 JJMIT AREA=2.5
I_PTL_S5_5|_RX|B1 0 _PTL_S5_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S5_5|_RX|B1 _PTL_S5_5|_RX|1 _PTL_S5_5|_RX|3  2.777e-12
I_PTL_S5_5|_RX|B2 0 _PTL_S5_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S5_5|_RX|B2 _PTL_S5_5|_RX|4 _PTL_S5_5|_RX|6  2.685e-12
I_PTL_S5_5|_RX|B3 0 _PTL_S5_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S5_5|_RX|B3 _PTL_S5_5|_RX|7 _PTL_S5_5|_RX|9  2.764e-12
L_PTL_S5_5|_RX|1 _PTL_S5_5|A_PTL _PTL_S5_5|_RX|1  1.346e-12
L_PTL_S5_5|_RX|2 _PTL_S5_5|_RX|1 _PTL_S5_5|_RX|4  6.348e-12
L_PTL_S5_5|_RX|3 _PTL_S5_5|_RX|4 _PTL_S5_5|_RX|7  5.197e-12
L_PTL_S5_5|_RX|4 _PTL_S5_5|_RX|7 S5_5  2.058e-12
L_PTL_S5_5|_RX|P1 _PTL_S5_5|_RX|2 0  4.795e-13
L_PTL_S5_5|_RX|P2 _PTL_S5_5|_RX|5 0  5.431e-13
L_PTL_S5_5|_RX|P3 _PTL_S5_5|_RX|8 0  5.339e-13
R_PTL_S5_5|_RX|B1 _PTL_S5_5|_RX|1 _PTL_S5_5|_RX|101  4.225701121488
R_PTL_S5_5|_RX|B2 _PTL_S5_5|_RX|4 _PTL_S5_5|_RX|104  3.429952209
R_PTL_S5_5|_RX|B3 _PTL_S5_5|_RX|7 _PTL_S5_5|_RX|107  2.7439617672
L_PTL_S5_5|_RX|RB1 _PTL_S5_5|_RX|101 0  2.38752113364072e-12
L_PTL_S5_5|_RX|RB2 _PTL_S5_5|_RX|104 0  1.937922998085e-12
L_PTL_S5_5|_RX|RB3 _PTL_S5_5|_RX|107 0  1.550338398468e-12
B_PTL_S6_5|_TX|1 _PTL_S6_5|_TX|1 _PTL_S6_5|_TX|2 JJMIT AREA=2.5
B_PTL_S6_5|_TX|2 _PTL_S6_5|_TX|4 _PTL_S6_5|_TX|5 JJMIT AREA=2.5
I_PTL_S6_5|_TX|B1 0 _PTL_S6_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S6_5|_TX|B2 0 _PTL_S6_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S6_5|_TX|B1 _PTL_S6_5|_TX|1 _PTL_S6_5|_TX|3  1.684e-12
L_PTL_S6_5|_TX|B2 _PTL_S6_5|_TX|4 _PTL_S6_5|_TX|6  3.596e-12
L_PTL_S6_5|_TX|1 S6_5_TX _PTL_S6_5|_TX|1  2.063e-12
L_PTL_S6_5|_TX|2 _PTL_S6_5|_TX|1 _PTL_S6_5|_TX|4  4.123e-12
L_PTL_S6_5|_TX|3 _PTL_S6_5|_TX|4 _PTL_S6_5|_TX|7  2.193e-12
R_PTL_S6_5|_TX|D _PTL_S6_5|_TX|7 _PTL_S6_5|A_PTL  1.36
L_PTL_S6_5|_TX|P1 _PTL_S6_5|_TX|2 0  5.254e-13
L_PTL_S6_5|_TX|P2 _PTL_S6_5|_TX|5 0  5.141e-13
R_PTL_S6_5|_TX|B1 _PTL_S6_5|_TX|1 _PTL_S6_5|_TX|101  2.7439617672
R_PTL_S6_5|_TX|B2 _PTL_S6_5|_TX|4 _PTL_S6_5|_TX|104  2.7439617672
L_PTL_S6_5|_TX|RB1 _PTL_S6_5|_TX|101 0  1.550338398468e-12
L_PTL_S6_5|_TX|RB2 _PTL_S6_5|_TX|104 0  1.550338398468e-12
B_PTL_S6_5|_RX|1 _PTL_S6_5|_RX|1 _PTL_S6_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S6_5|_RX|2 _PTL_S6_5|_RX|4 _PTL_S6_5|_RX|5 JJMIT AREA=2.0
B_PTL_S6_5|_RX|3 _PTL_S6_5|_RX|7 _PTL_S6_5|_RX|8 JJMIT AREA=2.5
I_PTL_S6_5|_RX|B1 0 _PTL_S6_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S6_5|_RX|B1 _PTL_S6_5|_RX|1 _PTL_S6_5|_RX|3  2.777e-12
I_PTL_S6_5|_RX|B2 0 _PTL_S6_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S6_5|_RX|B2 _PTL_S6_5|_RX|4 _PTL_S6_5|_RX|6  2.685e-12
I_PTL_S6_5|_RX|B3 0 _PTL_S6_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S6_5|_RX|B3 _PTL_S6_5|_RX|7 _PTL_S6_5|_RX|9  2.764e-12
L_PTL_S6_5|_RX|1 _PTL_S6_5|A_PTL _PTL_S6_5|_RX|1  1.346e-12
L_PTL_S6_5|_RX|2 _PTL_S6_5|_RX|1 _PTL_S6_5|_RX|4  6.348e-12
L_PTL_S6_5|_RX|3 _PTL_S6_5|_RX|4 _PTL_S6_5|_RX|7  5.197e-12
L_PTL_S6_5|_RX|4 _PTL_S6_5|_RX|7 S6_5  2.058e-12
L_PTL_S6_5|_RX|P1 _PTL_S6_5|_RX|2 0  4.795e-13
L_PTL_S6_5|_RX|P2 _PTL_S6_5|_RX|5 0  5.431e-13
L_PTL_S6_5|_RX|P3 _PTL_S6_5|_RX|8 0  5.339e-13
R_PTL_S6_5|_RX|B1 _PTL_S6_5|_RX|1 _PTL_S6_5|_RX|101  4.225701121488
R_PTL_S6_5|_RX|B2 _PTL_S6_5|_RX|4 _PTL_S6_5|_RX|104  3.429952209
R_PTL_S6_5|_RX|B3 _PTL_S6_5|_RX|7 _PTL_S6_5|_RX|107  2.7439617672
L_PTL_S6_5|_RX|RB1 _PTL_S6_5|_RX|101 0  2.38752113364072e-12
L_PTL_S6_5|_RX|RB2 _PTL_S6_5|_RX|104 0  1.937922998085e-12
L_PTL_S6_5|_RX|RB3 _PTL_S6_5|_RX|107 0  1.550338398468e-12
B_PTL_S7_5|_TX|1 _PTL_S7_5|_TX|1 _PTL_S7_5|_TX|2 JJMIT AREA=2.5
B_PTL_S7_5|_TX|2 _PTL_S7_5|_TX|4 _PTL_S7_5|_TX|5 JJMIT AREA=2.5
I_PTL_S7_5|_TX|B1 0 _PTL_S7_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S7_5|_TX|B2 0 _PTL_S7_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S7_5|_TX|B1 _PTL_S7_5|_TX|1 _PTL_S7_5|_TX|3  1.684e-12
L_PTL_S7_5|_TX|B2 _PTL_S7_5|_TX|4 _PTL_S7_5|_TX|6  3.596e-12
L_PTL_S7_5|_TX|1 S7_5_TX _PTL_S7_5|_TX|1  2.063e-12
L_PTL_S7_5|_TX|2 _PTL_S7_5|_TX|1 _PTL_S7_5|_TX|4  4.123e-12
L_PTL_S7_5|_TX|3 _PTL_S7_5|_TX|4 _PTL_S7_5|_TX|7  2.193e-12
R_PTL_S7_5|_TX|D _PTL_S7_5|_TX|7 _PTL_S7_5|A_PTL  1.36
L_PTL_S7_5|_TX|P1 _PTL_S7_5|_TX|2 0  5.254e-13
L_PTL_S7_5|_TX|P2 _PTL_S7_5|_TX|5 0  5.141e-13
R_PTL_S7_5|_TX|B1 _PTL_S7_5|_TX|1 _PTL_S7_5|_TX|101  2.7439617672
R_PTL_S7_5|_TX|B2 _PTL_S7_5|_TX|4 _PTL_S7_5|_TX|104  2.7439617672
L_PTL_S7_5|_TX|RB1 _PTL_S7_5|_TX|101 0  1.550338398468e-12
L_PTL_S7_5|_TX|RB2 _PTL_S7_5|_TX|104 0  1.550338398468e-12
B_PTL_S7_5|_RX|1 _PTL_S7_5|_RX|1 _PTL_S7_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S7_5|_RX|2 _PTL_S7_5|_RX|4 _PTL_S7_5|_RX|5 JJMIT AREA=2.0
B_PTL_S7_5|_RX|3 _PTL_S7_5|_RX|7 _PTL_S7_5|_RX|8 JJMIT AREA=2.5
I_PTL_S7_5|_RX|B1 0 _PTL_S7_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S7_5|_RX|B1 _PTL_S7_5|_RX|1 _PTL_S7_5|_RX|3  2.777e-12
I_PTL_S7_5|_RX|B2 0 _PTL_S7_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S7_5|_RX|B2 _PTL_S7_5|_RX|4 _PTL_S7_5|_RX|6  2.685e-12
I_PTL_S7_5|_RX|B3 0 _PTL_S7_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S7_5|_RX|B3 _PTL_S7_5|_RX|7 _PTL_S7_5|_RX|9  2.764e-12
L_PTL_S7_5|_RX|1 _PTL_S7_5|A_PTL _PTL_S7_5|_RX|1  1.346e-12
L_PTL_S7_5|_RX|2 _PTL_S7_5|_RX|1 _PTL_S7_5|_RX|4  6.348e-12
L_PTL_S7_5|_RX|3 _PTL_S7_5|_RX|4 _PTL_S7_5|_RX|7  5.197e-12
L_PTL_S7_5|_RX|4 _PTL_S7_5|_RX|7 S7_5  2.058e-12
L_PTL_S7_5|_RX|P1 _PTL_S7_5|_RX|2 0  4.795e-13
L_PTL_S7_5|_RX|P2 _PTL_S7_5|_RX|5 0  5.431e-13
L_PTL_S7_5|_RX|P3 _PTL_S7_5|_RX|8 0  5.339e-13
R_PTL_S7_5|_RX|B1 _PTL_S7_5|_RX|1 _PTL_S7_5|_RX|101  4.225701121488
R_PTL_S7_5|_RX|B2 _PTL_S7_5|_RX|4 _PTL_S7_5|_RX|104  3.429952209
R_PTL_S7_5|_RX|B3 _PTL_S7_5|_RX|7 _PTL_S7_5|_RX|107  2.7439617672
L_PTL_S7_5|_RX|RB1 _PTL_S7_5|_RX|101 0  2.38752113364072e-12
L_PTL_S7_5|_RX|RB2 _PTL_S7_5|_RX|104 0  1.937922998085e-12
L_PTL_S7_5|_RX|RB3 _PTL_S7_5|_RX|107 0  1.550338398468e-12
B_PTL_S8_5|_TX|1 _PTL_S8_5|_TX|1 _PTL_S8_5|_TX|2 JJMIT AREA=2.5
B_PTL_S8_5|_TX|2 _PTL_S8_5|_TX|4 _PTL_S8_5|_TX|5 JJMIT AREA=2.5
I_PTL_S8_5|_TX|B1 0 _PTL_S8_5|_TX|3  PWL(0 0 5e-12 0.000175)
I_PTL_S8_5|_TX|B2 0 _PTL_S8_5|_TX|6  PWL(0 0 5e-12 0.000175)
L_PTL_S8_5|_TX|B1 _PTL_S8_5|_TX|1 _PTL_S8_5|_TX|3  1.684e-12
L_PTL_S8_5|_TX|B2 _PTL_S8_5|_TX|4 _PTL_S8_5|_TX|6  3.596e-12
L_PTL_S8_5|_TX|1 S8_5_TX _PTL_S8_5|_TX|1  2.063e-12
L_PTL_S8_5|_TX|2 _PTL_S8_5|_TX|1 _PTL_S8_5|_TX|4  4.123e-12
L_PTL_S8_5|_TX|3 _PTL_S8_5|_TX|4 _PTL_S8_5|_TX|7  2.193e-12
R_PTL_S8_5|_TX|D _PTL_S8_5|_TX|7 _PTL_S8_5|A_PTL  1.36
L_PTL_S8_5|_TX|P1 _PTL_S8_5|_TX|2 0  5.254e-13
L_PTL_S8_5|_TX|P2 _PTL_S8_5|_TX|5 0  5.141e-13
R_PTL_S8_5|_TX|B1 _PTL_S8_5|_TX|1 _PTL_S8_5|_TX|101  2.7439617672
R_PTL_S8_5|_TX|B2 _PTL_S8_5|_TX|4 _PTL_S8_5|_TX|104  2.7439617672
L_PTL_S8_5|_TX|RB1 _PTL_S8_5|_TX|101 0  1.550338398468e-12
L_PTL_S8_5|_TX|RB2 _PTL_S8_5|_TX|104 0  1.550338398468e-12
B_PTL_S8_5|_RX|1 _PTL_S8_5|_RX|1 _PTL_S8_5|_RX|2 JJMIT AREA=1.6233766233766234
B_PTL_S8_5|_RX|2 _PTL_S8_5|_RX|4 _PTL_S8_5|_RX|5 JJMIT AREA=2.0
B_PTL_S8_5|_RX|3 _PTL_S8_5|_RX|7 _PTL_S8_5|_RX|8 JJMIT AREA=2.5
I_PTL_S8_5|_RX|B1 0 _PTL_S8_5|_RX|3  PWL(0 0 5e-12 0.000162338)
L_PTL_S8_5|_RX|B1 _PTL_S8_5|_RX|1 _PTL_S8_5|_RX|3  2.777e-12
I_PTL_S8_5|_RX|B2 0 _PTL_S8_5|_RX|6  PWL(0 0 5e-12 0.00014)
L_PTL_S8_5|_RX|B2 _PTL_S8_5|_RX|4 _PTL_S8_5|_RX|6  2.685e-12
I_PTL_S8_5|_RX|B3 0 _PTL_S8_5|_RX|9  PWL(0 0 5e-12 0.000175)
L_PTL_S8_5|_RX|B3 _PTL_S8_5|_RX|7 _PTL_S8_5|_RX|9  2.764e-12
L_PTL_S8_5|_RX|1 _PTL_S8_5|A_PTL _PTL_S8_5|_RX|1  1.346e-12
L_PTL_S8_5|_RX|2 _PTL_S8_5|_RX|1 _PTL_S8_5|_RX|4  6.348e-12
L_PTL_S8_5|_RX|3 _PTL_S8_5|_RX|4 _PTL_S8_5|_RX|7  5.197e-12
L_PTL_S8_5|_RX|4 _PTL_S8_5|_RX|7 S8_5  2.058e-12
L_PTL_S8_5|_RX|P1 _PTL_S8_5|_RX|2 0  4.795e-13
L_PTL_S8_5|_RX|P2 _PTL_S8_5|_RX|5 0  5.431e-13
L_PTL_S8_5|_RX|P3 _PTL_S8_5|_RX|8 0  5.339e-13
R_PTL_S8_5|_RX|B1 _PTL_S8_5|_RX|1 _PTL_S8_5|_RX|101  4.225701121488
R_PTL_S8_5|_RX|B2 _PTL_S8_5|_RX|4 _PTL_S8_5|_RX|104  3.429952209
R_PTL_S8_5|_RX|B3 _PTL_S8_5|_RX|7 _PTL_S8_5|_RX|107  2.7439617672
L_PTL_S8_5|_RX|RB1 _PTL_S8_5|_RX|101 0  2.38752113364072e-12
L_PTL_S8_5|_RX|RB2 _PTL_S8_5|_RX|104 0  1.937922998085e-12
L_PTL_S8_5|_RX|RB3 _PTL_S8_5|_RX|107 0  1.550338398468e-12
LI0|_SPL_A|I_D1|B I0|_SPL_A|D1 I0|_SPL_A|I_D1|MID  2e-12
II0|_SPL_A|I_D1|B 0 I0|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_D2|B I0|_SPL_A|D2 I0|_SPL_A|I_D2|MID  2e-12
II0|_SPL_A|I_D2|B 0 I0|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_A|I_Q1|B I0|_SPL_A|QA1 I0|_SPL_A|I_Q1|MID  2e-12
II0|_SPL_A|I_Q1|B 0 I0|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_Q2|B I0|_SPL_A|QB1 I0|_SPL_A|I_Q2|MID  2e-12
II0|_SPL_A|I_Q2|B 0 I0|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_A|1|1 I0|_SPL_A|D1 I0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|1|P I0|_SPL_A|1|MID_SERIES 0  2e-13
RI0|_SPL_A|1|B I0|_SPL_A|D1 I0|_SPL_A|1|MID_SHUNT  2.7439617672
LI0|_SPL_A|1|RB I0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|2|1 I0|_SPL_A|D2 I0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|2|P I0|_SPL_A|2|MID_SERIES 0  2e-13
RI0|_SPL_A|2|B I0|_SPL_A|D2 I0|_SPL_A|2|MID_SHUNT  2.7439617672
LI0|_SPL_A|2|RB I0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|A|1 I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|A|P I0|_SPL_A|A|MID_SERIES 0  2e-13
RI0|_SPL_A|A|B I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SHUNT  2.7439617672
LI0|_SPL_A|A|RB I0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|B|1 I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|B|P I0|_SPL_A|B|MID_SERIES 0  2e-13
RI0|_SPL_A|B|B I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SHUNT  2.7439617672
LI0|_SPL_A|B|RB I0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_B|I_D1|B I0|_SPL_B|D1 I0|_SPL_B|I_D1|MID  2e-12
II0|_SPL_B|I_D1|B 0 I0|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_D2|B I0|_SPL_B|D2 I0|_SPL_B|I_D2|MID  2e-12
II0|_SPL_B|I_D2|B 0 I0|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_B|I_Q1|B I0|_SPL_B|QA1 I0|_SPL_B|I_Q1|MID  2e-12
II0|_SPL_B|I_Q1|B 0 I0|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_Q2|B I0|_SPL_B|QB1 I0|_SPL_B|I_Q2|MID  2e-12
II0|_SPL_B|I_Q2|B 0 I0|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_B|1|1 I0|_SPL_B|D1 I0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|1|P I0|_SPL_B|1|MID_SERIES 0  2e-13
RI0|_SPL_B|1|B I0|_SPL_B|D1 I0|_SPL_B|1|MID_SHUNT  2.7439617672
LI0|_SPL_B|1|RB I0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|2|1 I0|_SPL_B|D2 I0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|2|P I0|_SPL_B|2|MID_SERIES 0  2e-13
RI0|_SPL_B|2|B I0|_SPL_B|D2 I0|_SPL_B|2|MID_SHUNT  2.7439617672
LI0|_SPL_B|2|RB I0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|A|1 I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|A|P I0|_SPL_B|A|MID_SERIES 0  2e-13
RI0|_SPL_B|A|B I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SHUNT  2.7439617672
LI0|_SPL_B|A|RB I0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|B|1 I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|B|P I0|_SPL_B|B|MID_SERIES 0  2e-13
RI0|_SPL_B|B|B I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SHUNT  2.7439617672
LI0|_SPL_B|B|RB I0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_A|I_1|B I0|_DFF_A|A1 I0|_DFF_A|I_1|MID  2e-12
II0|_DFF_A|I_1|B 0 I0|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_3|B I0|_DFF_A|A3 I0|_DFF_A|I_3|MID  2e-12
II0|_DFF_A|I_3|B 0 I0|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_A|I_T|B I0|_DFF_A|T1 I0|_DFF_A|I_T|MID  2e-12
II0|_DFF_A|I_T|B 0 I0|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_6|B I0|_DFF_A|Q1 I0|_DFF_A|I_6|MID  2e-12
II0|_DFF_A|I_6|B 0 I0|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_A|1|1 I0|_DFF_A|A1 I0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|1|P I0|_DFF_A|1|MID_SERIES 0  2e-13
RI0|_DFF_A|1|B I0|_DFF_A|A1 I0|_DFF_A|1|MID_SHUNT  2.7439617672
LI0|_DFF_A|1|RB I0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|23|1 I0|_DFF_A|A2 I0|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|23|B I0|_DFF_A|A2 I0|_DFF_A|23|MID_SHUNT  3.84154647408
LI0|_DFF_A|23|RB I0|_DFF_A|23|MID_SHUNT I0|_DFF_A|A3  2.1704737578552e-12
BI0|_DFF_A|3|1 I0|_DFF_A|A3 I0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|3|P I0|_DFF_A|3|MID_SERIES 0  2e-13
RI0|_DFF_A|3|B I0|_DFF_A|A3 I0|_DFF_A|3|MID_SHUNT  2.7439617672
LI0|_DFF_A|3|RB I0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|4|1 I0|_DFF_A|A4 I0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|4|P I0|_DFF_A|4|MID_SERIES 0  2e-13
RI0|_DFF_A|4|B I0|_DFF_A|A4 I0|_DFF_A|4|MID_SHUNT  2.7439617672
LI0|_DFF_A|4|RB I0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|T|1 I0|_DFF_A|T1 I0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|T|P I0|_DFF_A|T|MID_SERIES 0  2e-13
RI0|_DFF_A|T|B I0|_DFF_A|T1 I0|_DFF_A|T|MID_SHUNT  2.7439617672
LI0|_DFF_A|T|RB I0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|45|1 I0|_DFF_A|T2 I0|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|45|B I0|_DFF_A|T2 I0|_DFF_A|45|MID_SHUNT  3.84154647408
LI0|_DFF_A|45|RB I0|_DFF_A|45|MID_SHUNT I0|_DFF_A|A4  2.1704737578552e-12
BI0|_DFF_A|6|1 I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|6|P I0|_DFF_A|6|MID_SERIES 0  2e-13
RI0|_DFF_A|6|B I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SHUNT  2.7439617672
LI0|_DFF_A|6|RB I0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_B|I_1|B I0|_DFF_B|A1 I0|_DFF_B|I_1|MID  2e-12
II0|_DFF_B|I_1|B 0 I0|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_3|B I0|_DFF_B|A3 I0|_DFF_B|I_3|MID  2e-12
II0|_DFF_B|I_3|B 0 I0|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_B|I_T|B I0|_DFF_B|T1 I0|_DFF_B|I_T|MID  2e-12
II0|_DFF_B|I_T|B 0 I0|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_6|B I0|_DFF_B|Q1 I0|_DFF_B|I_6|MID  2e-12
II0|_DFF_B|I_6|B 0 I0|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_B|1|1 I0|_DFF_B|A1 I0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|1|P I0|_DFF_B|1|MID_SERIES 0  2e-13
RI0|_DFF_B|1|B I0|_DFF_B|A1 I0|_DFF_B|1|MID_SHUNT  2.7439617672
LI0|_DFF_B|1|RB I0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|23|1 I0|_DFF_B|A2 I0|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|23|B I0|_DFF_B|A2 I0|_DFF_B|23|MID_SHUNT  3.84154647408
LI0|_DFF_B|23|RB I0|_DFF_B|23|MID_SHUNT I0|_DFF_B|A3  2.1704737578552e-12
BI0|_DFF_B|3|1 I0|_DFF_B|A3 I0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|3|P I0|_DFF_B|3|MID_SERIES 0  2e-13
RI0|_DFF_B|3|B I0|_DFF_B|A3 I0|_DFF_B|3|MID_SHUNT  2.7439617672
LI0|_DFF_B|3|RB I0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|4|1 I0|_DFF_B|A4 I0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|4|P I0|_DFF_B|4|MID_SERIES 0  2e-13
RI0|_DFF_B|4|B I0|_DFF_B|A4 I0|_DFF_B|4|MID_SHUNT  2.7439617672
LI0|_DFF_B|4|RB I0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|T|1 I0|_DFF_B|T1 I0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|T|P I0|_DFF_B|T|MID_SERIES 0  2e-13
RI0|_DFF_B|T|B I0|_DFF_B|T1 I0|_DFF_B|T|MID_SHUNT  2.7439617672
LI0|_DFF_B|T|RB I0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|45|1 I0|_DFF_B|T2 I0|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|45|B I0|_DFF_B|T2 I0|_DFF_B|45|MID_SHUNT  3.84154647408
LI0|_DFF_B|45|RB I0|_DFF_B|45|MID_SHUNT I0|_DFF_B|A4  2.1704737578552e-12
BI0|_DFF_B|6|1 I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|6|P I0|_DFF_B|6|MID_SERIES 0  2e-13
RI0|_DFF_B|6|B I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SHUNT  2.7439617672
LI0|_DFF_B|6|RB I0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI0|_XOR|I_A1|B I0|_XOR|A1 I0|_XOR|I_A1|MID  2e-12
II0|_XOR|I_A1|B 0 I0|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_A3|B I0|_XOR|A3 I0|_XOR|I_A3|MID  2e-12
II0|_XOR|I_A3|B 0 I0|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B1|B I0|_XOR|B1 I0|_XOR|I_B1|MID  2e-12
II0|_XOR|I_B1|B 0 I0|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B3|B I0|_XOR|B3 I0|_XOR|I_B3|MID  2e-12
II0|_XOR|I_B3|B 0 I0|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_Q1|B I0|_XOR|Q1 I0|_XOR|I_Q1|MID  2e-12
II0|_XOR|I_Q1|B 0 I0|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_XOR|A1|1 I0|_XOR|A1 I0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A1|P I0|_XOR|A1|MID_SERIES 0  5e-13
RI0|_XOR|A1|B I0|_XOR|A1 I0|_XOR|A1|MID_SHUNT  2.7439617672
LI0|_XOR|A1|RB I0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A2|1 I0|_XOR|A2 I0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A2|P I0|_XOR|A2|MID_SERIES 0  5e-13
RI0|_XOR|A2|B I0|_XOR|A2 I0|_XOR|A2|MID_SHUNT  2.7439617672
LI0|_XOR|A2|RB I0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A3|1 I0|_XOR|A2 I0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A3|P I0|_XOR|A3|MID_SERIES I0|_XOR|A3  1.2e-12
RI0|_XOR|A3|B I0|_XOR|A2 I0|_XOR|A3|MID_SHUNT  2.7439617672
LI0|_XOR|A3|RB I0|_XOR|A3|MID_SHUNT I0|_XOR|A3  2.050338398468e-12
BI0|_XOR|B1|1 I0|_XOR|B1 I0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B1|P I0|_XOR|B1|MID_SERIES 0  5e-13
RI0|_XOR|B1|B I0|_XOR|B1 I0|_XOR|B1|MID_SHUNT  2.7439617672
LI0|_XOR|B1|RB I0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B2|1 I0|_XOR|B2 I0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B2|P I0|_XOR|B2|MID_SERIES 0  5e-13
RI0|_XOR|B2|B I0|_XOR|B2 I0|_XOR|B2|MID_SHUNT  2.7439617672
LI0|_XOR|B2|RB I0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B3|1 I0|_XOR|B2 I0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B3|P I0|_XOR|B3|MID_SERIES I0|_XOR|B3  1.2e-12
RI0|_XOR|B3|B I0|_XOR|B2 I0|_XOR|B3|MID_SHUNT  2.7439617672
LI0|_XOR|B3|RB I0|_XOR|B3|MID_SHUNT I0|_XOR|B3  2.050338398468e-12
BI0|_XOR|T1|1 I0|_XOR|T1 I0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|T1|P I0|_XOR|T1|MID_SERIES 0  5e-13
RI0|_XOR|T1|B I0|_XOR|T1 I0|_XOR|T1|MID_SHUNT  2.7439617672
LI0|_XOR|T1|RB I0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|T2|1 I0|_XOR|T2 I0|_XOR|ABTQ JJMIT AREA=2.0
RI0|_XOR|T2|B I0|_XOR|T2 I0|_XOR|T2|MID_SHUNT  3.429952209
LI0|_XOR|T2|RB I0|_XOR|T2|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|AB|1 I0|_XOR|AB I0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI0|_XOR|AB|P I0|_XOR|AB|MID_SERIES I0|_XOR|ABTQ  1.2e-12
RI0|_XOR|AB|B I0|_XOR|AB I0|_XOR|AB|MID_SHUNT  3.429952209
LI0|_XOR|AB|RB I0|_XOR|AB|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|ABTQ|1 I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|ABTQ|P I0|_XOR|ABTQ|MID_SERIES 0  5e-13
RI0|_XOR|ABTQ|B I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI0|_XOR|ABTQ|RB I0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|Q1|1 I0|_XOR|Q1 I0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|Q1|P I0|_XOR|Q1|MID_SERIES 0  5e-13
RI0|_XOR|Q1|B I0|_XOR|Q1 I0|_XOR|Q1|MID_SHUNT  2.7439617672
LI0|_XOR|Q1|RB I0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI0|_AND|I_A1|B I0|_AND|A1 I0|_AND|I_A1|MID  2e-12
II0|_AND|I_A1|B 0 I0|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_B1|B I0|_AND|B1 I0|_AND|I_B1|MID  2e-12
II0|_AND|I_B1|B 0 I0|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q3|B I0|_AND|Q3 I0|_AND|I_Q3|MID  2e-12
II0|_AND|I_Q3|B 0 I0|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0|_AND|I_Q2|B I0|_AND|Q2 I0|_AND|I_Q2|MID  2e-12
II0|_AND|I_Q2|B 0 I0|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q1|B I0|_AND|Q1 I0|_AND|I_Q1|MID  2e-12
II0|_AND|I_Q1|B 0 I0|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_AND|A1|1 I0|_AND|A1 I0|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A1|P I0|_AND|A1|MID_SERIES 0  2e-13
RI0|_AND|A1|B I0|_AND|A1 I0|_AND|A1|MID_SHUNT  2.7439617672
LI0|_AND|A1|RB I0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A2|1 I0|_AND|A2 I0|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A2|P I0|_AND|A2|MID_SERIES 0  2e-13
RI0|_AND|A2|B I0|_AND|A2 I0|_AND|A2|MID_SHUNT  2.7439617672
LI0|_AND|A2|RB I0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A12|1 I0|_AND|A2 I0|_AND|A3 JJMIT AREA=1.7857142857142858
RI0|_AND|A12|B I0|_AND|A2 I0|_AND|A12|MID_SHUNT  3.84154647408
LI0|_AND|A12|RB I0|_AND|A12|MID_SHUNT I0|_AND|A3  2.1704737578552e-12
BI0|_AND|B1|1 I0|_AND|B1 I0|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B1|P I0|_AND|B1|MID_SERIES 0  2e-13
RI0|_AND|B1|B I0|_AND|B1 I0|_AND|B1|MID_SHUNT  2.7439617672
LI0|_AND|B1|RB I0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B2|1 I0|_AND|B2 I0|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B2|P I0|_AND|B2|MID_SERIES 0  2e-13
RI0|_AND|B2|B I0|_AND|B2 I0|_AND|B2|MID_SHUNT  2.7439617672
LI0|_AND|B2|RB I0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B12|1 I0|_AND|B2 I0|_AND|B3 JJMIT AREA=1.7857142857142858
RI0|_AND|B12|B I0|_AND|B2 I0|_AND|B12|MID_SHUNT  3.84154647408
LI0|_AND|B12|RB I0|_AND|B12|MID_SHUNT I0|_AND|B3  2.1704737578552e-12
BI0|_AND|Q2|1 I0|_AND|Q2 I0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q2|P I0|_AND|Q2|MID_SERIES 0  2e-13
RI0|_AND|Q2|B I0|_AND|Q2 I0|_AND|Q2|MID_SHUNT  2.7439617672
LI0|_AND|Q2|RB I0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|Q1|1 I0|_AND|Q1 I0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q1|P I0|_AND|Q1|MID_SERIES 0  2e-13
RI0|_AND|Q1|B I0|_AND|Q1 I0|_AND|Q1|MID_SHUNT  2.7439617672
LI0|_AND|Q1|RB I0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_A|I_D1|B I1|_SPL_A|D1 I1|_SPL_A|I_D1|MID  2e-12
II1|_SPL_A|I_D1|B 0 I1|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_D2|B I1|_SPL_A|D2 I1|_SPL_A|I_D2|MID  2e-12
II1|_SPL_A|I_D2|B 0 I1|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_A|I_Q1|B I1|_SPL_A|QA1 I1|_SPL_A|I_Q1|MID  2e-12
II1|_SPL_A|I_Q1|B 0 I1|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_Q2|B I1|_SPL_A|QB1 I1|_SPL_A|I_Q2|MID  2e-12
II1|_SPL_A|I_Q2|B 0 I1|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_A|1|1 I1|_SPL_A|D1 I1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|1|P I1|_SPL_A|1|MID_SERIES 0  2e-13
RI1|_SPL_A|1|B I1|_SPL_A|D1 I1|_SPL_A|1|MID_SHUNT  2.7439617672
LI1|_SPL_A|1|RB I1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|2|1 I1|_SPL_A|D2 I1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|2|P I1|_SPL_A|2|MID_SERIES 0  2e-13
RI1|_SPL_A|2|B I1|_SPL_A|D2 I1|_SPL_A|2|MID_SHUNT  2.7439617672
LI1|_SPL_A|2|RB I1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|A|1 I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|A|P I1|_SPL_A|A|MID_SERIES 0  2e-13
RI1|_SPL_A|A|B I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SHUNT  2.7439617672
LI1|_SPL_A|A|RB I1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|B|1 I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|B|P I1|_SPL_A|B|MID_SERIES 0  2e-13
RI1|_SPL_A|B|B I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SHUNT  2.7439617672
LI1|_SPL_A|B|RB I1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_B|I_D1|B I1|_SPL_B|D1 I1|_SPL_B|I_D1|MID  2e-12
II1|_SPL_B|I_D1|B 0 I1|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_D2|B I1|_SPL_B|D2 I1|_SPL_B|I_D2|MID  2e-12
II1|_SPL_B|I_D2|B 0 I1|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_B|I_Q1|B I1|_SPL_B|QA1 I1|_SPL_B|I_Q1|MID  2e-12
II1|_SPL_B|I_Q1|B 0 I1|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_Q2|B I1|_SPL_B|QB1 I1|_SPL_B|I_Q2|MID  2e-12
II1|_SPL_B|I_Q2|B 0 I1|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_B|1|1 I1|_SPL_B|D1 I1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|1|P I1|_SPL_B|1|MID_SERIES 0  2e-13
RI1|_SPL_B|1|B I1|_SPL_B|D1 I1|_SPL_B|1|MID_SHUNT  2.7439617672
LI1|_SPL_B|1|RB I1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|2|1 I1|_SPL_B|D2 I1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|2|P I1|_SPL_B|2|MID_SERIES 0  2e-13
RI1|_SPL_B|2|B I1|_SPL_B|D2 I1|_SPL_B|2|MID_SHUNT  2.7439617672
LI1|_SPL_B|2|RB I1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|A|1 I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|A|P I1|_SPL_B|A|MID_SERIES 0  2e-13
RI1|_SPL_B|A|B I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SHUNT  2.7439617672
LI1|_SPL_B|A|RB I1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|B|1 I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|B|P I1|_SPL_B|B|MID_SERIES 0  2e-13
RI1|_SPL_B|B|B I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SHUNT  2.7439617672
LI1|_SPL_B|B|RB I1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_A|I_1|B I1|_DFF_A|A1 I1|_DFF_A|I_1|MID  2e-12
II1|_DFF_A|I_1|B 0 I1|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_3|B I1|_DFF_A|A3 I1|_DFF_A|I_3|MID  2e-12
II1|_DFF_A|I_3|B 0 I1|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_A|I_T|B I1|_DFF_A|T1 I1|_DFF_A|I_T|MID  2e-12
II1|_DFF_A|I_T|B 0 I1|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_6|B I1|_DFF_A|Q1 I1|_DFF_A|I_6|MID  2e-12
II1|_DFF_A|I_6|B 0 I1|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_A|1|1 I1|_DFF_A|A1 I1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|1|P I1|_DFF_A|1|MID_SERIES 0  2e-13
RI1|_DFF_A|1|B I1|_DFF_A|A1 I1|_DFF_A|1|MID_SHUNT  2.7439617672
LI1|_DFF_A|1|RB I1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|23|1 I1|_DFF_A|A2 I1|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|23|B I1|_DFF_A|A2 I1|_DFF_A|23|MID_SHUNT  3.84154647408
LI1|_DFF_A|23|RB I1|_DFF_A|23|MID_SHUNT I1|_DFF_A|A3  2.1704737578552e-12
BI1|_DFF_A|3|1 I1|_DFF_A|A3 I1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|3|P I1|_DFF_A|3|MID_SERIES 0  2e-13
RI1|_DFF_A|3|B I1|_DFF_A|A3 I1|_DFF_A|3|MID_SHUNT  2.7439617672
LI1|_DFF_A|3|RB I1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|4|1 I1|_DFF_A|A4 I1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|4|P I1|_DFF_A|4|MID_SERIES 0  2e-13
RI1|_DFF_A|4|B I1|_DFF_A|A4 I1|_DFF_A|4|MID_SHUNT  2.7439617672
LI1|_DFF_A|4|RB I1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|T|1 I1|_DFF_A|T1 I1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|T|P I1|_DFF_A|T|MID_SERIES 0  2e-13
RI1|_DFF_A|T|B I1|_DFF_A|T1 I1|_DFF_A|T|MID_SHUNT  2.7439617672
LI1|_DFF_A|T|RB I1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|45|1 I1|_DFF_A|T2 I1|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|45|B I1|_DFF_A|T2 I1|_DFF_A|45|MID_SHUNT  3.84154647408
LI1|_DFF_A|45|RB I1|_DFF_A|45|MID_SHUNT I1|_DFF_A|A4  2.1704737578552e-12
BI1|_DFF_A|6|1 I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|6|P I1|_DFF_A|6|MID_SERIES 0  2e-13
RI1|_DFF_A|6|B I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SHUNT  2.7439617672
LI1|_DFF_A|6|RB I1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_B|I_1|B I1|_DFF_B|A1 I1|_DFF_B|I_1|MID  2e-12
II1|_DFF_B|I_1|B 0 I1|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_3|B I1|_DFF_B|A3 I1|_DFF_B|I_3|MID  2e-12
II1|_DFF_B|I_3|B 0 I1|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_B|I_T|B I1|_DFF_B|T1 I1|_DFF_B|I_T|MID  2e-12
II1|_DFF_B|I_T|B 0 I1|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_6|B I1|_DFF_B|Q1 I1|_DFF_B|I_6|MID  2e-12
II1|_DFF_B|I_6|B 0 I1|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_B|1|1 I1|_DFF_B|A1 I1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|1|P I1|_DFF_B|1|MID_SERIES 0  2e-13
RI1|_DFF_B|1|B I1|_DFF_B|A1 I1|_DFF_B|1|MID_SHUNT  2.7439617672
LI1|_DFF_B|1|RB I1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|23|1 I1|_DFF_B|A2 I1|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|23|B I1|_DFF_B|A2 I1|_DFF_B|23|MID_SHUNT  3.84154647408
LI1|_DFF_B|23|RB I1|_DFF_B|23|MID_SHUNT I1|_DFF_B|A3  2.1704737578552e-12
BI1|_DFF_B|3|1 I1|_DFF_B|A3 I1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|3|P I1|_DFF_B|3|MID_SERIES 0  2e-13
RI1|_DFF_B|3|B I1|_DFF_B|A3 I1|_DFF_B|3|MID_SHUNT  2.7439617672
LI1|_DFF_B|3|RB I1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|4|1 I1|_DFF_B|A4 I1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|4|P I1|_DFF_B|4|MID_SERIES 0  2e-13
RI1|_DFF_B|4|B I1|_DFF_B|A4 I1|_DFF_B|4|MID_SHUNT  2.7439617672
LI1|_DFF_B|4|RB I1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|T|1 I1|_DFF_B|T1 I1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|T|P I1|_DFF_B|T|MID_SERIES 0  2e-13
RI1|_DFF_B|T|B I1|_DFF_B|T1 I1|_DFF_B|T|MID_SHUNT  2.7439617672
LI1|_DFF_B|T|RB I1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|45|1 I1|_DFF_B|T2 I1|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|45|B I1|_DFF_B|T2 I1|_DFF_B|45|MID_SHUNT  3.84154647408
LI1|_DFF_B|45|RB I1|_DFF_B|45|MID_SHUNT I1|_DFF_B|A4  2.1704737578552e-12
BI1|_DFF_B|6|1 I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|6|P I1|_DFF_B|6|MID_SERIES 0  2e-13
RI1|_DFF_B|6|B I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SHUNT  2.7439617672
LI1|_DFF_B|6|RB I1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI1|_XOR|I_A1|B I1|_XOR|A1 I1|_XOR|I_A1|MID  2e-12
II1|_XOR|I_A1|B 0 I1|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_A3|B I1|_XOR|A3 I1|_XOR|I_A3|MID  2e-12
II1|_XOR|I_A3|B 0 I1|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B1|B I1|_XOR|B1 I1|_XOR|I_B1|MID  2e-12
II1|_XOR|I_B1|B 0 I1|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B3|B I1|_XOR|B3 I1|_XOR|I_B3|MID  2e-12
II1|_XOR|I_B3|B 0 I1|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_Q1|B I1|_XOR|Q1 I1|_XOR|I_Q1|MID  2e-12
II1|_XOR|I_Q1|B 0 I1|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_XOR|A1|1 I1|_XOR|A1 I1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A1|P I1|_XOR|A1|MID_SERIES 0  5e-13
RI1|_XOR|A1|B I1|_XOR|A1 I1|_XOR|A1|MID_SHUNT  2.7439617672
LI1|_XOR|A1|RB I1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A2|1 I1|_XOR|A2 I1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A2|P I1|_XOR|A2|MID_SERIES 0  5e-13
RI1|_XOR|A2|B I1|_XOR|A2 I1|_XOR|A2|MID_SHUNT  2.7439617672
LI1|_XOR|A2|RB I1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A3|1 I1|_XOR|A2 I1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A3|P I1|_XOR|A3|MID_SERIES I1|_XOR|A3  1.2e-12
RI1|_XOR|A3|B I1|_XOR|A2 I1|_XOR|A3|MID_SHUNT  2.7439617672
LI1|_XOR|A3|RB I1|_XOR|A3|MID_SHUNT I1|_XOR|A3  2.050338398468e-12
BI1|_XOR|B1|1 I1|_XOR|B1 I1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B1|P I1|_XOR|B1|MID_SERIES 0  5e-13
RI1|_XOR|B1|B I1|_XOR|B1 I1|_XOR|B1|MID_SHUNT  2.7439617672
LI1|_XOR|B1|RB I1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B2|1 I1|_XOR|B2 I1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B2|P I1|_XOR|B2|MID_SERIES 0  5e-13
RI1|_XOR|B2|B I1|_XOR|B2 I1|_XOR|B2|MID_SHUNT  2.7439617672
LI1|_XOR|B2|RB I1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B3|1 I1|_XOR|B2 I1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B3|P I1|_XOR|B3|MID_SERIES I1|_XOR|B3  1.2e-12
RI1|_XOR|B3|B I1|_XOR|B2 I1|_XOR|B3|MID_SHUNT  2.7439617672
LI1|_XOR|B3|RB I1|_XOR|B3|MID_SHUNT I1|_XOR|B3  2.050338398468e-12
BI1|_XOR|T1|1 I1|_XOR|T1 I1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|T1|P I1|_XOR|T1|MID_SERIES 0  5e-13
RI1|_XOR|T1|B I1|_XOR|T1 I1|_XOR|T1|MID_SHUNT  2.7439617672
LI1|_XOR|T1|RB I1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|T2|1 I1|_XOR|T2 I1|_XOR|ABTQ JJMIT AREA=2.0
RI1|_XOR|T2|B I1|_XOR|T2 I1|_XOR|T2|MID_SHUNT  3.429952209
LI1|_XOR|T2|RB I1|_XOR|T2|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|AB|1 I1|_XOR|AB I1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI1|_XOR|AB|P I1|_XOR|AB|MID_SERIES I1|_XOR|ABTQ  1.2e-12
RI1|_XOR|AB|B I1|_XOR|AB I1|_XOR|AB|MID_SHUNT  3.429952209
LI1|_XOR|AB|RB I1|_XOR|AB|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|ABTQ|1 I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|ABTQ|P I1|_XOR|ABTQ|MID_SERIES 0  5e-13
RI1|_XOR|ABTQ|B I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI1|_XOR|ABTQ|RB I1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|Q1|1 I1|_XOR|Q1 I1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|Q1|P I1|_XOR|Q1|MID_SERIES 0  5e-13
RI1|_XOR|Q1|B I1|_XOR|Q1 I1|_XOR|Q1|MID_SHUNT  2.7439617672
LI1|_XOR|Q1|RB I1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI1|_AND|I_A1|B I1|_AND|A1 I1|_AND|I_A1|MID  2e-12
II1|_AND|I_A1|B 0 I1|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_B1|B I1|_AND|B1 I1|_AND|I_B1|MID  2e-12
II1|_AND|I_B1|B 0 I1|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q3|B I1|_AND|Q3 I1|_AND|I_Q3|MID  2e-12
II1|_AND|I_Q3|B 0 I1|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1|_AND|I_Q2|B I1|_AND|Q2 I1|_AND|I_Q2|MID  2e-12
II1|_AND|I_Q2|B 0 I1|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q1|B I1|_AND|Q1 I1|_AND|I_Q1|MID  2e-12
II1|_AND|I_Q1|B 0 I1|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_AND|A1|1 I1|_AND|A1 I1|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A1|P I1|_AND|A1|MID_SERIES 0  2e-13
RI1|_AND|A1|B I1|_AND|A1 I1|_AND|A1|MID_SHUNT  2.7439617672
LI1|_AND|A1|RB I1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A2|1 I1|_AND|A2 I1|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A2|P I1|_AND|A2|MID_SERIES 0  2e-13
RI1|_AND|A2|B I1|_AND|A2 I1|_AND|A2|MID_SHUNT  2.7439617672
LI1|_AND|A2|RB I1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A12|1 I1|_AND|A2 I1|_AND|A3 JJMIT AREA=1.7857142857142858
RI1|_AND|A12|B I1|_AND|A2 I1|_AND|A12|MID_SHUNT  3.84154647408
LI1|_AND|A12|RB I1|_AND|A12|MID_SHUNT I1|_AND|A3  2.1704737578552e-12
BI1|_AND|B1|1 I1|_AND|B1 I1|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B1|P I1|_AND|B1|MID_SERIES 0  2e-13
RI1|_AND|B1|B I1|_AND|B1 I1|_AND|B1|MID_SHUNT  2.7439617672
LI1|_AND|B1|RB I1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B2|1 I1|_AND|B2 I1|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B2|P I1|_AND|B2|MID_SERIES 0  2e-13
RI1|_AND|B2|B I1|_AND|B2 I1|_AND|B2|MID_SHUNT  2.7439617672
LI1|_AND|B2|RB I1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B12|1 I1|_AND|B2 I1|_AND|B3 JJMIT AREA=1.7857142857142858
RI1|_AND|B12|B I1|_AND|B2 I1|_AND|B12|MID_SHUNT  3.84154647408
LI1|_AND|B12|RB I1|_AND|B12|MID_SHUNT I1|_AND|B3  2.1704737578552e-12
BI1|_AND|Q2|1 I1|_AND|Q2 I1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q2|P I1|_AND|Q2|MID_SERIES 0  2e-13
RI1|_AND|Q2|B I1|_AND|Q2 I1|_AND|Q2|MID_SHUNT  2.7439617672
LI1|_AND|Q2|RB I1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|Q1|1 I1|_AND|Q1 I1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q1|P I1|_AND|Q1|MID_SERIES 0  2e-13
RI1|_AND|Q1|B I1|_AND|Q1 I1|_AND|Q1|MID_SHUNT  2.7439617672
LI1|_AND|Q1|RB I1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_A|I_D1|B I2|_SPL_A|D1 I2|_SPL_A|I_D1|MID  2e-12
II2|_SPL_A|I_D1|B 0 I2|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_D2|B I2|_SPL_A|D2 I2|_SPL_A|I_D2|MID  2e-12
II2|_SPL_A|I_D2|B 0 I2|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_A|I_Q1|B I2|_SPL_A|QA1 I2|_SPL_A|I_Q1|MID  2e-12
II2|_SPL_A|I_Q1|B 0 I2|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_Q2|B I2|_SPL_A|QB1 I2|_SPL_A|I_Q2|MID  2e-12
II2|_SPL_A|I_Q2|B 0 I2|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_A|1|1 I2|_SPL_A|D1 I2|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|1|P I2|_SPL_A|1|MID_SERIES 0  2e-13
RI2|_SPL_A|1|B I2|_SPL_A|D1 I2|_SPL_A|1|MID_SHUNT  2.7439617672
LI2|_SPL_A|1|RB I2|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|2|1 I2|_SPL_A|D2 I2|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|2|P I2|_SPL_A|2|MID_SERIES 0  2e-13
RI2|_SPL_A|2|B I2|_SPL_A|D2 I2|_SPL_A|2|MID_SHUNT  2.7439617672
LI2|_SPL_A|2|RB I2|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|A|1 I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|A|P I2|_SPL_A|A|MID_SERIES 0  2e-13
RI2|_SPL_A|A|B I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SHUNT  2.7439617672
LI2|_SPL_A|A|RB I2|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|B|1 I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|B|P I2|_SPL_A|B|MID_SERIES 0  2e-13
RI2|_SPL_A|B|B I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SHUNT  2.7439617672
LI2|_SPL_A|B|RB I2|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_B|I_D1|B I2|_SPL_B|D1 I2|_SPL_B|I_D1|MID  2e-12
II2|_SPL_B|I_D1|B 0 I2|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_D2|B I2|_SPL_B|D2 I2|_SPL_B|I_D2|MID  2e-12
II2|_SPL_B|I_D2|B 0 I2|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_B|I_Q1|B I2|_SPL_B|QA1 I2|_SPL_B|I_Q1|MID  2e-12
II2|_SPL_B|I_Q1|B 0 I2|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_Q2|B I2|_SPL_B|QB1 I2|_SPL_B|I_Q2|MID  2e-12
II2|_SPL_B|I_Q2|B 0 I2|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_B|1|1 I2|_SPL_B|D1 I2|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|1|P I2|_SPL_B|1|MID_SERIES 0  2e-13
RI2|_SPL_B|1|B I2|_SPL_B|D1 I2|_SPL_B|1|MID_SHUNT  2.7439617672
LI2|_SPL_B|1|RB I2|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|2|1 I2|_SPL_B|D2 I2|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|2|P I2|_SPL_B|2|MID_SERIES 0  2e-13
RI2|_SPL_B|2|B I2|_SPL_B|D2 I2|_SPL_B|2|MID_SHUNT  2.7439617672
LI2|_SPL_B|2|RB I2|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|A|1 I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|A|P I2|_SPL_B|A|MID_SERIES 0  2e-13
RI2|_SPL_B|A|B I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SHUNT  2.7439617672
LI2|_SPL_B|A|RB I2|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|B|1 I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|B|P I2|_SPL_B|B|MID_SERIES 0  2e-13
RI2|_SPL_B|B|B I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SHUNT  2.7439617672
LI2|_SPL_B|B|RB I2|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_A|I_1|B I2|_DFF_A|A1 I2|_DFF_A|I_1|MID  2e-12
II2|_DFF_A|I_1|B 0 I2|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_3|B I2|_DFF_A|A3 I2|_DFF_A|I_3|MID  2e-12
II2|_DFF_A|I_3|B 0 I2|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_A|I_T|B I2|_DFF_A|T1 I2|_DFF_A|I_T|MID  2e-12
II2|_DFF_A|I_T|B 0 I2|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_6|B I2|_DFF_A|Q1 I2|_DFF_A|I_6|MID  2e-12
II2|_DFF_A|I_6|B 0 I2|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_A|1|1 I2|_DFF_A|A1 I2|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|1|P I2|_DFF_A|1|MID_SERIES 0  2e-13
RI2|_DFF_A|1|B I2|_DFF_A|A1 I2|_DFF_A|1|MID_SHUNT  2.7439617672
LI2|_DFF_A|1|RB I2|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|23|1 I2|_DFF_A|A2 I2|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|23|B I2|_DFF_A|A2 I2|_DFF_A|23|MID_SHUNT  3.84154647408
LI2|_DFF_A|23|RB I2|_DFF_A|23|MID_SHUNT I2|_DFF_A|A3  2.1704737578552e-12
BI2|_DFF_A|3|1 I2|_DFF_A|A3 I2|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|3|P I2|_DFF_A|3|MID_SERIES 0  2e-13
RI2|_DFF_A|3|B I2|_DFF_A|A3 I2|_DFF_A|3|MID_SHUNT  2.7439617672
LI2|_DFF_A|3|RB I2|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|4|1 I2|_DFF_A|A4 I2|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|4|P I2|_DFF_A|4|MID_SERIES 0  2e-13
RI2|_DFF_A|4|B I2|_DFF_A|A4 I2|_DFF_A|4|MID_SHUNT  2.7439617672
LI2|_DFF_A|4|RB I2|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|T|1 I2|_DFF_A|T1 I2|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|T|P I2|_DFF_A|T|MID_SERIES 0  2e-13
RI2|_DFF_A|T|B I2|_DFF_A|T1 I2|_DFF_A|T|MID_SHUNT  2.7439617672
LI2|_DFF_A|T|RB I2|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|45|1 I2|_DFF_A|T2 I2|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|45|B I2|_DFF_A|T2 I2|_DFF_A|45|MID_SHUNT  3.84154647408
LI2|_DFF_A|45|RB I2|_DFF_A|45|MID_SHUNT I2|_DFF_A|A4  2.1704737578552e-12
BI2|_DFF_A|6|1 I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|6|P I2|_DFF_A|6|MID_SERIES 0  2e-13
RI2|_DFF_A|6|B I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SHUNT  2.7439617672
LI2|_DFF_A|6|RB I2|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_B|I_1|B I2|_DFF_B|A1 I2|_DFF_B|I_1|MID  2e-12
II2|_DFF_B|I_1|B 0 I2|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_3|B I2|_DFF_B|A3 I2|_DFF_B|I_3|MID  2e-12
II2|_DFF_B|I_3|B 0 I2|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_B|I_T|B I2|_DFF_B|T1 I2|_DFF_B|I_T|MID  2e-12
II2|_DFF_B|I_T|B 0 I2|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_6|B I2|_DFF_B|Q1 I2|_DFF_B|I_6|MID  2e-12
II2|_DFF_B|I_6|B 0 I2|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_B|1|1 I2|_DFF_B|A1 I2|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|1|P I2|_DFF_B|1|MID_SERIES 0  2e-13
RI2|_DFF_B|1|B I2|_DFF_B|A1 I2|_DFF_B|1|MID_SHUNT  2.7439617672
LI2|_DFF_B|1|RB I2|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|23|1 I2|_DFF_B|A2 I2|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|23|B I2|_DFF_B|A2 I2|_DFF_B|23|MID_SHUNT  3.84154647408
LI2|_DFF_B|23|RB I2|_DFF_B|23|MID_SHUNT I2|_DFF_B|A3  2.1704737578552e-12
BI2|_DFF_B|3|1 I2|_DFF_B|A3 I2|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|3|P I2|_DFF_B|3|MID_SERIES 0  2e-13
RI2|_DFF_B|3|B I2|_DFF_B|A3 I2|_DFF_B|3|MID_SHUNT  2.7439617672
LI2|_DFF_B|3|RB I2|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|4|1 I2|_DFF_B|A4 I2|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|4|P I2|_DFF_B|4|MID_SERIES 0  2e-13
RI2|_DFF_B|4|B I2|_DFF_B|A4 I2|_DFF_B|4|MID_SHUNT  2.7439617672
LI2|_DFF_B|4|RB I2|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|T|1 I2|_DFF_B|T1 I2|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|T|P I2|_DFF_B|T|MID_SERIES 0  2e-13
RI2|_DFF_B|T|B I2|_DFF_B|T1 I2|_DFF_B|T|MID_SHUNT  2.7439617672
LI2|_DFF_B|T|RB I2|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|45|1 I2|_DFF_B|T2 I2|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|45|B I2|_DFF_B|T2 I2|_DFF_B|45|MID_SHUNT  3.84154647408
LI2|_DFF_B|45|RB I2|_DFF_B|45|MID_SHUNT I2|_DFF_B|A4  2.1704737578552e-12
BI2|_DFF_B|6|1 I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|6|P I2|_DFF_B|6|MID_SERIES 0  2e-13
RI2|_DFF_B|6|B I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SHUNT  2.7439617672
LI2|_DFF_B|6|RB I2|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI2|_XOR|I_A1|B I2|_XOR|A1 I2|_XOR|I_A1|MID  2e-12
II2|_XOR|I_A1|B 0 I2|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_A3|B I2|_XOR|A3 I2|_XOR|I_A3|MID  2e-12
II2|_XOR|I_A3|B 0 I2|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B1|B I2|_XOR|B1 I2|_XOR|I_B1|MID  2e-12
II2|_XOR|I_B1|B 0 I2|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B3|B I2|_XOR|B3 I2|_XOR|I_B3|MID  2e-12
II2|_XOR|I_B3|B 0 I2|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_Q1|B I2|_XOR|Q1 I2|_XOR|I_Q1|MID  2e-12
II2|_XOR|I_Q1|B 0 I2|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_XOR|A1|1 I2|_XOR|A1 I2|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A1|P I2|_XOR|A1|MID_SERIES 0  5e-13
RI2|_XOR|A1|B I2|_XOR|A1 I2|_XOR|A1|MID_SHUNT  2.7439617672
LI2|_XOR|A1|RB I2|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A2|1 I2|_XOR|A2 I2|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A2|P I2|_XOR|A2|MID_SERIES 0  5e-13
RI2|_XOR|A2|B I2|_XOR|A2 I2|_XOR|A2|MID_SHUNT  2.7439617672
LI2|_XOR|A2|RB I2|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A3|1 I2|_XOR|A2 I2|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A3|P I2|_XOR|A3|MID_SERIES I2|_XOR|A3  1.2e-12
RI2|_XOR|A3|B I2|_XOR|A2 I2|_XOR|A3|MID_SHUNT  2.7439617672
LI2|_XOR|A3|RB I2|_XOR|A3|MID_SHUNT I2|_XOR|A3  2.050338398468e-12
BI2|_XOR|B1|1 I2|_XOR|B1 I2|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B1|P I2|_XOR|B1|MID_SERIES 0  5e-13
RI2|_XOR|B1|B I2|_XOR|B1 I2|_XOR|B1|MID_SHUNT  2.7439617672
LI2|_XOR|B1|RB I2|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B2|1 I2|_XOR|B2 I2|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B2|P I2|_XOR|B2|MID_SERIES 0  5e-13
RI2|_XOR|B2|B I2|_XOR|B2 I2|_XOR|B2|MID_SHUNT  2.7439617672
LI2|_XOR|B2|RB I2|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B3|1 I2|_XOR|B2 I2|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B3|P I2|_XOR|B3|MID_SERIES I2|_XOR|B3  1.2e-12
RI2|_XOR|B3|B I2|_XOR|B2 I2|_XOR|B3|MID_SHUNT  2.7439617672
LI2|_XOR|B3|RB I2|_XOR|B3|MID_SHUNT I2|_XOR|B3  2.050338398468e-12
BI2|_XOR|T1|1 I2|_XOR|T1 I2|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|T1|P I2|_XOR|T1|MID_SERIES 0  5e-13
RI2|_XOR|T1|B I2|_XOR|T1 I2|_XOR|T1|MID_SHUNT  2.7439617672
LI2|_XOR|T1|RB I2|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|T2|1 I2|_XOR|T2 I2|_XOR|ABTQ JJMIT AREA=2.0
RI2|_XOR|T2|B I2|_XOR|T2 I2|_XOR|T2|MID_SHUNT  3.429952209
LI2|_XOR|T2|RB I2|_XOR|T2|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|AB|1 I2|_XOR|AB I2|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI2|_XOR|AB|P I2|_XOR|AB|MID_SERIES I2|_XOR|ABTQ  1.2e-12
RI2|_XOR|AB|B I2|_XOR|AB I2|_XOR|AB|MID_SHUNT  3.429952209
LI2|_XOR|AB|RB I2|_XOR|AB|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|ABTQ|1 I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|ABTQ|P I2|_XOR|ABTQ|MID_SERIES 0  5e-13
RI2|_XOR|ABTQ|B I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI2|_XOR|ABTQ|RB I2|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|Q1|1 I2|_XOR|Q1 I2|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|Q1|P I2|_XOR|Q1|MID_SERIES 0  5e-13
RI2|_XOR|Q1|B I2|_XOR|Q1 I2|_XOR|Q1|MID_SHUNT  2.7439617672
LI2|_XOR|Q1|RB I2|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI2|_AND|I_A1|B I2|_AND|A1 I2|_AND|I_A1|MID  2e-12
II2|_AND|I_A1|B 0 I2|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_B1|B I2|_AND|B1 I2|_AND|I_B1|MID  2e-12
II2|_AND|I_B1|B 0 I2|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q3|B I2|_AND|Q3 I2|_AND|I_Q3|MID  2e-12
II2|_AND|I_Q3|B 0 I2|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2|_AND|I_Q2|B I2|_AND|Q2 I2|_AND|I_Q2|MID  2e-12
II2|_AND|I_Q2|B 0 I2|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q1|B I2|_AND|Q1 I2|_AND|I_Q1|MID  2e-12
II2|_AND|I_Q1|B 0 I2|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_AND|A1|1 I2|_AND|A1 I2|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A1|P I2|_AND|A1|MID_SERIES 0  2e-13
RI2|_AND|A1|B I2|_AND|A1 I2|_AND|A1|MID_SHUNT  2.7439617672
LI2|_AND|A1|RB I2|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A2|1 I2|_AND|A2 I2|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A2|P I2|_AND|A2|MID_SERIES 0  2e-13
RI2|_AND|A2|B I2|_AND|A2 I2|_AND|A2|MID_SHUNT  2.7439617672
LI2|_AND|A2|RB I2|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A12|1 I2|_AND|A2 I2|_AND|A3 JJMIT AREA=1.7857142857142858
RI2|_AND|A12|B I2|_AND|A2 I2|_AND|A12|MID_SHUNT  3.84154647408
LI2|_AND|A12|RB I2|_AND|A12|MID_SHUNT I2|_AND|A3  2.1704737578552e-12
BI2|_AND|B1|1 I2|_AND|B1 I2|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B1|P I2|_AND|B1|MID_SERIES 0  2e-13
RI2|_AND|B1|B I2|_AND|B1 I2|_AND|B1|MID_SHUNT  2.7439617672
LI2|_AND|B1|RB I2|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B2|1 I2|_AND|B2 I2|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B2|P I2|_AND|B2|MID_SERIES 0  2e-13
RI2|_AND|B2|B I2|_AND|B2 I2|_AND|B2|MID_SHUNT  2.7439617672
LI2|_AND|B2|RB I2|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B12|1 I2|_AND|B2 I2|_AND|B3 JJMIT AREA=1.7857142857142858
RI2|_AND|B12|B I2|_AND|B2 I2|_AND|B12|MID_SHUNT  3.84154647408
LI2|_AND|B12|RB I2|_AND|B12|MID_SHUNT I2|_AND|B3  2.1704737578552e-12
BI2|_AND|Q2|1 I2|_AND|Q2 I2|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q2|P I2|_AND|Q2|MID_SERIES 0  2e-13
RI2|_AND|Q2|B I2|_AND|Q2 I2|_AND|Q2|MID_SHUNT  2.7439617672
LI2|_AND|Q2|RB I2|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|Q1|1 I2|_AND|Q1 I2|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q1|P I2|_AND|Q1|MID_SERIES 0  2e-13
RI2|_AND|Q1|B I2|_AND|Q1 I2|_AND|Q1|MID_SHUNT  2.7439617672
LI2|_AND|Q1|RB I2|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_A|I_D1|B I3|_SPL_A|D1 I3|_SPL_A|I_D1|MID  2e-12
II3|_SPL_A|I_D1|B 0 I3|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_D2|B I3|_SPL_A|D2 I3|_SPL_A|I_D2|MID  2e-12
II3|_SPL_A|I_D2|B 0 I3|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_A|I_Q1|B I3|_SPL_A|QA1 I3|_SPL_A|I_Q1|MID  2e-12
II3|_SPL_A|I_Q1|B 0 I3|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_Q2|B I3|_SPL_A|QB1 I3|_SPL_A|I_Q2|MID  2e-12
II3|_SPL_A|I_Q2|B 0 I3|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_A|1|1 I3|_SPL_A|D1 I3|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|1|P I3|_SPL_A|1|MID_SERIES 0  2e-13
RI3|_SPL_A|1|B I3|_SPL_A|D1 I3|_SPL_A|1|MID_SHUNT  2.7439617672
LI3|_SPL_A|1|RB I3|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|2|1 I3|_SPL_A|D2 I3|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|2|P I3|_SPL_A|2|MID_SERIES 0  2e-13
RI3|_SPL_A|2|B I3|_SPL_A|D2 I3|_SPL_A|2|MID_SHUNT  2.7439617672
LI3|_SPL_A|2|RB I3|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|A|1 I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|A|P I3|_SPL_A|A|MID_SERIES 0  2e-13
RI3|_SPL_A|A|B I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SHUNT  2.7439617672
LI3|_SPL_A|A|RB I3|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|B|1 I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|B|P I3|_SPL_A|B|MID_SERIES 0  2e-13
RI3|_SPL_A|B|B I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SHUNT  2.7439617672
LI3|_SPL_A|B|RB I3|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_B|I_D1|B I3|_SPL_B|D1 I3|_SPL_B|I_D1|MID  2e-12
II3|_SPL_B|I_D1|B 0 I3|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_D2|B I3|_SPL_B|D2 I3|_SPL_B|I_D2|MID  2e-12
II3|_SPL_B|I_D2|B 0 I3|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_B|I_Q1|B I3|_SPL_B|QA1 I3|_SPL_B|I_Q1|MID  2e-12
II3|_SPL_B|I_Q1|B 0 I3|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_Q2|B I3|_SPL_B|QB1 I3|_SPL_B|I_Q2|MID  2e-12
II3|_SPL_B|I_Q2|B 0 I3|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_B|1|1 I3|_SPL_B|D1 I3|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|1|P I3|_SPL_B|1|MID_SERIES 0  2e-13
RI3|_SPL_B|1|B I3|_SPL_B|D1 I3|_SPL_B|1|MID_SHUNT  2.7439617672
LI3|_SPL_B|1|RB I3|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|2|1 I3|_SPL_B|D2 I3|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|2|P I3|_SPL_B|2|MID_SERIES 0  2e-13
RI3|_SPL_B|2|B I3|_SPL_B|D2 I3|_SPL_B|2|MID_SHUNT  2.7439617672
LI3|_SPL_B|2|RB I3|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|A|1 I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|A|P I3|_SPL_B|A|MID_SERIES 0  2e-13
RI3|_SPL_B|A|B I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SHUNT  2.7439617672
LI3|_SPL_B|A|RB I3|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|B|1 I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|B|P I3|_SPL_B|B|MID_SERIES 0  2e-13
RI3|_SPL_B|B|B I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SHUNT  2.7439617672
LI3|_SPL_B|B|RB I3|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_A|I_1|B I3|_DFF_A|A1 I3|_DFF_A|I_1|MID  2e-12
II3|_DFF_A|I_1|B 0 I3|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_3|B I3|_DFF_A|A3 I3|_DFF_A|I_3|MID  2e-12
II3|_DFF_A|I_3|B 0 I3|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_A|I_T|B I3|_DFF_A|T1 I3|_DFF_A|I_T|MID  2e-12
II3|_DFF_A|I_T|B 0 I3|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_6|B I3|_DFF_A|Q1 I3|_DFF_A|I_6|MID  2e-12
II3|_DFF_A|I_6|B 0 I3|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_A|1|1 I3|_DFF_A|A1 I3|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|1|P I3|_DFF_A|1|MID_SERIES 0  2e-13
RI3|_DFF_A|1|B I3|_DFF_A|A1 I3|_DFF_A|1|MID_SHUNT  2.7439617672
LI3|_DFF_A|1|RB I3|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|23|1 I3|_DFF_A|A2 I3|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|23|B I3|_DFF_A|A2 I3|_DFF_A|23|MID_SHUNT  3.84154647408
LI3|_DFF_A|23|RB I3|_DFF_A|23|MID_SHUNT I3|_DFF_A|A3  2.1704737578552e-12
BI3|_DFF_A|3|1 I3|_DFF_A|A3 I3|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|3|P I3|_DFF_A|3|MID_SERIES 0  2e-13
RI3|_DFF_A|3|B I3|_DFF_A|A3 I3|_DFF_A|3|MID_SHUNT  2.7439617672
LI3|_DFF_A|3|RB I3|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|4|1 I3|_DFF_A|A4 I3|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|4|P I3|_DFF_A|4|MID_SERIES 0  2e-13
RI3|_DFF_A|4|B I3|_DFF_A|A4 I3|_DFF_A|4|MID_SHUNT  2.7439617672
LI3|_DFF_A|4|RB I3|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|T|1 I3|_DFF_A|T1 I3|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|T|P I3|_DFF_A|T|MID_SERIES 0  2e-13
RI3|_DFF_A|T|B I3|_DFF_A|T1 I3|_DFF_A|T|MID_SHUNT  2.7439617672
LI3|_DFF_A|T|RB I3|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|45|1 I3|_DFF_A|T2 I3|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|45|B I3|_DFF_A|T2 I3|_DFF_A|45|MID_SHUNT  3.84154647408
LI3|_DFF_A|45|RB I3|_DFF_A|45|MID_SHUNT I3|_DFF_A|A4  2.1704737578552e-12
BI3|_DFF_A|6|1 I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|6|P I3|_DFF_A|6|MID_SERIES 0  2e-13
RI3|_DFF_A|6|B I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SHUNT  2.7439617672
LI3|_DFF_A|6|RB I3|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_B|I_1|B I3|_DFF_B|A1 I3|_DFF_B|I_1|MID  2e-12
II3|_DFF_B|I_1|B 0 I3|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_3|B I3|_DFF_B|A3 I3|_DFF_B|I_3|MID  2e-12
II3|_DFF_B|I_3|B 0 I3|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_B|I_T|B I3|_DFF_B|T1 I3|_DFF_B|I_T|MID  2e-12
II3|_DFF_B|I_T|B 0 I3|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_6|B I3|_DFF_B|Q1 I3|_DFF_B|I_6|MID  2e-12
II3|_DFF_B|I_6|B 0 I3|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_B|1|1 I3|_DFF_B|A1 I3|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|1|P I3|_DFF_B|1|MID_SERIES 0  2e-13
RI3|_DFF_B|1|B I3|_DFF_B|A1 I3|_DFF_B|1|MID_SHUNT  2.7439617672
LI3|_DFF_B|1|RB I3|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|23|1 I3|_DFF_B|A2 I3|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|23|B I3|_DFF_B|A2 I3|_DFF_B|23|MID_SHUNT  3.84154647408
LI3|_DFF_B|23|RB I3|_DFF_B|23|MID_SHUNT I3|_DFF_B|A3  2.1704737578552e-12
BI3|_DFF_B|3|1 I3|_DFF_B|A3 I3|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|3|P I3|_DFF_B|3|MID_SERIES 0  2e-13
RI3|_DFF_B|3|B I3|_DFF_B|A3 I3|_DFF_B|3|MID_SHUNT  2.7439617672
LI3|_DFF_B|3|RB I3|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|4|1 I3|_DFF_B|A4 I3|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|4|P I3|_DFF_B|4|MID_SERIES 0  2e-13
RI3|_DFF_B|4|B I3|_DFF_B|A4 I3|_DFF_B|4|MID_SHUNT  2.7439617672
LI3|_DFF_B|4|RB I3|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|T|1 I3|_DFF_B|T1 I3|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|T|P I3|_DFF_B|T|MID_SERIES 0  2e-13
RI3|_DFF_B|T|B I3|_DFF_B|T1 I3|_DFF_B|T|MID_SHUNT  2.7439617672
LI3|_DFF_B|T|RB I3|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|45|1 I3|_DFF_B|T2 I3|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|45|B I3|_DFF_B|T2 I3|_DFF_B|45|MID_SHUNT  3.84154647408
LI3|_DFF_B|45|RB I3|_DFF_B|45|MID_SHUNT I3|_DFF_B|A4  2.1704737578552e-12
BI3|_DFF_B|6|1 I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|6|P I3|_DFF_B|6|MID_SERIES 0  2e-13
RI3|_DFF_B|6|B I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SHUNT  2.7439617672
LI3|_DFF_B|6|RB I3|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI3|_XOR|I_A1|B I3|_XOR|A1 I3|_XOR|I_A1|MID  2e-12
II3|_XOR|I_A1|B 0 I3|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_A3|B I3|_XOR|A3 I3|_XOR|I_A3|MID  2e-12
II3|_XOR|I_A3|B 0 I3|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B1|B I3|_XOR|B1 I3|_XOR|I_B1|MID  2e-12
II3|_XOR|I_B1|B 0 I3|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B3|B I3|_XOR|B3 I3|_XOR|I_B3|MID  2e-12
II3|_XOR|I_B3|B 0 I3|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_Q1|B I3|_XOR|Q1 I3|_XOR|I_Q1|MID  2e-12
II3|_XOR|I_Q1|B 0 I3|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_XOR|A1|1 I3|_XOR|A1 I3|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A1|P I3|_XOR|A1|MID_SERIES 0  5e-13
RI3|_XOR|A1|B I3|_XOR|A1 I3|_XOR|A1|MID_SHUNT  2.7439617672
LI3|_XOR|A1|RB I3|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A2|1 I3|_XOR|A2 I3|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A2|P I3|_XOR|A2|MID_SERIES 0  5e-13
RI3|_XOR|A2|B I3|_XOR|A2 I3|_XOR|A2|MID_SHUNT  2.7439617672
LI3|_XOR|A2|RB I3|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A3|1 I3|_XOR|A2 I3|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A3|P I3|_XOR|A3|MID_SERIES I3|_XOR|A3  1.2e-12
RI3|_XOR|A3|B I3|_XOR|A2 I3|_XOR|A3|MID_SHUNT  2.7439617672
LI3|_XOR|A3|RB I3|_XOR|A3|MID_SHUNT I3|_XOR|A3  2.050338398468e-12
BI3|_XOR|B1|1 I3|_XOR|B1 I3|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B1|P I3|_XOR|B1|MID_SERIES 0  5e-13
RI3|_XOR|B1|B I3|_XOR|B1 I3|_XOR|B1|MID_SHUNT  2.7439617672
LI3|_XOR|B1|RB I3|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B2|1 I3|_XOR|B2 I3|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B2|P I3|_XOR|B2|MID_SERIES 0  5e-13
RI3|_XOR|B2|B I3|_XOR|B2 I3|_XOR|B2|MID_SHUNT  2.7439617672
LI3|_XOR|B2|RB I3|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B3|1 I3|_XOR|B2 I3|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B3|P I3|_XOR|B3|MID_SERIES I3|_XOR|B3  1.2e-12
RI3|_XOR|B3|B I3|_XOR|B2 I3|_XOR|B3|MID_SHUNT  2.7439617672
LI3|_XOR|B3|RB I3|_XOR|B3|MID_SHUNT I3|_XOR|B3  2.050338398468e-12
BI3|_XOR|T1|1 I3|_XOR|T1 I3|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|T1|P I3|_XOR|T1|MID_SERIES 0  5e-13
RI3|_XOR|T1|B I3|_XOR|T1 I3|_XOR|T1|MID_SHUNT  2.7439617672
LI3|_XOR|T1|RB I3|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|T2|1 I3|_XOR|T2 I3|_XOR|ABTQ JJMIT AREA=2.0
RI3|_XOR|T2|B I3|_XOR|T2 I3|_XOR|T2|MID_SHUNT  3.429952209
LI3|_XOR|T2|RB I3|_XOR|T2|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|AB|1 I3|_XOR|AB I3|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI3|_XOR|AB|P I3|_XOR|AB|MID_SERIES I3|_XOR|ABTQ  1.2e-12
RI3|_XOR|AB|B I3|_XOR|AB I3|_XOR|AB|MID_SHUNT  3.429952209
LI3|_XOR|AB|RB I3|_XOR|AB|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|ABTQ|1 I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|ABTQ|P I3|_XOR|ABTQ|MID_SERIES 0  5e-13
RI3|_XOR|ABTQ|B I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI3|_XOR|ABTQ|RB I3|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|Q1|1 I3|_XOR|Q1 I3|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|Q1|P I3|_XOR|Q1|MID_SERIES 0  5e-13
RI3|_XOR|Q1|B I3|_XOR|Q1 I3|_XOR|Q1|MID_SHUNT  2.7439617672
LI3|_XOR|Q1|RB I3|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI3|_AND|I_A1|B I3|_AND|A1 I3|_AND|I_A1|MID  2e-12
II3|_AND|I_A1|B 0 I3|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_B1|B I3|_AND|B1 I3|_AND|I_B1|MID  2e-12
II3|_AND|I_B1|B 0 I3|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q3|B I3|_AND|Q3 I3|_AND|I_Q3|MID  2e-12
II3|_AND|I_Q3|B 0 I3|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3|_AND|I_Q2|B I3|_AND|Q2 I3|_AND|I_Q2|MID  2e-12
II3|_AND|I_Q2|B 0 I3|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q1|B I3|_AND|Q1 I3|_AND|I_Q1|MID  2e-12
II3|_AND|I_Q1|B 0 I3|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_AND|A1|1 I3|_AND|A1 I3|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A1|P I3|_AND|A1|MID_SERIES 0  2e-13
RI3|_AND|A1|B I3|_AND|A1 I3|_AND|A1|MID_SHUNT  2.7439617672
LI3|_AND|A1|RB I3|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A2|1 I3|_AND|A2 I3|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A2|P I3|_AND|A2|MID_SERIES 0  2e-13
RI3|_AND|A2|B I3|_AND|A2 I3|_AND|A2|MID_SHUNT  2.7439617672
LI3|_AND|A2|RB I3|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A12|1 I3|_AND|A2 I3|_AND|A3 JJMIT AREA=1.7857142857142858
RI3|_AND|A12|B I3|_AND|A2 I3|_AND|A12|MID_SHUNT  3.84154647408
LI3|_AND|A12|RB I3|_AND|A12|MID_SHUNT I3|_AND|A3  2.1704737578552e-12
BI3|_AND|B1|1 I3|_AND|B1 I3|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B1|P I3|_AND|B1|MID_SERIES 0  2e-13
RI3|_AND|B1|B I3|_AND|B1 I3|_AND|B1|MID_SHUNT  2.7439617672
LI3|_AND|B1|RB I3|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B2|1 I3|_AND|B2 I3|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B2|P I3|_AND|B2|MID_SERIES 0  2e-13
RI3|_AND|B2|B I3|_AND|B2 I3|_AND|B2|MID_SHUNT  2.7439617672
LI3|_AND|B2|RB I3|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B12|1 I3|_AND|B2 I3|_AND|B3 JJMIT AREA=1.7857142857142858
RI3|_AND|B12|B I3|_AND|B2 I3|_AND|B12|MID_SHUNT  3.84154647408
LI3|_AND|B12|RB I3|_AND|B12|MID_SHUNT I3|_AND|B3  2.1704737578552e-12
BI3|_AND|Q2|1 I3|_AND|Q2 I3|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q2|P I3|_AND|Q2|MID_SERIES 0  2e-13
RI3|_AND|Q2|B I3|_AND|Q2 I3|_AND|Q2|MID_SHUNT  2.7439617672
LI3|_AND|Q2|RB I3|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|Q1|1 I3|_AND|Q1 I3|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q1|P I3|_AND|Q1|MID_SERIES 0  2e-13
RI3|_AND|Q1|B I3|_AND|Q1 I3|_AND|Q1|MID_SHUNT  2.7439617672
LI3|_AND|Q1|RB I3|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI4|_SPL_A|I_D1|B I4|_SPL_A|D1 I4|_SPL_A|I_D1|MID  2e-12
II4|_SPL_A|I_D1|B 0 I4|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI4|_SPL_A|I_D2|B I4|_SPL_A|D2 I4|_SPL_A|I_D2|MID  2e-12
II4|_SPL_A|I_D2|B 0 I4|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI4|_SPL_A|I_Q1|B I4|_SPL_A|QA1 I4|_SPL_A|I_Q1|MID  2e-12
II4|_SPL_A|I_Q1|B 0 I4|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI4|_SPL_A|I_Q2|B I4|_SPL_A|QB1 I4|_SPL_A|I_Q2|MID  2e-12
II4|_SPL_A|I_Q2|B 0 I4|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI4|_SPL_A|1|1 I4|_SPL_A|D1 I4|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_A|1|P I4|_SPL_A|1|MID_SERIES 0  2e-13
RI4|_SPL_A|1|B I4|_SPL_A|D1 I4|_SPL_A|1|MID_SHUNT  2.7439617672
LI4|_SPL_A|1|RB I4|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI4|_SPL_A|2|1 I4|_SPL_A|D2 I4|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_A|2|P I4|_SPL_A|2|MID_SERIES 0  2e-13
RI4|_SPL_A|2|B I4|_SPL_A|D2 I4|_SPL_A|2|MID_SHUNT  2.7439617672
LI4|_SPL_A|2|RB I4|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI4|_SPL_A|A|1 I4|_SPL_A|QA1 I4|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_A|A|P I4|_SPL_A|A|MID_SERIES 0  2e-13
RI4|_SPL_A|A|B I4|_SPL_A|QA1 I4|_SPL_A|A|MID_SHUNT  2.7439617672
LI4|_SPL_A|A|RB I4|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI4|_SPL_A|B|1 I4|_SPL_A|QB1 I4|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_A|B|P I4|_SPL_A|B|MID_SERIES 0  2e-13
RI4|_SPL_A|B|B I4|_SPL_A|QB1 I4|_SPL_A|B|MID_SHUNT  2.7439617672
LI4|_SPL_A|B|RB I4|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI4|_SPL_B|I_D1|B I4|_SPL_B|D1 I4|_SPL_B|I_D1|MID  2e-12
II4|_SPL_B|I_D1|B 0 I4|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI4|_SPL_B|I_D2|B I4|_SPL_B|D2 I4|_SPL_B|I_D2|MID  2e-12
II4|_SPL_B|I_D2|B 0 I4|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI4|_SPL_B|I_Q1|B I4|_SPL_B|QA1 I4|_SPL_B|I_Q1|MID  2e-12
II4|_SPL_B|I_Q1|B 0 I4|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI4|_SPL_B|I_Q2|B I4|_SPL_B|QB1 I4|_SPL_B|I_Q2|MID  2e-12
II4|_SPL_B|I_Q2|B 0 I4|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI4|_SPL_B|1|1 I4|_SPL_B|D1 I4|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_B|1|P I4|_SPL_B|1|MID_SERIES 0  2e-13
RI4|_SPL_B|1|B I4|_SPL_B|D1 I4|_SPL_B|1|MID_SHUNT  2.7439617672
LI4|_SPL_B|1|RB I4|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI4|_SPL_B|2|1 I4|_SPL_B|D2 I4|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_B|2|P I4|_SPL_B|2|MID_SERIES 0  2e-13
RI4|_SPL_B|2|B I4|_SPL_B|D2 I4|_SPL_B|2|MID_SHUNT  2.7439617672
LI4|_SPL_B|2|RB I4|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI4|_SPL_B|A|1 I4|_SPL_B|QA1 I4|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_B|A|P I4|_SPL_B|A|MID_SERIES 0  2e-13
RI4|_SPL_B|A|B I4|_SPL_B|QA1 I4|_SPL_B|A|MID_SHUNT  2.7439617672
LI4|_SPL_B|A|RB I4|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI4|_SPL_B|B|1 I4|_SPL_B|QB1 I4|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI4|_SPL_B|B|P I4|_SPL_B|B|MID_SERIES 0  2e-13
RI4|_SPL_B|B|B I4|_SPL_B|QB1 I4|_SPL_B|B|MID_SHUNT  2.7439617672
LI4|_SPL_B|B|RB I4|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI4|_DFF_A|I_1|B I4|_DFF_A|A1 I4|_DFF_A|I_1|MID  2e-12
II4|_DFF_A|I_1|B 0 I4|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI4|_DFF_A|I_3|B I4|_DFF_A|A3 I4|_DFF_A|I_3|MID  2e-12
II4|_DFF_A|I_3|B 0 I4|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI4|_DFF_A|I_T|B I4|_DFF_A|T1 I4|_DFF_A|I_T|MID  2e-12
II4|_DFF_A|I_T|B 0 I4|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI4|_DFF_A|I_6|B I4|_DFF_A|Q1 I4|_DFF_A|I_6|MID  2e-12
II4|_DFF_A|I_6|B 0 I4|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI4|_DFF_A|1|1 I4|_DFF_A|A1 I4|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_A|1|P I4|_DFF_A|1|MID_SERIES 0  2e-13
RI4|_DFF_A|1|B I4|_DFF_A|A1 I4|_DFF_A|1|MID_SHUNT  2.7439617672
LI4|_DFF_A|1|RB I4|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_A|23|1 I4|_DFF_A|A2 I4|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI4|_DFF_A|23|B I4|_DFF_A|A2 I4|_DFF_A|23|MID_SHUNT  3.84154647408
LI4|_DFF_A|23|RB I4|_DFF_A|23|MID_SHUNT I4|_DFF_A|A3  2.1704737578552e-12
BI4|_DFF_A|3|1 I4|_DFF_A|A3 I4|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_A|3|P I4|_DFF_A|3|MID_SERIES 0  2e-13
RI4|_DFF_A|3|B I4|_DFF_A|A3 I4|_DFF_A|3|MID_SHUNT  2.7439617672
LI4|_DFF_A|3|RB I4|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_A|4|1 I4|_DFF_A|A4 I4|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_A|4|P I4|_DFF_A|4|MID_SERIES 0  2e-13
RI4|_DFF_A|4|B I4|_DFF_A|A4 I4|_DFF_A|4|MID_SHUNT  2.7439617672
LI4|_DFF_A|4|RB I4|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_A|T|1 I4|_DFF_A|T1 I4|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_A|T|P I4|_DFF_A|T|MID_SERIES 0  2e-13
RI4|_DFF_A|T|B I4|_DFF_A|T1 I4|_DFF_A|T|MID_SHUNT  2.7439617672
LI4|_DFF_A|T|RB I4|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_A|45|1 I4|_DFF_A|T2 I4|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI4|_DFF_A|45|B I4|_DFF_A|T2 I4|_DFF_A|45|MID_SHUNT  3.84154647408
LI4|_DFF_A|45|RB I4|_DFF_A|45|MID_SHUNT I4|_DFF_A|A4  2.1704737578552e-12
BI4|_DFF_A|6|1 I4|_DFF_A|Q1 I4|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_A|6|P I4|_DFF_A|6|MID_SERIES 0  2e-13
RI4|_DFF_A|6|B I4|_DFF_A|Q1 I4|_DFF_A|6|MID_SHUNT  2.7439617672
LI4|_DFF_A|6|RB I4|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI4|_DFF_B|I_1|B I4|_DFF_B|A1 I4|_DFF_B|I_1|MID  2e-12
II4|_DFF_B|I_1|B 0 I4|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI4|_DFF_B|I_3|B I4|_DFF_B|A3 I4|_DFF_B|I_3|MID  2e-12
II4|_DFF_B|I_3|B 0 I4|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI4|_DFF_B|I_T|B I4|_DFF_B|T1 I4|_DFF_B|I_T|MID  2e-12
II4|_DFF_B|I_T|B 0 I4|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI4|_DFF_B|I_6|B I4|_DFF_B|Q1 I4|_DFF_B|I_6|MID  2e-12
II4|_DFF_B|I_6|B 0 I4|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI4|_DFF_B|1|1 I4|_DFF_B|A1 I4|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_B|1|P I4|_DFF_B|1|MID_SERIES 0  2e-13
RI4|_DFF_B|1|B I4|_DFF_B|A1 I4|_DFF_B|1|MID_SHUNT  2.7439617672
LI4|_DFF_B|1|RB I4|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_B|23|1 I4|_DFF_B|A2 I4|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI4|_DFF_B|23|B I4|_DFF_B|A2 I4|_DFF_B|23|MID_SHUNT  3.84154647408
LI4|_DFF_B|23|RB I4|_DFF_B|23|MID_SHUNT I4|_DFF_B|A3  2.1704737578552e-12
BI4|_DFF_B|3|1 I4|_DFF_B|A3 I4|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_B|3|P I4|_DFF_B|3|MID_SERIES 0  2e-13
RI4|_DFF_B|3|B I4|_DFF_B|A3 I4|_DFF_B|3|MID_SHUNT  2.7439617672
LI4|_DFF_B|3|RB I4|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_B|4|1 I4|_DFF_B|A4 I4|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_B|4|P I4|_DFF_B|4|MID_SERIES 0  2e-13
RI4|_DFF_B|4|B I4|_DFF_B|A4 I4|_DFF_B|4|MID_SHUNT  2.7439617672
LI4|_DFF_B|4|RB I4|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_B|T|1 I4|_DFF_B|T1 I4|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_B|T|P I4|_DFF_B|T|MID_SERIES 0  2e-13
RI4|_DFF_B|T|B I4|_DFF_B|T1 I4|_DFF_B|T|MID_SHUNT  2.7439617672
LI4|_DFF_B|T|RB I4|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI4|_DFF_B|45|1 I4|_DFF_B|T2 I4|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI4|_DFF_B|45|B I4|_DFF_B|T2 I4|_DFF_B|45|MID_SHUNT  3.84154647408
LI4|_DFF_B|45|RB I4|_DFF_B|45|MID_SHUNT I4|_DFF_B|A4  2.1704737578552e-12
BI4|_DFF_B|6|1 I4|_DFF_B|Q1 I4|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI4|_DFF_B|6|P I4|_DFF_B|6|MID_SERIES 0  2e-13
RI4|_DFF_B|6|B I4|_DFF_B|Q1 I4|_DFF_B|6|MID_SHUNT  2.7439617672
LI4|_DFF_B|6|RB I4|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI4|_XOR|I_A1|B I4|_XOR|A1 I4|_XOR|I_A1|MID  2e-12
II4|_XOR|I_A1|B 0 I4|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI4|_XOR|I_A3|B I4|_XOR|A3 I4|_XOR|I_A3|MID  2e-12
II4|_XOR|I_A3|B 0 I4|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI4|_XOR|I_B1|B I4|_XOR|B1 I4|_XOR|I_B1|MID  2e-12
II4|_XOR|I_B1|B 0 I4|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI4|_XOR|I_B3|B I4|_XOR|B3 I4|_XOR|I_B3|MID  2e-12
II4|_XOR|I_B3|B 0 I4|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI4|_XOR|I_Q1|B I4|_XOR|Q1 I4|_XOR|I_Q1|MID  2e-12
II4|_XOR|I_Q1|B 0 I4|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI4|_XOR|A1|1 I4|_XOR|A1 I4|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|A1|P I4|_XOR|A1|MID_SERIES 0  5e-13
RI4|_XOR|A1|B I4|_XOR|A1 I4|_XOR|A1|MID_SHUNT  2.7439617672
LI4|_XOR|A1|RB I4|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI4|_XOR|A2|1 I4|_XOR|A2 I4|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|A2|P I4|_XOR|A2|MID_SERIES 0  5e-13
RI4|_XOR|A2|B I4|_XOR|A2 I4|_XOR|A2|MID_SHUNT  2.7439617672
LI4|_XOR|A2|RB I4|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI4|_XOR|A3|1 I4|_XOR|A2 I4|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|A3|P I4|_XOR|A3|MID_SERIES I4|_XOR|A3  1.2e-12
RI4|_XOR|A3|B I4|_XOR|A2 I4|_XOR|A3|MID_SHUNT  2.7439617672
LI4|_XOR|A3|RB I4|_XOR|A3|MID_SHUNT I4|_XOR|A3  2.050338398468e-12
BI4|_XOR|B1|1 I4|_XOR|B1 I4|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|B1|P I4|_XOR|B1|MID_SERIES 0  5e-13
RI4|_XOR|B1|B I4|_XOR|B1 I4|_XOR|B1|MID_SHUNT  2.7439617672
LI4|_XOR|B1|RB I4|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI4|_XOR|B2|1 I4|_XOR|B2 I4|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|B2|P I4|_XOR|B2|MID_SERIES 0  5e-13
RI4|_XOR|B2|B I4|_XOR|B2 I4|_XOR|B2|MID_SHUNT  2.7439617672
LI4|_XOR|B2|RB I4|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI4|_XOR|B3|1 I4|_XOR|B2 I4|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|B3|P I4|_XOR|B3|MID_SERIES I4|_XOR|B3  1.2e-12
RI4|_XOR|B3|B I4|_XOR|B2 I4|_XOR|B3|MID_SHUNT  2.7439617672
LI4|_XOR|B3|RB I4|_XOR|B3|MID_SHUNT I4|_XOR|B3  2.050338398468e-12
BI4|_XOR|T1|1 I4|_XOR|T1 I4|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|T1|P I4|_XOR|T1|MID_SERIES 0  5e-13
RI4|_XOR|T1|B I4|_XOR|T1 I4|_XOR|T1|MID_SHUNT  2.7439617672
LI4|_XOR|T1|RB I4|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI4|_XOR|T2|1 I4|_XOR|T2 I4|_XOR|ABTQ JJMIT AREA=2.0
RI4|_XOR|T2|B I4|_XOR|T2 I4|_XOR|T2|MID_SHUNT  3.429952209
LI4|_XOR|T2|RB I4|_XOR|T2|MID_SHUNT I4|_XOR|ABTQ  2.437922998085e-12
BI4|_XOR|AB|1 I4|_XOR|AB I4|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI4|_XOR|AB|P I4|_XOR|AB|MID_SERIES I4|_XOR|ABTQ  1.2e-12
RI4|_XOR|AB|B I4|_XOR|AB I4|_XOR|AB|MID_SHUNT  3.429952209
LI4|_XOR|AB|RB I4|_XOR|AB|MID_SHUNT I4|_XOR|ABTQ  2.437922998085e-12
BI4|_XOR|ABTQ|1 I4|_XOR|ABTQ I4|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|ABTQ|P I4|_XOR|ABTQ|MID_SERIES 0  5e-13
RI4|_XOR|ABTQ|B I4|_XOR|ABTQ I4|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI4|_XOR|ABTQ|RB I4|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI4|_XOR|Q1|1 I4|_XOR|Q1 I4|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI4|_XOR|Q1|P I4|_XOR|Q1|MID_SERIES 0  5e-13
RI4|_XOR|Q1|B I4|_XOR|Q1 I4|_XOR|Q1|MID_SHUNT  2.7439617672
LI4|_XOR|Q1|RB I4|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI4|_AND|I_A1|B I4|_AND|A1 I4|_AND|I_A1|MID  2e-12
II4|_AND|I_A1|B 0 I4|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI4|_AND|I_B1|B I4|_AND|B1 I4|_AND|I_B1|MID  2e-12
II4|_AND|I_B1|B 0 I4|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI4|_AND|I_Q3|B I4|_AND|Q3 I4|_AND|I_Q3|MID  2e-12
II4|_AND|I_Q3|B 0 I4|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI4|_AND|I_Q2|B I4|_AND|Q2 I4|_AND|I_Q2|MID  2e-12
II4|_AND|I_Q2|B 0 I4|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI4|_AND|I_Q1|B I4|_AND|Q1 I4|_AND|I_Q1|MID  2e-12
II4|_AND|I_Q1|B 0 I4|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI4|_AND|A1|1 I4|_AND|A1 I4|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI4|_AND|A1|P I4|_AND|A1|MID_SERIES 0  2e-13
RI4|_AND|A1|B I4|_AND|A1 I4|_AND|A1|MID_SHUNT  2.7439617672
LI4|_AND|A1|RB I4|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI4|_AND|A2|1 I4|_AND|A2 I4|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI4|_AND|A2|P I4|_AND|A2|MID_SERIES 0  2e-13
RI4|_AND|A2|B I4|_AND|A2 I4|_AND|A2|MID_SHUNT  2.7439617672
LI4|_AND|A2|RB I4|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI4|_AND|A12|1 I4|_AND|A2 I4|_AND|A3 JJMIT AREA=1.7857142857142858
RI4|_AND|A12|B I4|_AND|A2 I4|_AND|A12|MID_SHUNT  3.84154647408
LI4|_AND|A12|RB I4|_AND|A12|MID_SHUNT I4|_AND|A3  2.1704737578552e-12
BI4|_AND|B1|1 I4|_AND|B1 I4|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI4|_AND|B1|P I4|_AND|B1|MID_SERIES 0  2e-13
RI4|_AND|B1|B I4|_AND|B1 I4|_AND|B1|MID_SHUNT  2.7439617672
LI4|_AND|B1|RB I4|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI4|_AND|B2|1 I4|_AND|B2 I4|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI4|_AND|B2|P I4|_AND|B2|MID_SERIES 0  2e-13
RI4|_AND|B2|B I4|_AND|B2 I4|_AND|B2|MID_SHUNT  2.7439617672
LI4|_AND|B2|RB I4|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI4|_AND|B12|1 I4|_AND|B2 I4|_AND|B3 JJMIT AREA=1.7857142857142858
RI4|_AND|B12|B I4|_AND|B2 I4|_AND|B12|MID_SHUNT  3.84154647408
LI4|_AND|B12|RB I4|_AND|B12|MID_SHUNT I4|_AND|B3  2.1704737578552e-12
BI4|_AND|Q2|1 I4|_AND|Q2 I4|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI4|_AND|Q2|P I4|_AND|Q2|MID_SERIES 0  2e-13
RI4|_AND|Q2|B I4|_AND|Q2 I4|_AND|Q2|MID_SHUNT  2.7439617672
LI4|_AND|Q2|RB I4|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI4|_AND|Q1|1 I4|_AND|Q1 I4|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI4|_AND|Q1|P I4|_AND|Q1|MID_SERIES 0  2e-13
RI4|_AND|Q1|B I4|_AND|Q1 I4|_AND|Q1|MID_SHUNT  2.7439617672
LI4|_AND|Q1|RB I4|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI5|_SPL_A|I_D1|B I5|_SPL_A|D1 I5|_SPL_A|I_D1|MID  2e-12
II5|_SPL_A|I_D1|B 0 I5|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI5|_SPL_A|I_D2|B I5|_SPL_A|D2 I5|_SPL_A|I_D2|MID  2e-12
II5|_SPL_A|I_D2|B 0 I5|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI5|_SPL_A|I_Q1|B I5|_SPL_A|QA1 I5|_SPL_A|I_Q1|MID  2e-12
II5|_SPL_A|I_Q1|B 0 I5|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI5|_SPL_A|I_Q2|B I5|_SPL_A|QB1 I5|_SPL_A|I_Q2|MID  2e-12
II5|_SPL_A|I_Q2|B 0 I5|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI5|_SPL_A|1|1 I5|_SPL_A|D1 I5|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_A|1|P I5|_SPL_A|1|MID_SERIES 0  2e-13
RI5|_SPL_A|1|B I5|_SPL_A|D1 I5|_SPL_A|1|MID_SHUNT  2.7439617672
LI5|_SPL_A|1|RB I5|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI5|_SPL_A|2|1 I5|_SPL_A|D2 I5|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_A|2|P I5|_SPL_A|2|MID_SERIES 0  2e-13
RI5|_SPL_A|2|B I5|_SPL_A|D2 I5|_SPL_A|2|MID_SHUNT  2.7439617672
LI5|_SPL_A|2|RB I5|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI5|_SPL_A|A|1 I5|_SPL_A|QA1 I5|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_A|A|P I5|_SPL_A|A|MID_SERIES 0  2e-13
RI5|_SPL_A|A|B I5|_SPL_A|QA1 I5|_SPL_A|A|MID_SHUNT  2.7439617672
LI5|_SPL_A|A|RB I5|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI5|_SPL_A|B|1 I5|_SPL_A|QB1 I5|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_A|B|P I5|_SPL_A|B|MID_SERIES 0  2e-13
RI5|_SPL_A|B|B I5|_SPL_A|QB1 I5|_SPL_A|B|MID_SHUNT  2.7439617672
LI5|_SPL_A|B|RB I5|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI5|_SPL_B|I_D1|B I5|_SPL_B|D1 I5|_SPL_B|I_D1|MID  2e-12
II5|_SPL_B|I_D1|B 0 I5|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI5|_SPL_B|I_D2|B I5|_SPL_B|D2 I5|_SPL_B|I_D2|MID  2e-12
II5|_SPL_B|I_D2|B 0 I5|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI5|_SPL_B|I_Q1|B I5|_SPL_B|QA1 I5|_SPL_B|I_Q1|MID  2e-12
II5|_SPL_B|I_Q1|B 0 I5|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI5|_SPL_B|I_Q2|B I5|_SPL_B|QB1 I5|_SPL_B|I_Q2|MID  2e-12
II5|_SPL_B|I_Q2|B 0 I5|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI5|_SPL_B|1|1 I5|_SPL_B|D1 I5|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_B|1|P I5|_SPL_B|1|MID_SERIES 0  2e-13
RI5|_SPL_B|1|B I5|_SPL_B|D1 I5|_SPL_B|1|MID_SHUNT  2.7439617672
LI5|_SPL_B|1|RB I5|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI5|_SPL_B|2|1 I5|_SPL_B|D2 I5|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_B|2|P I5|_SPL_B|2|MID_SERIES 0  2e-13
RI5|_SPL_B|2|B I5|_SPL_B|D2 I5|_SPL_B|2|MID_SHUNT  2.7439617672
LI5|_SPL_B|2|RB I5|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI5|_SPL_B|A|1 I5|_SPL_B|QA1 I5|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_B|A|P I5|_SPL_B|A|MID_SERIES 0  2e-13
RI5|_SPL_B|A|B I5|_SPL_B|QA1 I5|_SPL_B|A|MID_SHUNT  2.7439617672
LI5|_SPL_B|A|RB I5|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI5|_SPL_B|B|1 I5|_SPL_B|QB1 I5|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI5|_SPL_B|B|P I5|_SPL_B|B|MID_SERIES 0  2e-13
RI5|_SPL_B|B|B I5|_SPL_B|QB1 I5|_SPL_B|B|MID_SHUNT  2.7439617672
LI5|_SPL_B|B|RB I5|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI5|_DFF_A|I_1|B I5|_DFF_A|A1 I5|_DFF_A|I_1|MID  2e-12
II5|_DFF_A|I_1|B 0 I5|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI5|_DFF_A|I_3|B I5|_DFF_A|A3 I5|_DFF_A|I_3|MID  2e-12
II5|_DFF_A|I_3|B 0 I5|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI5|_DFF_A|I_T|B I5|_DFF_A|T1 I5|_DFF_A|I_T|MID  2e-12
II5|_DFF_A|I_T|B 0 I5|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI5|_DFF_A|I_6|B I5|_DFF_A|Q1 I5|_DFF_A|I_6|MID  2e-12
II5|_DFF_A|I_6|B 0 I5|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI5|_DFF_A|1|1 I5|_DFF_A|A1 I5|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_A|1|P I5|_DFF_A|1|MID_SERIES 0  2e-13
RI5|_DFF_A|1|B I5|_DFF_A|A1 I5|_DFF_A|1|MID_SHUNT  2.7439617672
LI5|_DFF_A|1|RB I5|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_A|23|1 I5|_DFF_A|A2 I5|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI5|_DFF_A|23|B I5|_DFF_A|A2 I5|_DFF_A|23|MID_SHUNT  3.84154647408
LI5|_DFF_A|23|RB I5|_DFF_A|23|MID_SHUNT I5|_DFF_A|A3  2.1704737578552e-12
BI5|_DFF_A|3|1 I5|_DFF_A|A3 I5|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_A|3|P I5|_DFF_A|3|MID_SERIES 0  2e-13
RI5|_DFF_A|3|B I5|_DFF_A|A3 I5|_DFF_A|3|MID_SHUNT  2.7439617672
LI5|_DFF_A|3|RB I5|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_A|4|1 I5|_DFF_A|A4 I5|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_A|4|P I5|_DFF_A|4|MID_SERIES 0  2e-13
RI5|_DFF_A|4|B I5|_DFF_A|A4 I5|_DFF_A|4|MID_SHUNT  2.7439617672
LI5|_DFF_A|4|RB I5|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_A|T|1 I5|_DFF_A|T1 I5|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_A|T|P I5|_DFF_A|T|MID_SERIES 0  2e-13
RI5|_DFF_A|T|B I5|_DFF_A|T1 I5|_DFF_A|T|MID_SHUNT  2.7439617672
LI5|_DFF_A|T|RB I5|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_A|45|1 I5|_DFF_A|T2 I5|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI5|_DFF_A|45|B I5|_DFF_A|T2 I5|_DFF_A|45|MID_SHUNT  3.84154647408
LI5|_DFF_A|45|RB I5|_DFF_A|45|MID_SHUNT I5|_DFF_A|A4  2.1704737578552e-12
BI5|_DFF_A|6|1 I5|_DFF_A|Q1 I5|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_A|6|P I5|_DFF_A|6|MID_SERIES 0  2e-13
RI5|_DFF_A|6|B I5|_DFF_A|Q1 I5|_DFF_A|6|MID_SHUNT  2.7439617672
LI5|_DFF_A|6|RB I5|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI5|_DFF_B|I_1|B I5|_DFF_B|A1 I5|_DFF_B|I_1|MID  2e-12
II5|_DFF_B|I_1|B 0 I5|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI5|_DFF_B|I_3|B I5|_DFF_B|A3 I5|_DFF_B|I_3|MID  2e-12
II5|_DFF_B|I_3|B 0 I5|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI5|_DFF_B|I_T|B I5|_DFF_B|T1 I5|_DFF_B|I_T|MID  2e-12
II5|_DFF_B|I_T|B 0 I5|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI5|_DFF_B|I_6|B I5|_DFF_B|Q1 I5|_DFF_B|I_6|MID  2e-12
II5|_DFF_B|I_6|B 0 I5|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI5|_DFF_B|1|1 I5|_DFF_B|A1 I5|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_B|1|P I5|_DFF_B|1|MID_SERIES 0  2e-13
RI5|_DFF_B|1|B I5|_DFF_B|A1 I5|_DFF_B|1|MID_SHUNT  2.7439617672
LI5|_DFF_B|1|RB I5|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_B|23|1 I5|_DFF_B|A2 I5|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI5|_DFF_B|23|B I5|_DFF_B|A2 I5|_DFF_B|23|MID_SHUNT  3.84154647408
LI5|_DFF_B|23|RB I5|_DFF_B|23|MID_SHUNT I5|_DFF_B|A3  2.1704737578552e-12
BI5|_DFF_B|3|1 I5|_DFF_B|A3 I5|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_B|3|P I5|_DFF_B|3|MID_SERIES 0  2e-13
RI5|_DFF_B|3|B I5|_DFF_B|A3 I5|_DFF_B|3|MID_SHUNT  2.7439617672
LI5|_DFF_B|3|RB I5|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_B|4|1 I5|_DFF_B|A4 I5|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_B|4|P I5|_DFF_B|4|MID_SERIES 0  2e-13
RI5|_DFF_B|4|B I5|_DFF_B|A4 I5|_DFF_B|4|MID_SHUNT  2.7439617672
LI5|_DFF_B|4|RB I5|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_B|T|1 I5|_DFF_B|T1 I5|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_B|T|P I5|_DFF_B|T|MID_SERIES 0  2e-13
RI5|_DFF_B|T|B I5|_DFF_B|T1 I5|_DFF_B|T|MID_SHUNT  2.7439617672
LI5|_DFF_B|T|RB I5|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI5|_DFF_B|45|1 I5|_DFF_B|T2 I5|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI5|_DFF_B|45|B I5|_DFF_B|T2 I5|_DFF_B|45|MID_SHUNT  3.84154647408
LI5|_DFF_B|45|RB I5|_DFF_B|45|MID_SHUNT I5|_DFF_B|A4  2.1704737578552e-12
BI5|_DFF_B|6|1 I5|_DFF_B|Q1 I5|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI5|_DFF_B|6|P I5|_DFF_B|6|MID_SERIES 0  2e-13
RI5|_DFF_B|6|B I5|_DFF_B|Q1 I5|_DFF_B|6|MID_SHUNT  2.7439617672
LI5|_DFF_B|6|RB I5|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI5|_XOR|I_A1|B I5|_XOR|A1 I5|_XOR|I_A1|MID  2e-12
II5|_XOR|I_A1|B 0 I5|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI5|_XOR|I_A3|B I5|_XOR|A3 I5|_XOR|I_A3|MID  2e-12
II5|_XOR|I_A3|B 0 I5|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI5|_XOR|I_B1|B I5|_XOR|B1 I5|_XOR|I_B1|MID  2e-12
II5|_XOR|I_B1|B 0 I5|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI5|_XOR|I_B3|B I5|_XOR|B3 I5|_XOR|I_B3|MID  2e-12
II5|_XOR|I_B3|B 0 I5|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI5|_XOR|I_Q1|B I5|_XOR|Q1 I5|_XOR|I_Q1|MID  2e-12
II5|_XOR|I_Q1|B 0 I5|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI5|_XOR|A1|1 I5|_XOR|A1 I5|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|A1|P I5|_XOR|A1|MID_SERIES 0  5e-13
RI5|_XOR|A1|B I5|_XOR|A1 I5|_XOR|A1|MID_SHUNT  2.7439617672
LI5|_XOR|A1|RB I5|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI5|_XOR|A2|1 I5|_XOR|A2 I5|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|A2|P I5|_XOR|A2|MID_SERIES 0  5e-13
RI5|_XOR|A2|B I5|_XOR|A2 I5|_XOR|A2|MID_SHUNT  2.7439617672
LI5|_XOR|A2|RB I5|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI5|_XOR|A3|1 I5|_XOR|A2 I5|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|A3|P I5|_XOR|A3|MID_SERIES I5|_XOR|A3  1.2e-12
RI5|_XOR|A3|B I5|_XOR|A2 I5|_XOR|A3|MID_SHUNT  2.7439617672
LI5|_XOR|A3|RB I5|_XOR|A3|MID_SHUNT I5|_XOR|A3  2.050338398468e-12
BI5|_XOR|B1|1 I5|_XOR|B1 I5|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|B1|P I5|_XOR|B1|MID_SERIES 0  5e-13
RI5|_XOR|B1|B I5|_XOR|B1 I5|_XOR|B1|MID_SHUNT  2.7439617672
LI5|_XOR|B1|RB I5|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI5|_XOR|B2|1 I5|_XOR|B2 I5|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|B2|P I5|_XOR|B2|MID_SERIES 0  5e-13
RI5|_XOR|B2|B I5|_XOR|B2 I5|_XOR|B2|MID_SHUNT  2.7439617672
LI5|_XOR|B2|RB I5|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI5|_XOR|B3|1 I5|_XOR|B2 I5|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|B3|P I5|_XOR|B3|MID_SERIES I5|_XOR|B3  1.2e-12
RI5|_XOR|B3|B I5|_XOR|B2 I5|_XOR|B3|MID_SHUNT  2.7439617672
LI5|_XOR|B3|RB I5|_XOR|B3|MID_SHUNT I5|_XOR|B3  2.050338398468e-12
BI5|_XOR|T1|1 I5|_XOR|T1 I5|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|T1|P I5|_XOR|T1|MID_SERIES 0  5e-13
RI5|_XOR|T1|B I5|_XOR|T1 I5|_XOR|T1|MID_SHUNT  2.7439617672
LI5|_XOR|T1|RB I5|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI5|_XOR|T2|1 I5|_XOR|T2 I5|_XOR|ABTQ JJMIT AREA=2.0
RI5|_XOR|T2|B I5|_XOR|T2 I5|_XOR|T2|MID_SHUNT  3.429952209
LI5|_XOR|T2|RB I5|_XOR|T2|MID_SHUNT I5|_XOR|ABTQ  2.437922998085e-12
BI5|_XOR|AB|1 I5|_XOR|AB I5|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI5|_XOR|AB|P I5|_XOR|AB|MID_SERIES I5|_XOR|ABTQ  1.2e-12
RI5|_XOR|AB|B I5|_XOR|AB I5|_XOR|AB|MID_SHUNT  3.429952209
LI5|_XOR|AB|RB I5|_XOR|AB|MID_SHUNT I5|_XOR|ABTQ  2.437922998085e-12
BI5|_XOR|ABTQ|1 I5|_XOR|ABTQ I5|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|ABTQ|P I5|_XOR|ABTQ|MID_SERIES 0  5e-13
RI5|_XOR|ABTQ|B I5|_XOR|ABTQ I5|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI5|_XOR|ABTQ|RB I5|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI5|_XOR|Q1|1 I5|_XOR|Q1 I5|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI5|_XOR|Q1|P I5|_XOR|Q1|MID_SERIES 0  5e-13
RI5|_XOR|Q1|B I5|_XOR|Q1 I5|_XOR|Q1|MID_SHUNT  2.7439617672
LI5|_XOR|Q1|RB I5|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI5|_AND|I_A1|B I5|_AND|A1 I5|_AND|I_A1|MID  2e-12
II5|_AND|I_A1|B 0 I5|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI5|_AND|I_B1|B I5|_AND|B1 I5|_AND|I_B1|MID  2e-12
II5|_AND|I_B1|B 0 I5|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI5|_AND|I_Q3|B I5|_AND|Q3 I5|_AND|I_Q3|MID  2e-12
II5|_AND|I_Q3|B 0 I5|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI5|_AND|I_Q2|B I5|_AND|Q2 I5|_AND|I_Q2|MID  2e-12
II5|_AND|I_Q2|B 0 I5|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI5|_AND|I_Q1|B I5|_AND|Q1 I5|_AND|I_Q1|MID  2e-12
II5|_AND|I_Q1|B 0 I5|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI5|_AND|A1|1 I5|_AND|A1 I5|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI5|_AND|A1|P I5|_AND|A1|MID_SERIES 0  2e-13
RI5|_AND|A1|B I5|_AND|A1 I5|_AND|A1|MID_SHUNT  2.7439617672
LI5|_AND|A1|RB I5|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI5|_AND|A2|1 I5|_AND|A2 I5|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI5|_AND|A2|P I5|_AND|A2|MID_SERIES 0  2e-13
RI5|_AND|A2|B I5|_AND|A2 I5|_AND|A2|MID_SHUNT  2.7439617672
LI5|_AND|A2|RB I5|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI5|_AND|A12|1 I5|_AND|A2 I5|_AND|A3 JJMIT AREA=1.7857142857142858
RI5|_AND|A12|B I5|_AND|A2 I5|_AND|A12|MID_SHUNT  3.84154647408
LI5|_AND|A12|RB I5|_AND|A12|MID_SHUNT I5|_AND|A3  2.1704737578552e-12
BI5|_AND|B1|1 I5|_AND|B1 I5|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI5|_AND|B1|P I5|_AND|B1|MID_SERIES 0  2e-13
RI5|_AND|B1|B I5|_AND|B1 I5|_AND|B1|MID_SHUNT  2.7439617672
LI5|_AND|B1|RB I5|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI5|_AND|B2|1 I5|_AND|B2 I5|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI5|_AND|B2|P I5|_AND|B2|MID_SERIES 0  2e-13
RI5|_AND|B2|B I5|_AND|B2 I5|_AND|B2|MID_SHUNT  2.7439617672
LI5|_AND|B2|RB I5|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI5|_AND|B12|1 I5|_AND|B2 I5|_AND|B3 JJMIT AREA=1.7857142857142858
RI5|_AND|B12|B I5|_AND|B2 I5|_AND|B12|MID_SHUNT  3.84154647408
LI5|_AND|B12|RB I5|_AND|B12|MID_SHUNT I5|_AND|B3  2.1704737578552e-12
BI5|_AND|Q2|1 I5|_AND|Q2 I5|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI5|_AND|Q2|P I5|_AND|Q2|MID_SERIES 0  2e-13
RI5|_AND|Q2|B I5|_AND|Q2 I5|_AND|Q2|MID_SHUNT  2.7439617672
LI5|_AND|Q2|RB I5|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI5|_AND|Q1|1 I5|_AND|Q1 I5|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI5|_AND|Q1|P I5|_AND|Q1|MID_SERIES 0  2e-13
RI5|_AND|Q1|B I5|_AND|Q1 I5|_AND|Q1|MID_SHUNT  2.7439617672
LI5|_AND|Q1|RB I5|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI6|_SPL_A|I_D1|B I6|_SPL_A|D1 I6|_SPL_A|I_D1|MID  2e-12
II6|_SPL_A|I_D1|B 0 I6|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI6|_SPL_A|I_D2|B I6|_SPL_A|D2 I6|_SPL_A|I_D2|MID  2e-12
II6|_SPL_A|I_D2|B 0 I6|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI6|_SPL_A|I_Q1|B I6|_SPL_A|QA1 I6|_SPL_A|I_Q1|MID  2e-12
II6|_SPL_A|I_Q1|B 0 I6|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI6|_SPL_A|I_Q2|B I6|_SPL_A|QB1 I6|_SPL_A|I_Q2|MID  2e-12
II6|_SPL_A|I_Q2|B 0 I6|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI6|_SPL_A|1|1 I6|_SPL_A|D1 I6|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_A|1|P I6|_SPL_A|1|MID_SERIES 0  2e-13
RI6|_SPL_A|1|B I6|_SPL_A|D1 I6|_SPL_A|1|MID_SHUNT  2.7439617672
LI6|_SPL_A|1|RB I6|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI6|_SPL_A|2|1 I6|_SPL_A|D2 I6|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_A|2|P I6|_SPL_A|2|MID_SERIES 0  2e-13
RI6|_SPL_A|2|B I6|_SPL_A|D2 I6|_SPL_A|2|MID_SHUNT  2.7439617672
LI6|_SPL_A|2|RB I6|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI6|_SPL_A|A|1 I6|_SPL_A|QA1 I6|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_A|A|P I6|_SPL_A|A|MID_SERIES 0  2e-13
RI6|_SPL_A|A|B I6|_SPL_A|QA1 I6|_SPL_A|A|MID_SHUNT  2.7439617672
LI6|_SPL_A|A|RB I6|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI6|_SPL_A|B|1 I6|_SPL_A|QB1 I6|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_A|B|P I6|_SPL_A|B|MID_SERIES 0  2e-13
RI6|_SPL_A|B|B I6|_SPL_A|QB1 I6|_SPL_A|B|MID_SHUNT  2.7439617672
LI6|_SPL_A|B|RB I6|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI6|_SPL_B|I_D1|B I6|_SPL_B|D1 I6|_SPL_B|I_D1|MID  2e-12
II6|_SPL_B|I_D1|B 0 I6|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI6|_SPL_B|I_D2|B I6|_SPL_B|D2 I6|_SPL_B|I_D2|MID  2e-12
II6|_SPL_B|I_D2|B 0 I6|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI6|_SPL_B|I_Q1|B I6|_SPL_B|QA1 I6|_SPL_B|I_Q1|MID  2e-12
II6|_SPL_B|I_Q1|B 0 I6|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI6|_SPL_B|I_Q2|B I6|_SPL_B|QB1 I6|_SPL_B|I_Q2|MID  2e-12
II6|_SPL_B|I_Q2|B 0 I6|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI6|_SPL_B|1|1 I6|_SPL_B|D1 I6|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_B|1|P I6|_SPL_B|1|MID_SERIES 0  2e-13
RI6|_SPL_B|1|B I6|_SPL_B|D1 I6|_SPL_B|1|MID_SHUNT  2.7439617672
LI6|_SPL_B|1|RB I6|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI6|_SPL_B|2|1 I6|_SPL_B|D2 I6|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_B|2|P I6|_SPL_B|2|MID_SERIES 0  2e-13
RI6|_SPL_B|2|B I6|_SPL_B|D2 I6|_SPL_B|2|MID_SHUNT  2.7439617672
LI6|_SPL_B|2|RB I6|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI6|_SPL_B|A|1 I6|_SPL_B|QA1 I6|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_B|A|P I6|_SPL_B|A|MID_SERIES 0  2e-13
RI6|_SPL_B|A|B I6|_SPL_B|QA1 I6|_SPL_B|A|MID_SHUNT  2.7439617672
LI6|_SPL_B|A|RB I6|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI6|_SPL_B|B|1 I6|_SPL_B|QB1 I6|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI6|_SPL_B|B|P I6|_SPL_B|B|MID_SERIES 0  2e-13
RI6|_SPL_B|B|B I6|_SPL_B|QB1 I6|_SPL_B|B|MID_SHUNT  2.7439617672
LI6|_SPL_B|B|RB I6|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI6|_DFF_A|I_1|B I6|_DFF_A|A1 I6|_DFF_A|I_1|MID  2e-12
II6|_DFF_A|I_1|B 0 I6|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI6|_DFF_A|I_3|B I6|_DFF_A|A3 I6|_DFF_A|I_3|MID  2e-12
II6|_DFF_A|I_3|B 0 I6|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI6|_DFF_A|I_T|B I6|_DFF_A|T1 I6|_DFF_A|I_T|MID  2e-12
II6|_DFF_A|I_T|B 0 I6|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI6|_DFF_A|I_6|B I6|_DFF_A|Q1 I6|_DFF_A|I_6|MID  2e-12
II6|_DFF_A|I_6|B 0 I6|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI6|_DFF_A|1|1 I6|_DFF_A|A1 I6|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_A|1|P I6|_DFF_A|1|MID_SERIES 0  2e-13
RI6|_DFF_A|1|B I6|_DFF_A|A1 I6|_DFF_A|1|MID_SHUNT  2.7439617672
LI6|_DFF_A|1|RB I6|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_A|23|1 I6|_DFF_A|A2 I6|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI6|_DFF_A|23|B I6|_DFF_A|A2 I6|_DFF_A|23|MID_SHUNT  3.84154647408
LI6|_DFF_A|23|RB I6|_DFF_A|23|MID_SHUNT I6|_DFF_A|A3  2.1704737578552e-12
BI6|_DFF_A|3|1 I6|_DFF_A|A3 I6|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_A|3|P I6|_DFF_A|3|MID_SERIES 0  2e-13
RI6|_DFF_A|3|B I6|_DFF_A|A3 I6|_DFF_A|3|MID_SHUNT  2.7439617672
LI6|_DFF_A|3|RB I6|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_A|4|1 I6|_DFF_A|A4 I6|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_A|4|P I6|_DFF_A|4|MID_SERIES 0  2e-13
RI6|_DFF_A|4|B I6|_DFF_A|A4 I6|_DFF_A|4|MID_SHUNT  2.7439617672
LI6|_DFF_A|4|RB I6|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_A|T|1 I6|_DFF_A|T1 I6|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_A|T|P I6|_DFF_A|T|MID_SERIES 0  2e-13
RI6|_DFF_A|T|B I6|_DFF_A|T1 I6|_DFF_A|T|MID_SHUNT  2.7439617672
LI6|_DFF_A|T|RB I6|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_A|45|1 I6|_DFF_A|T2 I6|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI6|_DFF_A|45|B I6|_DFF_A|T2 I6|_DFF_A|45|MID_SHUNT  3.84154647408
LI6|_DFF_A|45|RB I6|_DFF_A|45|MID_SHUNT I6|_DFF_A|A4  2.1704737578552e-12
BI6|_DFF_A|6|1 I6|_DFF_A|Q1 I6|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_A|6|P I6|_DFF_A|6|MID_SERIES 0  2e-13
RI6|_DFF_A|6|B I6|_DFF_A|Q1 I6|_DFF_A|6|MID_SHUNT  2.7439617672
LI6|_DFF_A|6|RB I6|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI6|_DFF_B|I_1|B I6|_DFF_B|A1 I6|_DFF_B|I_1|MID  2e-12
II6|_DFF_B|I_1|B 0 I6|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI6|_DFF_B|I_3|B I6|_DFF_B|A3 I6|_DFF_B|I_3|MID  2e-12
II6|_DFF_B|I_3|B 0 I6|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI6|_DFF_B|I_T|B I6|_DFF_B|T1 I6|_DFF_B|I_T|MID  2e-12
II6|_DFF_B|I_T|B 0 I6|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI6|_DFF_B|I_6|B I6|_DFF_B|Q1 I6|_DFF_B|I_6|MID  2e-12
II6|_DFF_B|I_6|B 0 I6|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI6|_DFF_B|1|1 I6|_DFF_B|A1 I6|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_B|1|P I6|_DFF_B|1|MID_SERIES 0  2e-13
RI6|_DFF_B|1|B I6|_DFF_B|A1 I6|_DFF_B|1|MID_SHUNT  2.7439617672
LI6|_DFF_B|1|RB I6|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_B|23|1 I6|_DFF_B|A2 I6|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI6|_DFF_B|23|B I6|_DFF_B|A2 I6|_DFF_B|23|MID_SHUNT  3.84154647408
LI6|_DFF_B|23|RB I6|_DFF_B|23|MID_SHUNT I6|_DFF_B|A3  2.1704737578552e-12
BI6|_DFF_B|3|1 I6|_DFF_B|A3 I6|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_B|3|P I6|_DFF_B|3|MID_SERIES 0  2e-13
RI6|_DFF_B|3|B I6|_DFF_B|A3 I6|_DFF_B|3|MID_SHUNT  2.7439617672
LI6|_DFF_B|3|RB I6|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_B|4|1 I6|_DFF_B|A4 I6|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_B|4|P I6|_DFF_B|4|MID_SERIES 0  2e-13
RI6|_DFF_B|4|B I6|_DFF_B|A4 I6|_DFF_B|4|MID_SHUNT  2.7439617672
LI6|_DFF_B|4|RB I6|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_B|T|1 I6|_DFF_B|T1 I6|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_B|T|P I6|_DFF_B|T|MID_SERIES 0  2e-13
RI6|_DFF_B|T|B I6|_DFF_B|T1 I6|_DFF_B|T|MID_SHUNT  2.7439617672
LI6|_DFF_B|T|RB I6|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI6|_DFF_B|45|1 I6|_DFF_B|T2 I6|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI6|_DFF_B|45|B I6|_DFF_B|T2 I6|_DFF_B|45|MID_SHUNT  3.84154647408
LI6|_DFF_B|45|RB I6|_DFF_B|45|MID_SHUNT I6|_DFF_B|A4  2.1704737578552e-12
BI6|_DFF_B|6|1 I6|_DFF_B|Q1 I6|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI6|_DFF_B|6|P I6|_DFF_B|6|MID_SERIES 0  2e-13
RI6|_DFF_B|6|B I6|_DFF_B|Q1 I6|_DFF_B|6|MID_SHUNT  2.7439617672
LI6|_DFF_B|6|RB I6|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI6|_XOR|I_A1|B I6|_XOR|A1 I6|_XOR|I_A1|MID  2e-12
II6|_XOR|I_A1|B 0 I6|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI6|_XOR|I_A3|B I6|_XOR|A3 I6|_XOR|I_A3|MID  2e-12
II6|_XOR|I_A3|B 0 I6|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI6|_XOR|I_B1|B I6|_XOR|B1 I6|_XOR|I_B1|MID  2e-12
II6|_XOR|I_B1|B 0 I6|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI6|_XOR|I_B3|B I6|_XOR|B3 I6|_XOR|I_B3|MID  2e-12
II6|_XOR|I_B3|B 0 I6|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI6|_XOR|I_Q1|B I6|_XOR|Q1 I6|_XOR|I_Q1|MID  2e-12
II6|_XOR|I_Q1|B 0 I6|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI6|_XOR|A1|1 I6|_XOR|A1 I6|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|A1|P I6|_XOR|A1|MID_SERIES 0  5e-13
RI6|_XOR|A1|B I6|_XOR|A1 I6|_XOR|A1|MID_SHUNT  2.7439617672
LI6|_XOR|A1|RB I6|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI6|_XOR|A2|1 I6|_XOR|A2 I6|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|A2|P I6|_XOR|A2|MID_SERIES 0  5e-13
RI6|_XOR|A2|B I6|_XOR|A2 I6|_XOR|A2|MID_SHUNT  2.7439617672
LI6|_XOR|A2|RB I6|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI6|_XOR|A3|1 I6|_XOR|A2 I6|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|A3|P I6|_XOR|A3|MID_SERIES I6|_XOR|A3  1.2e-12
RI6|_XOR|A3|B I6|_XOR|A2 I6|_XOR|A3|MID_SHUNT  2.7439617672
LI6|_XOR|A3|RB I6|_XOR|A3|MID_SHUNT I6|_XOR|A3  2.050338398468e-12
BI6|_XOR|B1|1 I6|_XOR|B1 I6|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|B1|P I6|_XOR|B1|MID_SERIES 0  5e-13
RI6|_XOR|B1|B I6|_XOR|B1 I6|_XOR|B1|MID_SHUNT  2.7439617672
LI6|_XOR|B1|RB I6|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI6|_XOR|B2|1 I6|_XOR|B2 I6|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|B2|P I6|_XOR|B2|MID_SERIES 0  5e-13
RI6|_XOR|B2|B I6|_XOR|B2 I6|_XOR|B2|MID_SHUNT  2.7439617672
LI6|_XOR|B2|RB I6|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI6|_XOR|B3|1 I6|_XOR|B2 I6|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|B3|P I6|_XOR|B3|MID_SERIES I6|_XOR|B3  1.2e-12
RI6|_XOR|B3|B I6|_XOR|B2 I6|_XOR|B3|MID_SHUNT  2.7439617672
LI6|_XOR|B3|RB I6|_XOR|B3|MID_SHUNT I6|_XOR|B3  2.050338398468e-12
BI6|_XOR|T1|1 I6|_XOR|T1 I6|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|T1|P I6|_XOR|T1|MID_SERIES 0  5e-13
RI6|_XOR|T1|B I6|_XOR|T1 I6|_XOR|T1|MID_SHUNT  2.7439617672
LI6|_XOR|T1|RB I6|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI6|_XOR|T2|1 I6|_XOR|T2 I6|_XOR|ABTQ JJMIT AREA=2.0
RI6|_XOR|T2|B I6|_XOR|T2 I6|_XOR|T2|MID_SHUNT  3.429952209
LI6|_XOR|T2|RB I6|_XOR|T2|MID_SHUNT I6|_XOR|ABTQ  2.437922998085e-12
BI6|_XOR|AB|1 I6|_XOR|AB I6|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI6|_XOR|AB|P I6|_XOR|AB|MID_SERIES I6|_XOR|ABTQ  1.2e-12
RI6|_XOR|AB|B I6|_XOR|AB I6|_XOR|AB|MID_SHUNT  3.429952209
LI6|_XOR|AB|RB I6|_XOR|AB|MID_SHUNT I6|_XOR|ABTQ  2.437922998085e-12
BI6|_XOR|ABTQ|1 I6|_XOR|ABTQ I6|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|ABTQ|P I6|_XOR|ABTQ|MID_SERIES 0  5e-13
RI6|_XOR|ABTQ|B I6|_XOR|ABTQ I6|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI6|_XOR|ABTQ|RB I6|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI6|_XOR|Q1|1 I6|_XOR|Q1 I6|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI6|_XOR|Q1|P I6|_XOR|Q1|MID_SERIES 0  5e-13
RI6|_XOR|Q1|B I6|_XOR|Q1 I6|_XOR|Q1|MID_SHUNT  2.7439617672
LI6|_XOR|Q1|RB I6|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI6|_AND|I_A1|B I6|_AND|A1 I6|_AND|I_A1|MID  2e-12
II6|_AND|I_A1|B 0 I6|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI6|_AND|I_B1|B I6|_AND|B1 I6|_AND|I_B1|MID  2e-12
II6|_AND|I_B1|B 0 I6|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI6|_AND|I_Q3|B I6|_AND|Q3 I6|_AND|I_Q3|MID  2e-12
II6|_AND|I_Q3|B 0 I6|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI6|_AND|I_Q2|B I6|_AND|Q2 I6|_AND|I_Q2|MID  2e-12
II6|_AND|I_Q2|B 0 I6|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI6|_AND|I_Q1|B I6|_AND|Q1 I6|_AND|I_Q1|MID  2e-12
II6|_AND|I_Q1|B 0 I6|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI6|_AND|A1|1 I6|_AND|A1 I6|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI6|_AND|A1|P I6|_AND|A1|MID_SERIES 0  2e-13
RI6|_AND|A1|B I6|_AND|A1 I6|_AND|A1|MID_SHUNT  2.7439617672
LI6|_AND|A1|RB I6|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI6|_AND|A2|1 I6|_AND|A2 I6|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI6|_AND|A2|P I6|_AND|A2|MID_SERIES 0  2e-13
RI6|_AND|A2|B I6|_AND|A2 I6|_AND|A2|MID_SHUNT  2.7439617672
LI6|_AND|A2|RB I6|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI6|_AND|A12|1 I6|_AND|A2 I6|_AND|A3 JJMIT AREA=1.7857142857142858
RI6|_AND|A12|B I6|_AND|A2 I6|_AND|A12|MID_SHUNT  3.84154647408
LI6|_AND|A12|RB I6|_AND|A12|MID_SHUNT I6|_AND|A3  2.1704737578552e-12
BI6|_AND|B1|1 I6|_AND|B1 I6|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI6|_AND|B1|P I6|_AND|B1|MID_SERIES 0  2e-13
RI6|_AND|B1|B I6|_AND|B1 I6|_AND|B1|MID_SHUNT  2.7439617672
LI6|_AND|B1|RB I6|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI6|_AND|B2|1 I6|_AND|B2 I6|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI6|_AND|B2|P I6|_AND|B2|MID_SERIES 0  2e-13
RI6|_AND|B2|B I6|_AND|B2 I6|_AND|B2|MID_SHUNT  2.7439617672
LI6|_AND|B2|RB I6|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI6|_AND|B12|1 I6|_AND|B2 I6|_AND|B3 JJMIT AREA=1.7857142857142858
RI6|_AND|B12|B I6|_AND|B2 I6|_AND|B12|MID_SHUNT  3.84154647408
LI6|_AND|B12|RB I6|_AND|B12|MID_SHUNT I6|_AND|B3  2.1704737578552e-12
BI6|_AND|Q2|1 I6|_AND|Q2 I6|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI6|_AND|Q2|P I6|_AND|Q2|MID_SERIES 0  2e-13
RI6|_AND|Q2|B I6|_AND|Q2 I6|_AND|Q2|MID_SHUNT  2.7439617672
LI6|_AND|Q2|RB I6|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI6|_AND|Q1|1 I6|_AND|Q1 I6|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI6|_AND|Q1|P I6|_AND|Q1|MID_SERIES 0  2e-13
RI6|_AND|Q1|B I6|_AND|Q1 I6|_AND|Q1|MID_SHUNT  2.7439617672
LI6|_AND|Q1|RB I6|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI7|_SPL_A|I_D1|B I7|_SPL_A|D1 I7|_SPL_A|I_D1|MID  2e-12
II7|_SPL_A|I_D1|B 0 I7|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI7|_SPL_A|I_D2|B I7|_SPL_A|D2 I7|_SPL_A|I_D2|MID  2e-12
II7|_SPL_A|I_D2|B 0 I7|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI7|_SPL_A|I_Q1|B I7|_SPL_A|QA1 I7|_SPL_A|I_Q1|MID  2e-12
II7|_SPL_A|I_Q1|B 0 I7|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI7|_SPL_A|I_Q2|B I7|_SPL_A|QB1 I7|_SPL_A|I_Q2|MID  2e-12
II7|_SPL_A|I_Q2|B 0 I7|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI7|_SPL_A|1|1 I7|_SPL_A|D1 I7|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_A|1|P I7|_SPL_A|1|MID_SERIES 0  2e-13
RI7|_SPL_A|1|B I7|_SPL_A|D1 I7|_SPL_A|1|MID_SHUNT  2.7439617672
LI7|_SPL_A|1|RB I7|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI7|_SPL_A|2|1 I7|_SPL_A|D2 I7|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_A|2|P I7|_SPL_A|2|MID_SERIES 0  2e-13
RI7|_SPL_A|2|B I7|_SPL_A|D2 I7|_SPL_A|2|MID_SHUNT  2.7439617672
LI7|_SPL_A|2|RB I7|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI7|_SPL_A|A|1 I7|_SPL_A|QA1 I7|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_A|A|P I7|_SPL_A|A|MID_SERIES 0  2e-13
RI7|_SPL_A|A|B I7|_SPL_A|QA1 I7|_SPL_A|A|MID_SHUNT  2.7439617672
LI7|_SPL_A|A|RB I7|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI7|_SPL_A|B|1 I7|_SPL_A|QB1 I7|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_A|B|P I7|_SPL_A|B|MID_SERIES 0  2e-13
RI7|_SPL_A|B|B I7|_SPL_A|QB1 I7|_SPL_A|B|MID_SHUNT  2.7439617672
LI7|_SPL_A|B|RB I7|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI7|_SPL_B|I_D1|B I7|_SPL_B|D1 I7|_SPL_B|I_D1|MID  2e-12
II7|_SPL_B|I_D1|B 0 I7|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI7|_SPL_B|I_D2|B I7|_SPL_B|D2 I7|_SPL_B|I_D2|MID  2e-12
II7|_SPL_B|I_D2|B 0 I7|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI7|_SPL_B|I_Q1|B I7|_SPL_B|QA1 I7|_SPL_B|I_Q1|MID  2e-12
II7|_SPL_B|I_Q1|B 0 I7|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI7|_SPL_B|I_Q2|B I7|_SPL_B|QB1 I7|_SPL_B|I_Q2|MID  2e-12
II7|_SPL_B|I_Q2|B 0 I7|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI7|_SPL_B|1|1 I7|_SPL_B|D1 I7|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_B|1|P I7|_SPL_B|1|MID_SERIES 0  2e-13
RI7|_SPL_B|1|B I7|_SPL_B|D1 I7|_SPL_B|1|MID_SHUNT  2.7439617672
LI7|_SPL_B|1|RB I7|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI7|_SPL_B|2|1 I7|_SPL_B|D2 I7|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_B|2|P I7|_SPL_B|2|MID_SERIES 0  2e-13
RI7|_SPL_B|2|B I7|_SPL_B|D2 I7|_SPL_B|2|MID_SHUNT  2.7439617672
LI7|_SPL_B|2|RB I7|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI7|_SPL_B|A|1 I7|_SPL_B|QA1 I7|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_B|A|P I7|_SPL_B|A|MID_SERIES 0  2e-13
RI7|_SPL_B|A|B I7|_SPL_B|QA1 I7|_SPL_B|A|MID_SHUNT  2.7439617672
LI7|_SPL_B|A|RB I7|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI7|_SPL_B|B|1 I7|_SPL_B|QB1 I7|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI7|_SPL_B|B|P I7|_SPL_B|B|MID_SERIES 0  2e-13
RI7|_SPL_B|B|B I7|_SPL_B|QB1 I7|_SPL_B|B|MID_SHUNT  2.7439617672
LI7|_SPL_B|B|RB I7|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI7|_DFF_A|I_1|B I7|_DFF_A|A1 I7|_DFF_A|I_1|MID  2e-12
II7|_DFF_A|I_1|B 0 I7|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI7|_DFF_A|I_3|B I7|_DFF_A|A3 I7|_DFF_A|I_3|MID  2e-12
II7|_DFF_A|I_3|B 0 I7|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI7|_DFF_A|I_T|B I7|_DFF_A|T1 I7|_DFF_A|I_T|MID  2e-12
II7|_DFF_A|I_T|B 0 I7|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI7|_DFF_A|I_6|B I7|_DFF_A|Q1 I7|_DFF_A|I_6|MID  2e-12
II7|_DFF_A|I_6|B 0 I7|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI7|_DFF_A|1|1 I7|_DFF_A|A1 I7|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_A|1|P I7|_DFF_A|1|MID_SERIES 0  2e-13
RI7|_DFF_A|1|B I7|_DFF_A|A1 I7|_DFF_A|1|MID_SHUNT  2.7439617672
LI7|_DFF_A|1|RB I7|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_A|23|1 I7|_DFF_A|A2 I7|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI7|_DFF_A|23|B I7|_DFF_A|A2 I7|_DFF_A|23|MID_SHUNT  3.84154647408
LI7|_DFF_A|23|RB I7|_DFF_A|23|MID_SHUNT I7|_DFF_A|A3  2.1704737578552e-12
BI7|_DFF_A|3|1 I7|_DFF_A|A3 I7|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_A|3|P I7|_DFF_A|3|MID_SERIES 0  2e-13
RI7|_DFF_A|3|B I7|_DFF_A|A3 I7|_DFF_A|3|MID_SHUNT  2.7439617672
LI7|_DFF_A|3|RB I7|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_A|4|1 I7|_DFF_A|A4 I7|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_A|4|P I7|_DFF_A|4|MID_SERIES 0  2e-13
RI7|_DFF_A|4|B I7|_DFF_A|A4 I7|_DFF_A|4|MID_SHUNT  2.7439617672
LI7|_DFF_A|4|RB I7|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_A|T|1 I7|_DFF_A|T1 I7|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_A|T|P I7|_DFF_A|T|MID_SERIES 0  2e-13
RI7|_DFF_A|T|B I7|_DFF_A|T1 I7|_DFF_A|T|MID_SHUNT  2.7439617672
LI7|_DFF_A|T|RB I7|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_A|45|1 I7|_DFF_A|T2 I7|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI7|_DFF_A|45|B I7|_DFF_A|T2 I7|_DFF_A|45|MID_SHUNT  3.84154647408
LI7|_DFF_A|45|RB I7|_DFF_A|45|MID_SHUNT I7|_DFF_A|A4  2.1704737578552e-12
BI7|_DFF_A|6|1 I7|_DFF_A|Q1 I7|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_A|6|P I7|_DFF_A|6|MID_SERIES 0  2e-13
RI7|_DFF_A|6|B I7|_DFF_A|Q1 I7|_DFF_A|6|MID_SHUNT  2.7439617672
LI7|_DFF_A|6|RB I7|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI7|_DFF_B|I_1|B I7|_DFF_B|A1 I7|_DFF_B|I_1|MID  2e-12
II7|_DFF_B|I_1|B 0 I7|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI7|_DFF_B|I_3|B I7|_DFF_B|A3 I7|_DFF_B|I_3|MID  2e-12
II7|_DFF_B|I_3|B 0 I7|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI7|_DFF_B|I_T|B I7|_DFF_B|T1 I7|_DFF_B|I_T|MID  2e-12
II7|_DFF_B|I_T|B 0 I7|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI7|_DFF_B|I_6|B I7|_DFF_B|Q1 I7|_DFF_B|I_6|MID  2e-12
II7|_DFF_B|I_6|B 0 I7|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI7|_DFF_B|1|1 I7|_DFF_B|A1 I7|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_B|1|P I7|_DFF_B|1|MID_SERIES 0  2e-13
RI7|_DFF_B|1|B I7|_DFF_B|A1 I7|_DFF_B|1|MID_SHUNT  2.7439617672
LI7|_DFF_B|1|RB I7|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_B|23|1 I7|_DFF_B|A2 I7|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI7|_DFF_B|23|B I7|_DFF_B|A2 I7|_DFF_B|23|MID_SHUNT  3.84154647408
LI7|_DFF_B|23|RB I7|_DFF_B|23|MID_SHUNT I7|_DFF_B|A3  2.1704737578552e-12
BI7|_DFF_B|3|1 I7|_DFF_B|A3 I7|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_B|3|P I7|_DFF_B|3|MID_SERIES 0  2e-13
RI7|_DFF_B|3|B I7|_DFF_B|A3 I7|_DFF_B|3|MID_SHUNT  2.7439617672
LI7|_DFF_B|3|RB I7|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_B|4|1 I7|_DFF_B|A4 I7|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_B|4|P I7|_DFF_B|4|MID_SERIES 0  2e-13
RI7|_DFF_B|4|B I7|_DFF_B|A4 I7|_DFF_B|4|MID_SHUNT  2.7439617672
LI7|_DFF_B|4|RB I7|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_B|T|1 I7|_DFF_B|T1 I7|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_B|T|P I7|_DFF_B|T|MID_SERIES 0  2e-13
RI7|_DFF_B|T|B I7|_DFF_B|T1 I7|_DFF_B|T|MID_SHUNT  2.7439617672
LI7|_DFF_B|T|RB I7|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI7|_DFF_B|45|1 I7|_DFF_B|T2 I7|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI7|_DFF_B|45|B I7|_DFF_B|T2 I7|_DFF_B|45|MID_SHUNT  3.84154647408
LI7|_DFF_B|45|RB I7|_DFF_B|45|MID_SHUNT I7|_DFF_B|A4  2.1704737578552e-12
BI7|_DFF_B|6|1 I7|_DFF_B|Q1 I7|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI7|_DFF_B|6|P I7|_DFF_B|6|MID_SERIES 0  2e-13
RI7|_DFF_B|6|B I7|_DFF_B|Q1 I7|_DFF_B|6|MID_SHUNT  2.7439617672
LI7|_DFF_B|6|RB I7|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI7|_XOR|I_A1|B I7|_XOR|A1 I7|_XOR|I_A1|MID  2e-12
II7|_XOR|I_A1|B 0 I7|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI7|_XOR|I_A3|B I7|_XOR|A3 I7|_XOR|I_A3|MID  2e-12
II7|_XOR|I_A3|B 0 I7|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI7|_XOR|I_B1|B I7|_XOR|B1 I7|_XOR|I_B1|MID  2e-12
II7|_XOR|I_B1|B 0 I7|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI7|_XOR|I_B3|B I7|_XOR|B3 I7|_XOR|I_B3|MID  2e-12
II7|_XOR|I_B3|B 0 I7|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI7|_XOR|I_Q1|B I7|_XOR|Q1 I7|_XOR|I_Q1|MID  2e-12
II7|_XOR|I_Q1|B 0 I7|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI7|_XOR|A1|1 I7|_XOR|A1 I7|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|A1|P I7|_XOR|A1|MID_SERIES 0  5e-13
RI7|_XOR|A1|B I7|_XOR|A1 I7|_XOR|A1|MID_SHUNT  2.7439617672
LI7|_XOR|A1|RB I7|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI7|_XOR|A2|1 I7|_XOR|A2 I7|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|A2|P I7|_XOR|A2|MID_SERIES 0  5e-13
RI7|_XOR|A2|B I7|_XOR|A2 I7|_XOR|A2|MID_SHUNT  2.7439617672
LI7|_XOR|A2|RB I7|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI7|_XOR|A3|1 I7|_XOR|A2 I7|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|A3|P I7|_XOR|A3|MID_SERIES I7|_XOR|A3  1.2e-12
RI7|_XOR|A3|B I7|_XOR|A2 I7|_XOR|A3|MID_SHUNT  2.7439617672
LI7|_XOR|A3|RB I7|_XOR|A3|MID_SHUNT I7|_XOR|A3  2.050338398468e-12
BI7|_XOR|B1|1 I7|_XOR|B1 I7|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|B1|P I7|_XOR|B1|MID_SERIES 0  5e-13
RI7|_XOR|B1|B I7|_XOR|B1 I7|_XOR|B1|MID_SHUNT  2.7439617672
LI7|_XOR|B1|RB I7|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI7|_XOR|B2|1 I7|_XOR|B2 I7|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|B2|P I7|_XOR|B2|MID_SERIES 0  5e-13
RI7|_XOR|B2|B I7|_XOR|B2 I7|_XOR|B2|MID_SHUNT  2.7439617672
LI7|_XOR|B2|RB I7|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI7|_XOR|B3|1 I7|_XOR|B2 I7|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|B3|P I7|_XOR|B3|MID_SERIES I7|_XOR|B3  1.2e-12
RI7|_XOR|B3|B I7|_XOR|B2 I7|_XOR|B3|MID_SHUNT  2.7439617672
LI7|_XOR|B3|RB I7|_XOR|B3|MID_SHUNT I7|_XOR|B3  2.050338398468e-12
BI7|_XOR|T1|1 I7|_XOR|T1 I7|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|T1|P I7|_XOR|T1|MID_SERIES 0  5e-13
RI7|_XOR|T1|B I7|_XOR|T1 I7|_XOR|T1|MID_SHUNT  2.7439617672
LI7|_XOR|T1|RB I7|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI7|_XOR|T2|1 I7|_XOR|T2 I7|_XOR|ABTQ JJMIT AREA=2.0
RI7|_XOR|T2|B I7|_XOR|T2 I7|_XOR|T2|MID_SHUNT  3.429952209
LI7|_XOR|T2|RB I7|_XOR|T2|MID_SHUNT I7|_XOR|ABTQ  2.437922998085e-12
BI7|_XOR|AB|1 I7|_XOR|AB I7|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI7|_XOR|AB|P I7|_XOR|AB|MID_SERIES I7|_XOR|ABTQ  1.2e-12
RI7|_XOR|AB|B I7|_XOR|AB I7|_XOR|AB|MID_SHUNT  3.429952209
LI7|_XOR|AB|RB I7|_XOR|AB|MID_SHUNT I7|_XOR|ABTQ  2.437922998085e-12
BI7|_XOR|ABTQ|1 I7|_XOR|ABTQ I7|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|ABTQ|P I7|_XOR|ABTQ|MID_SERIES 0  5e-13
RI7|_XOR|ABTQ|B I7|_XOR|ABTQ I7|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI7|_XOR|ABTQ|RB I7|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI7|_XOR|Q1|1 I7|_XOR|Q1 I7|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI7|_XOR|Q1|P I7|_XOR|Q1|MID_SERIES 0  5e-13
RI7|_XOR|Q1|B I7|_XOR|Q1 I7|_XOR|Q1|MID_SHUNT  2.7439617672
LI7|_XOR|Q1|RB I7|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI7|_AND|I_A1|B I7|_AND|A1 I7|_AND|I_A1|MID  2e-12
II7|_AND|I_A1|B 0 I7|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI7|_AND|I_B1|B I7|_AND|B1 I7|_AND|I_B1|MID  2e-12
II7|_AND|I_B1|B 0 I7|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI7|_AND|I_Q3|B I7|_AND|Q3 I7|_AND|I_Q3|MID  2e-12
II7|_AND|I_Q3|B 0 I7|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI7|_AND|I_Q2|B I7|_AND|Q2 I7|_AND|I_Q2|MID  2e-12
II7|_AND|I_Q2|B 0 I7|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI7|_AND|I_Q1|B I7|_AND|Q1 I7|_AND|I_Q1|MID  2e-12
II7|_AND|I_Q1|B 0 I7|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI7|_AND|A1|1 I7|_AND|A1 I7|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI7|_AND|A1|P I7|_AND|A1|MID_SERIES 0  2e-13
RI7|_AND|A1|B I7|_AND|A1 I7|_AND|A1|MID_SHUNT  2.7439617672
LI7|_AND|A1|RB I7|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI7|_AND|A2|1 I7|_AND|A2 I7|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI7|_AND|A2|P I7|_AND|A2|MID_SERIES 0  2e-13
RI7|_AND|A2|B I7|_AND|A2 I7|_AND|A2|MID_SHUNT  2.7439617672
LI7|_AND|A2|RB I7|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI7|_AND|A12|1 I7|_AND|A2 I7|_AND|A3 JJMIT AREA=1.7857142857142858
RI7|_AND|A12|B I7|_AND|A2 I7|_AND|A12|MID_SHUNT  3.84154647408
LI7|_AND|A12|RB I7|_AND|A12|MID_SHUNT I7|_AND|A3  2.1704737578552e-12
BI7|_AND|B1|1 I7|_AND|B1 I7|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI7|_AND|B1|P I7|_AND|B1|MID_SERIES 0  2e-13
RI7|_AND|B1|B I7|_AND|B1 I7|_AND|B1|MID_SHUNT  2.7439617672
LI7|_AND|B1|RB I7|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI7|_AND|B2|1 I7|_AND|B2 I7|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI7|_AND|B2|P I7|_AND|B2|MID_SERIES 0  2e-13
RI7|_AND|B2|B I7|_AND|B2 I7|_AND|B2|MID_SHUNT  2.7439617672
LI7|_AND|B2|RB I7|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI7|_AND|B12|1 I7|_AND|B2 I7|_AND|B3 JJMIT AREA=1.7857142857142858
RI7|_AND|B12|B I7|_AND|B2 I7|_AND|B12|MID_SHUNT  3.84154647408
LI7|_AND|B12|RB I7|_AND|B12|MID_SHUNT I7|_AND|B3  2.1704737578552e-12
BI7|_AND|Q2|1 I7|_AND|Q2 I7|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI7|_AND|Q2|P I7|_AND|Q2|MID_SERIES 0  2e-13
RI7|_AND|Q2|B I7|_AND|Q2 I7|_AND|Q2|MID_SHUNT  2.7439617672
LI7|_AND|Q2|RB I7|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI7|_AND|Q1|1 I7|_AND|Q1 I7|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI7|_AND|Q1|P I7|_AND|Q1|MID_SERIES 0  2e-13
RI7|_AND|Q1|B I7|_AND|Q1 I7|_AND|Q1|MID_SHUNT  2.7439617672
LI7|_AND|Q1|RB I7|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP0_0|_SPL|I_D1|B _PTL_IP0_0|_SPL|D1 _PTL_IP0_0|_SPL|I_D1|MID  2e-12
I_PTL_IP0_0|_SPL|I_D1|B 0 _PTL_IP0_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_SPL|I_D2|B _PTL_IP0_0|_SPL|D2 _PTL_IP0_0|_SPL|I_D2|MID  2e-12
I_PTL_IP0_0|_SPL|I_D2|B 0 _PTL_IP0_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP0_0|_SPL|I_Q1|B _PTL_IP0_0|_SPL|QA1 _PTL_IP0_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP0_0|_SPL|I_Q1|B 0 _PTL_IP0_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP0_0|_SPL|I_Q2|B _PTL_IP0_0|_SPL|QB1 _PTL_IP0_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP0_0|_SPL|I_Q2|B 0 _PTL_IP0_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP0_0|_SPL|1|1 _PTL_IP0_0|_SPL|D1 _PTL_IP0_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP0_0|_SPL|1|P _PTL_IP0_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP0_0|_SPL|1|B _PTL_IP0_0|_SPL|D1 _PTL_IP0_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP0_0|_SPL|1|RB _PTL_IP0_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP0_0|_SPL|2|1 _PTL_IP0_0|_SPL|D2 _PTL_IP0_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP0_0|_SPL|2|P _PTL_IP0_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP0_0|_SPL|2|B _PTL_IP0_0|_SPL|D2 _PTL_IP0_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP0_0|_SPL|2|RB _PTL_IP0_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP0_0|_SPL|A|1 _PTL_IP0_0|_SPL|QA1 _PTL_IP0_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP0_0|_SPL|A|P _PTL_IP0_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP0_0|_SPL|A|B _PTL_IP0_0|_SPL|QA1 _PTL_IP0_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP0_0|_SPL|A|RB _PTL_IP0_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP0_0|_SPL|B|1 _PTL_IP0_0|_SPL|QB1 _PTL_IP0_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP0_0|_SPL|B|P _PTL_IP0_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP0_0|_SPL|B|B _PTL_IP0_0|_SPL|QB1 _PTL_IP0_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP0_0|_SPL|B|RB _PTL_IP0_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IG0_0|_SPL|I_D1|B _PTL_IG0_0|_SPL|D1 _PTL_IG0_0|_SPL|I_D1|MID  2e-12
I_PTL_IG0_0|_SPL|I_D1|B 0 _PTL_IG0_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_SPL|I_D2|B _PTL_IG0_0|_SPL|D2 _PTL_IG0_0|_SPL|I_D2|MID  2e-12
I_PTL_IG0_0|_SPL|I_D2|B 0 _PTL_IG0_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IG0_0|_SPL|I_Q1|B _PTL_IG0_0|_SPL|QA1 _PTL_IG0_0|_SPL|I_Q1|MID  2e-12
I_PTL_IG0_0|_SPL|I_Q1|B 0 _PTL_IG0_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG0_0|_SPL|I_Q2|B _PTL_IG0_0|_SPL|QB1 _PTL_IG0_0|_SPL|I_Q2|MID  2e-12
I_PTL_IG0_0|_SPL|I_Q2|B 0 _PTL_IG0_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IG0_0|_SPL|1|1 _PTL_IG0_0|_SPL|D1 _PTL_IG0_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IG0_0|_SPL|1|P _PTL_IG0_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IG0_0|_SPL|1|B _PTL_IG0_0|_SPL|D1 _PTL_IG0_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IG0_0|_SPL|1|RB _PTL_IG0_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG0_0|_SPL|2|1 _PTL_IG0_0|_SPL|D2 _PTL_IG0_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IG0_0|_SPL|2|P _PTL_IG0_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IG0_0|_SPL|2|B _PTL_IG0_0|_SPL|D2 _PTL_IG0_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IG0_0|_SPL|2|RB _PTL_IG0_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG0_0|_SPL|A|1 _PTL_IG0_0|_SPL|QA1 _PTL_IG0_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IG0_0|_SPL|A|P _PTL_IG0_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IG0_0|_SPL|A|B _PTL_IG0_0|_SPL|QA1 _PTL_IG0_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IG0_0|_SPL|A|RB _PTL_IG0_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG0_0|_SPL|B|1 _PTL_IG0_0|_SPL|QB1 _PTL_IG0_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IG0_0|_SPL|B|P _PTL_IG0_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IG0_0|_SPL|B|B _PTL_IG0_0|_SPL|QB1 _PTL_IG0_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IG0_0|_SPL|B|RB _PTL_IG0_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP1_0|_SPL|I_D1|B _PTL_IP1_0|_SPL|D1 _PTL_IP1_0|_SPL|I_D1|MID  2e-12
I_PTL_IP1_0|_SPL|I_D1|B 0 _PTL_IP1_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_SPL|I_D2|B _PTL_IP1_0|_SPL|D2 _PTL_IP1_0|_SPL|I_D2|MID  2e-12
I_PTL_IP1_0|_SPL|I_D2|B 0 _PTL_IP1_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP1_0|_SPL|I_Q1|B _PTL_IP1_0|_SPL|QA1 _PTL_IP1_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP1_0|_SPL|I_Q1|B 0 _PTL_IP1_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP1_0|_SPL|I_Q2|B _PTL_IP1_0|_SPL|QB1 _PTL_IP1_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP1_0|_SPL|I_Q2|B 0 _PTL_IP1_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP1_0|_SPL|1|1 _PTL_IP1_0|_SPL|D1 _PTL_IP1_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP1_0|_SPL|1|P _PTL_IP1_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP1_0|_SPL|1|B _PTL_IP1_0|_SPL|D1 _PTL_IP1_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP1_0|_SPL|1|RB _PTL_IP1_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP1_0|_SPL|2|1 _PTL_IP1_0|_SPL|D2 _PTL_IP1_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP1_0|_SPL|2|P _PTL_IP1_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP1_0|_SPL|2|B _PTL_IP1_0|_SPL|D2 _PTL_IP1_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP1_0|_SPL|2|RB _PTL_IP1_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP1_0|_SPL|A|1 _PTL_IP1_0|_SPL|QA1 _PTL_IP1_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP1_0|_SPL|A|P _PTL_IP1_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP1_0|_SPL|A|B _PTL_IP1_0|_SPL|QA1 _PTL_IP1_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP1_0|_SPL|A|RB _PTL_IP1_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP1_0|_SPL|B|1 _PTL_IP1_0|_SPL|QB1 _PTL_IP1_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP1_0|_SPL|B|P _PTL_IP1_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP1_0|_SPL|B|B _PTL_IP1_0|_SPL|QB1 _PTL_IP1_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP1_0|_SPL|B|RB _PTL_IP1_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP2_0|_SPL|I_D1|B _PTL_IP2_0|_SPL|D1 _PTL_IP2_0|_SPL|I_D1|MID  2e-12
I_PTL_IP2_0|_SPL|I_D1|B 0 _PTL_IP2_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_SPL|I_D2|B _PTL_IP2_0|_SPL|D2 _PTL_IP2_0|_SPL|I_D2|MID  2e-12
I_PTL_IP2_0|_SPL|I_D2|B 0 _PTL_IP2_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP2_0|_SPL|I_Q1|B _PTL_IP2_0|_SPL|QA1 _PTL_IP2_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP2_0|_SPL|I_Q1|B 0 _PTL_IP2_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP2_0|_SPL|I_Q2|B _PTL_IP2_0|_SPL|QB1 _PTL_IP2_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP2_0|_SPL|I_Q2|B 0 _PTL_IP2_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP2_0|_SPL|1|1 _PTL_IP2_0|_SPL|D1 _PTL_IP2_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP2_0|_SPL|1|P _PTL_IP2_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP2_0|_SPL|1|B _PTL_IP2_0|_SPL|D1 _PTL_IP2_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP2_0|_SPL|1|RB _PTL_IP2_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP2_0|_SPL|2|1 _PTL_IP2_0|_SPL|D2 _PTL_IP2_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP2_0|_SPL|2|P _PTL_IP2_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP2_0|_SPL|2|B _PTL_IP2_0|_SPL|D2 _PTL_IP2_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP2_0|_SPL|2|RB _PTL_IP2_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP2_0|_SPL|A|1 _PTL_IP2_0|_SPL|QA1 _PTL_IP2_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP2_0|_SPL|A|P _PTL_IP2_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP2_0|_SPL|A|B _PTL_IP2_0|_SPL|QA1 _PTL_IP2_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP2_0|_SPL|A|RB _PTL_IP2_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP2_0|_SPL|B|1 _PTL_IP2_0|_SPL|QB1 _PTL_IP2_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP2_0|_SPL|B|P _PTL_IP2_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP2_0|_SPL|B|B _PTL_IP2_0|_SPL|QB1 _PTL_IP2_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP2_0|_SPL|B|RB _PTL_IP2_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IG2_0|_SPL|I_D1|B _PTL_IG2_0|_SPL|D1 _PTL_IG2_0|_SPL|I_D1|MID  2e-12
I_PTL_IG2_0|_SPL|I_D1|B 0 _PTL_IG2_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_SPL|I_D2|B _PTL_IG2_0|_SPL|D2 _PTL_IG2_0|_SPL|I_D2|MID  2e-12
I_PTL_IG2_0|_SPL|I_D2|B 0 _PTL_IG2_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IG2_0|_SPL|I_Q1|B _PTL_IG2_0|_SPL|QA1 _PTL_IG2_0|_SPL|I_Q1|MID  2e-12
I_PTL_IG2_0|_SPL|I_Q1|B 0 _PTL_IG2_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG2_0|_SPL|I_Q2|B _PTL_IG2_0|_SPL|QB1 _PTL_IG2_0|_SPL|I_Q2|MID  2e-12
I_PTL_IG2_0|_SPL|I_Q2|B 0 _PTL_IG2_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IG2_0|_SPL|1|1 _PTL_IG2_0|_SPL|D1 _PTL_IG2_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IG2_0|_SPL|1|P _PTL_IG2_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IG2_0|_SPL|1|B _PTL_IG2_0|_SPL|D1 _PTL_IG2_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IG2_0|_SPL|1|RB _PTL_IG2_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG2_0|_SPL|2|1 _PTL_IG2_0|_SPL|D2 _PTL_IG2_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IG2_0|_SPL|2|P _PTL_IG2_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IG2_0|_SPL|2|B _PTL_IG2_0|_SPL|D2 _PTL_IG2_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IG2_0|_SPL|2|RB _PTL_IG2_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG2_0|_SPL|A|1 _PTL_IG2_0|_SPL|QA1 _PTL_IG2_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IG2_0|_SPL|A|P _PTL_IG2_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IG2_0|_SPL|A|B _PTL_IG2_0|_SPL|QA1 _PTL_IG2_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IG2_0|_SPL|A|RB _PTL_IG2_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG2_0|_SPL|B|1 _PTL_IG2_0|_SPL|QB1 _PTL_IG2_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IG2_0|_SPL|B|P _PTL_IG2_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IG2_0|_SPL|B|B _PTL_IG2_0|_SPL|QB1 _PTL_IG2_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IG2_0|_SPL|B|RB _PTL_IG2_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP3_0|_SPL|I_D1|B _PTL_IP3_0|_SPL|D1 _PTL_IP3_0|_SPL|I_D1|MID  2e-12
I_PTL_IP3_0|_SPL|I_D1|B 0 _PTL_IP3_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_SPL|I_D2|B _PTL_IP3_0|_SPL|D2 _PTL_IP3_0|_SPL|I_D2|MID  2e-12
I_PTL_IP3_0|_SPL|I_D2|B 0 _PTL_IP3_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP3_0|_SPL|I_Q1|B _PTL_IP3_0|_SPL|QA1 _PTL_IP3_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP3_0|_SPL|I_Q1|B 0 _PTL_IP3_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP3_0|_SPL|I_Q2|B _PTL_IP3_0|_SPL|QB1 _PTL_IP3_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP3_0|_SPL|I_Q2|B 0 _PTL_IP3_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP3_0|_SPL|1|1 _PTL_IP3_0|_SPL|D1 _PTL_IP3_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP3_0|_SPL|1|P _PTL_IP3_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP3_0|_SPL|1|B _PTL_IP3_0|_SPL|D1 _PTL_IP3_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP3_0|_SPL|1|RB _PTL_IP3_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP3_0|_SPL|2|1 _PTL_IP3_0|_SPL|D2 _PTL_IP3_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP3_0|_SPL|2|P _PTL_IP3_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP3_0|_SPL|2|B _PTL_IP3_0|_SPL|D2 _PTL_IP3_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP3_0|_SPL|2|RB _PTL_IP3_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP3_0|_SPL|A|1 _PTL_IP3_0|_SPL|QA1 _PTL_IP3_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP3_0|_SPL|A|P _PTL_IP3_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP3_0|_SPL|A|B _PTL_IP3_0|_SPL|QA1 _PTL_IP3_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP3_0|_SPL|A|RB _PTL_IP3_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP3_0|_SPL|B|1 _PTL_IP3_0|_SPL|QB1 _PTL_IP3_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP3_0|_SPL|B|P _PTL_IP3_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP3_0|_SPL|B|B _PTL_IP3_0|_SPL|QB1 _PTL_IP3_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP3_0|_SPL|B|RB _PTL_IP3_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP4_0|_SPL|I_D1|B _PTL_IP4_0|_SPL|D1 _PTL_IP4_0|_SPL|I_D1|MID  2e-12
I_PTL_IP4_0|_SPL|I_D1|B 0 _PTL_IP4_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP4_0|_SPL|I_D2|B _PTL_IP4_0|_SPL|D2 _PTL_IP4_0|_SPL|I_D2|MID  2e-12
I_PTL_IP4_0|_SPL|I_D2|B 0 _PTL_IP4_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP4_0|_SPL|I_Q1|B _PTL_IP4_0|_SPL|QA1 _PTL_IP4_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP4_0|_SPL|I_Q1|B 0 _PTL_IP4_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP4_0|_SPL|I_Q2|B _PTL_IP4_0|_SPL|QB1 _PTL_IP4_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP4_0|_SPL|I_Q2|B 0 _PTL_IP4_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP4_0|_SPL|1|1 _PTL_IP4_0|_SPL|D1 _PTL_IP4_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP4_0|_SPL|1|P _PTL_IP4_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP4_0|_SPL|1|B _PTL_IP4_0|_SPL|D1 _PTL_IP4_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP4_0|_SPL|1|RB _PTL_IP4_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP4_0|_SPL|2|1 _PTL_IP4_0|_SPL|D2 _PTL_IP4_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP4_0|_SPL|2|P _PTL_IP4_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP4_0|_SPL|2|B _PTL_IP4_0|_SPL|D2 _PTL_IP4_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP4_0|_SPL|2|RB _PTL_IP4_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP4_0|_SPL|A|1 _PTL_IP4_0|_SPL|QA1 _PTL_IP4_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP4_0|_SPL|A|P _PTL_IP4_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP4_0|_SPL|A|B _PTL_IP4_0|_SPL|QA1 _PTL_IP4_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP4_0|_SPL|A|RB _PTL_IP4_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP4_0|_SPL|B|1 _PTL_IP4_0|_SPL|QB1 _PTL_IP4_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP4_0|_SPL|B|P _PTL_IP4_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP4_0|_SPL|B|B _PTL_IP4_0|_SPL|QB1 _PTL_IP4_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP4_0|_SPL|B|RB _PTL_IP4_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IG4_0|_SPL|I_D1|B _PTL_IG4_0|_SPL|D1 _PTL_IG4_0|_SPL|I_D1|MID  2e-12
I_PTL_IG4_0|_SPL|I_D1|B 0 _PTL_IG4_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG4_0|_SPL|I_D2|B _PTL_IG4_0|_SPL|D2 _PTL_IG4_0|_SPL|I_D2|MID  2e-12
I_PTL_IG4_0|_SPL|I_D2|B 0 _PTL_IG4_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IG4_0|_SPL|I_Q1|B _PTL_IG4_0|_SPL|QA1 _PTL_IG4_0|_SPL|I_Q1|MID  2e-12
I_PTL_IG4_0|_SPL|I_Q1|B 0 _PTL_IG4_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG4_0|_SPL|I_Q2|B _PTL_IG4_0|_SPL|QB1 _PTL_IG4_0|_SPL|I_Q2|MID  2e-12
I_PTL_IG4_0|_SPL|I_Q2|B 0 _PTL_IG4_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IG4_0|_SPL|1|1 _PTL_IG4_0|_SPL|D1 _PTL_IG4_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IG4_0|_SPL|1|P _PTL_IG4_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IG4_0|_SPL|1|B _PTL_IG4_0|_SPL|D1 _PTL_IG4_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IG4_0|_SPL|1|RB _PTL_IG4_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG4_0|_SPL|2|1 _PTL_IG4_0|_SPL|D2 _PTL_IG4_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IG4_0|_SPL|2|P _PTL_IG4_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IG4_0|_SPL|2|B _PTL_IG4_0|_SPL|D2 _PTL_IG4_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IG4_0|_SPL|2|RB _PTL_IG4_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG4_0|_SPL|A|1 _PTL_IG4_0|_SPL|QA1 _PTL_IG4_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IG4_0|_SPL|A|P _PTL_IG4_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IG4_0|_SPL|A|B _PTL_IG4_0|_SPL|QA1 _PTL_IG4_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IG4_0|_SPL|A|RB _PTL_IG4_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG4_0|_SPL|B|1 _PTL_IG4_0|_SPL|QB1 _PTL_IG4_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IG4_0|_SPL|B|P _PTL_IG4_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IG4_0|_SPL|B|B _PTL_IG4_0|_SPL|QB1 _PTL_IG4_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IG4_0|_SPL|B|RB _PTL_IG4_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP5_0|_SPL|I_D1|B _PTL_IP5_0|_SPL|D1 _PTL_IP5_0|_SPL|I_D1|MID  2e-12
I_PTL_IP5_0|_SPL|I_D1|B 0 _PTL_IP5_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_0|_SPL|I_D2|B _PTL_IP5_0|_SPL|D2 _PTL_IP5_0|_SPL|I_D2|MID  2e-12
I_PTL_IP5_0|_SPL|I_D2|B 0 _PTL_IP5_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP5_0|_SPL|I_Q1|B _PTL_IP5_0|_SPL|QA1 _PTL_IP5_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP5_0|_SPL|I_Q1|B 0 _PTL_IP5_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP5_0|_SPL|I_Q2|B _PTL_IP5_0|_SPL|QB1 _PTL_IP5_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP5_0|_SPL|I_Q2|B 0 _PTL_IP5_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP5_0|_SPL|1|1 _PTL_IP5_0|_SPL|D1 _PTL_IP5_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP5_0|_SPL|1|P _PTL_IP5_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP5_0|_SPL|1|B _PTL_IP5_0|_SPL|D1 _PTL_IP5_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP5_0|_SPL|1|RB _PTL_IP5_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP5_0|_SPL|2|1 _PTL_IP5_0|_SPL|D2 _PTL_IP5_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP5_0|_SPL|2|P _PTL_IP5_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP5_0|_SPL|2|B _PTL_IP5_0|_SPL|D2 _PTL_IP5_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP5_0|_SPL|2|RB _PTL_IP5_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP5_0|_SPL|A|1 _PTL_IP5_0|_SPL|QA1 _PTL_IP5_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP5_0|_SPL|A|P _PTL_IP5_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP5_0|_SPL|A|B _PTL_IP5_0|_SPL|QA1 _PTL_IP5_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP5_0|_SPL|A|RB _PTL_IP5_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP5_0|_SPL|B|1 _PTL_IP5_0|_SPL|QB1 _PTL_IP5_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP5_0|_SPL|B|P _PTL_IP5_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP5_0|_SPL|B|B _PTL_IP5_0|_SPL|QB1 _PTL_IP5_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP5_0|_SPL|B|RB _PTL_IP5_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP6_0|_SPL|I_D1|B _PTL_IP6_0|_SPL|D1 _PTL_IP6_0|_SPL|I_D1|MID  2e-12
I_PTL_IP6_0|_SPL|I_D1|B 0 _PTL_IP6_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP6_0|_SPL|I_D2|B _PTL_IP6_0|_SPL|D2 _PTL_IP6_0|_SPL|I_D2|MID  2e-12
I_PTL_IP6_0|_SPL|I_D2|B 0 _PTL_IP6_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP6_0|_SPL|I_Q1|B _PTL_IP6_0|_SPL|QA1 _PTL_IP6_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP6_0|_SPL|I_Q1|B 0 _PTL_IP6_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP6_0|_SPL|I_Q2|B _PTL_IP6_0|_SPL|QB1 _PTL_IP6_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP6_0|_SPL|I_Q2|B 0 _PTL_IP6_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP6_0|_SPL|1|1 _PTL_IP6_0|_SPL|D1 _PTL_IP6_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP6_0|_SPL|1|P _PTL_IP6_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP6_0|_SPL|1|B _PTL_IP6_0|_SPL|D1 _PTL_IP6_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP6_0|_SPL|1|RB _PTL_IP6_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP6_0|_SPL|2|1 _PTL_IP6_0|_SPL|D2 _PTL_IP6_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP6_0|_SPL|2|P _PTL_IP6_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP6_0|_SPL|2|B _PTL_IP6_0|_SPL|D2 _PTL_IP6_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP6_0|_SPL|2|RB _PTL_IP6_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP6_0|_SPL|A|1 _PTL_IP6_0|_SPL|QA1 _PTL_IP6_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP6_0|_SPL|A|P _PTL_IP6_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP6_0|_SPL|A|B _PTL_IP6_0|_SPL|QA1 _PTL_IP6_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP6_0|_SPL|A|RB _PTL_IP6_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP6_0|_SPL|B|1 _PTL_IP6_0|_SPL|QB1 _PTL_IP6_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP6_0|_SPL|B|P _PTL_IP6_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP6_0|_SPL|B|B _PTL_IP6_0|_SPL|QB1 _PTL_IP6_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP6_0|_SPL|B|RB _PTL_IP6_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IG6_0|_SPL|I_D1|B _PTL_IG6_0|_SPL|D1 _PTL_IG6_0|_SPL|I_D1|MID  2e-12
I_PTL_IG6_0|_SPL|I_D1|B 0 _PTL_IG6_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG6_0|_SPL|I_D2|B _PTL_IG6_0|_SPL|D2 _PTL_IG6_0|_SPL|I_D2|MID  2e-12
I_PTL_IG6_0|_SPL|I_D2|B 0 _PTL_IG6_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IG6_0|_SPL|I_Q1|B _PTL_IG6_0|_SPL|QA1 _PTL_IG6_0|_SPL|I_Q1|MID  2e-12
I_PTL_IG6_0|_SPL|I_Q1|B 0 _PTL_IG6_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IG6_0|_SPL|I_Q2|B _PTL_IG6_0|_SPL|QB1 _PTL_IG6_0|_SPL|I_Q2|MID  2e-12
I_PTL_IG6_0|_SPL|I_Q2|B 0 _PTL_IG6_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IG6_0|_SPL|1|1 _PTL_IG6_0|_SPL|D1 _PTL_IG6_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IG6_0|_SPL|1|P _PTL_IG6_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IG6_0|_SPL|1|B _PTL_IG6_0|_SPL|D1 _PTL_IG6_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IG6_0|_SPL|1|RB _PTL_IG6_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG6_0|_SPL|2|1 _PTL_IG6_0|_SPL|D2 _PTL_IG6_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IG6_0|_SPL|2|P _PTL_IG6_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IG6_0|_SPL|2|B _PTL_IG6_0|_SPL|D2 _PTL_IG6_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IG6_0|_SPL|2|RB _PTL_IG6_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG6_0|_SPL|A|1 _PTL_IG6_0|_SPL|QA1 _PTL_IG6_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IG6_0|_SPL|A|P _PTL_IG6_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IG6_0|_SPL|A|B _PTL_IG6_0|_SPL|QA1 _PTL_IG6_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IG6_0|_SPL|A|RB _PTL_IG6_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IG6_0|_SPL|B|1 _PTL_IG6_0|_SPL|QB1 _PTL_IG6_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IG6_0|_SPL|B|P _PTL_IG6_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IG6_0|_SPL|B|B _PTL_IG6_0|_SPL|QB1 _PTL_IG6_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IG6_0|_SPL|B|RB _PTL_IG6_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_IP7_0|_SPL|I_D1|B _PTL_IP7_0|_SPL|D1 _PTL_IP7_0|_SPL|I_D1|MID  2e-12
I_PTL_IP7_0|_SPL|I_D1|B 0 _PTL_IP7_0|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_0|_SPL|I_D2|B _PTL_IP7_0|_SPL|D2 _PTL_IP7_0|_SPL|I_D2|MID  2e-12
I_PTL_IP7_0|_SPL|I_D2|B 0 _PTL_IP7_0|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_IP7_0|_SPL|I_Q1|B _PTL_IP7_0|_SPL|QA1 _PTL_IP7_0|_SPL|I_Q1|MID  2e-12
I_PTL_IP7_0|_SPL|I_Q1|B 0 _PTL_IP7_0|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_IP7_0|_SPL|I_Q2|B _PTL_IP7_0|_SPL|QB1 _PTL_IP7_0|_SPL|I_Q2|MID  2e-12
I_PTL_IP7_0|_SPL|I_Q2|B 0 _PTL_IP7_0|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_IP7_0|_SPL|1|1 _PTL_IP7_0|_SPL|D1 _PTL_IP7_0|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_IP7_0|_SPL|1|P _PTL_IP7_0|_SPL|1|MID_SERIES 0  2e-13
R_PTL_IP7_0|_SPL|1|B _PTL_IP7_0|_SPL|D1 _PTL_IP7_0|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_IP7_0|_SPL|1|RB _PTL_IP7_0|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP7_0|_SPL|2|1 _PTL_IP7_0|_SPL|D2 _PTL_IP7_0|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_IP7_0|_SPL|2|P _PTL_IP7_0|_SPL|2|MID_SERIES 0  2e-13
R_PTL_IP7_0|_SPL|2|B _PTL_IP7_0|_SPL|D2 _PTL_IP7_0|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_IP7_0|_SPL|2|RB _PTL_IP7_0|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP7_0|_SPL|A|1 _PTL_IP7_0|_SPL|QA1 _PTL_IP7_0|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_IP7_0|_SPL|A|P _PTL_IP7_0|_SPL|A|MID_SERIES 0  2e-13
R_PTL_IP7_0|_SPL|A|B _PTL_IP7_0|_SPL|QA1 _PTL_IP7_0|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_IP7_0|_SPL|A|RB _PTL_IP7_0|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_IP7_0|_SPL|B|1 _PTL_IP7_0|_SPL|QB1 _PTL_IP7_0|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_IP7_0|_SPL|B|P _PTL_IP7_0|_SPL|B|MID_SERIES 0  2e-13
R_PTL_IP7_0|_SPL|B|B _PTL_IP7_0|_SPL|QB1 _PTL_IP7_0|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_IP7_0|_SPL|B|RB _PTL_IP7_0|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_SPL_G1|I_D1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|I_D1|MID  2e-12
I_PG1_01|_SPL_G1|I_D1|B 0 _PG1_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_D2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|I_D2|MID  2e-12
I_PG1_01|_SPL_G1|I_D2|B 0 _PG1_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG1_01|_SPL_G1|I_Q1|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|I_Q1|MID  2e-12
I_PG1_01|_SPL_G1|I_Q1|B 0 _PG1_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_Q2|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|I_Q2|MID  2e-12
I_PG1_01|_SPL_G1|I_Q2|B 0 _PG1_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG1_01|_SPL_G1|1|1 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|1|P _PG1_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|1|RB _PG1_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|2|1 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|2|P _PG1_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|2|RB _PG1_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|A|1 _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|A|P _PG1_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|A|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|A|RB _PG1_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|B|1 _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|B|P _PG1_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|B|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|B|RB _PG1_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_SPL_P1|I_D1|B _PG1_01|_SPL_P1|D1 _PG1_01|_SPL_P1|I_D1|MID  2e-12
I_PG1_01|_SPL_P1|I_D1|B 0 _PG1_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_P1|I_D2|B _PG1_01|_SPL_P1|D2 _PG1_01|_SPL_P1|I_D2|MID  2e-12
I_PG1_01|_SPL_P1|I_D2|B 0 _PG1_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG1_01|_SPL_P1|I_Q1|B _PG1_01|_SPL_P1|QA1 _PG1_01|_SPL_P1|I_Q1|MID  2e-12
I_PG1_01|_SPL_P1|I_Q1|B 0 _PG1_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_P1|I_Q2|B _PG1_01|_SPL_P1|QB1 _PG1_01|_SPL_P1|I_Q2|MID  2e-12
I_PG1_01|_SPL_P1|I_Q2|B 0 _PG1_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG1_01|_SPL_P1|1|1 _PG1_01|_SPL_P1|D1 _PG1_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_P1|1|P _PG1_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG1_01|_SPL_P1|1|B _PG1_01|_SPL_P1|D1 _PG1_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_P1|1|RB _PG1_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_P1|2|1 _PG1_01|_SPL_P1|D2 _PG1_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_P1|2|P _PG1_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG1_01|_SPL_P1|2|B _PG1_01|_SPL_P1|D2 _PG1_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_P1|2|RB _PG1_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_P1|A|1 _PG1_01|_SPL_P1|QA1 _PG1_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_P1|A|P _PG1_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG1_01|_SPL_P1|A|B _PG1_01|_SPL_P1|QA1 _PG1_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_P1|A|RB _PG1_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_P1|B|1 _PG1_01|_SPL_P1|QB1 _PG1_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_P1|B|P _PG1_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG1_01|_SPL_P1|B|B _PG1_01|_SPL_P1|QB1 _PG1_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_P1|B|RB _PG1_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_PG|I_A1|B _PG1_01|_PG|A1 _PG1_01|_PG|I_A1|MID  2e-12
I_PG1_01|_PG|I_A1|B 0 _PG1_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_B1|B _PG1_01|_PG|B1 _PG1_01|_PG|I_B1|MID  2e-12
I_PG1_01|_PG|I_B1|B 0 _PG1_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q3|B _PG1_01|_PG|Q3 _PG1_01|_PG|I_Q3|MID  2e-12
I_PG1_01|_PG|I_Q3|B 0 _PG1_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_PG|I_Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|I_Q2|MID  2e-12
I_PG1_01|_PG|I_Q2|B 0 _PG1_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|I_Q1|MID  2e-12
I_PG1_01|_PG|I_Q1|B 0 _PG1_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_PG|A1|1 _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A1|P _PG1_01|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01|_PG|A1|B _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A1|RB _PG1_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A2|1 _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A2|P _PG1_01|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01|_PG|A2|B _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A2|RB _PG1_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A12|1 _PG1_01|_PG|A2 _PG1_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|A12|B _PG1_01|_PG|A2 _PG1_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|A12|RB _PG1_01|_PG|A12|MID_SHUNT _PG1_01|_PG|A3  2.1704737578552e-12
B_PG1_01|_PG|B1|1 _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B1|P _PG1_01|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01|_PG|B1|B _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B1|RB _PG1_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B2|1 _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B2|P _PG1_01|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01|_PG|B2|B _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B2|RB _PG1_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B12|1 _PG1_01|_PG|B2 _PG1_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|B12|B _PG1_01|_PG|B2 _PG1_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|B12|RB _PG1_01|_PG|B12|MID_SHUNT _PG1_01|_PG|B3  2.1704737578552e-12
B_PG1_01|_PG|Q2|1 _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q2|P _PG1_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q2|RB _PG1_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|Q1|1 _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q1|P _PG1_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q1|RB _PG1_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_GG|I_A1|B _PG1_01|_GG|A1 _PG1_01|_GG|I_A1|MID  2e-12
I_PG1_01|_GG|I_A1|B 0 _PG1_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_B1|B _PG1_01|_GG|B1 _PG1_01|_GG|I_B1|MID  2e-12
I_PG1_01|_GG|I_B1|B 0 _PG1_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q3|B _PG1_01|_GG|Q3 _PG1_01|_GG|I_Q3|MID  2e-12
I_PG1_01|_GG|I_Q3|B 0 _PG1_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_GG|I_Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|I_Q2|MID  2e-12
I_PG1_01|_GG|I_Q2|B 0 _PG1_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|I_Q1|MID  2e-12
I_PG1_01|_GG|I_Q1|B 0 _PG1_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_GG|A1|1 _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A1|P _PG1_01|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01|_GG|A1|B _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A1|RB _PG1_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A2|1 _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A2|P _PG1_01|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01|_GG|A2|B _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A2|RB _PG1_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A12|1 _PG1_01|_GG|A2 _PG1_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|A12|B _PG1_01|_GG|A2 _PG1_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|A12|RB _PG1_01|_GG|A12|MID_SHUNT _PG1_01|_GG|A3  2.1704737578552e-12
B_PG1_01|_GG|B1|1 _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B1|P _PG1_01|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01|_GG|B1|B _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B1|RB _PG1_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B2|1 _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B2|P _PG1_01|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01|_GG|B2|B _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B2|RB _PG1_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B12|1 _PG1_01|_GG|B2 _PG1_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|B12|B _PG1_01|_GG|B2 _PG1_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|B12|RB _PG1_01|_GG|B12|MID_SHUNT _PG1_01|_GG|B3  2.1704737578552e-12
B_PG1_01|_GG|Q2|1 _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q2|P _PG1_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q2|RB _PG1_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|Q1|1 _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q1|P _PG1_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q1|RB _PG1_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_P0|I_1|B _PG1_01|_DFF_P0|A1 _PG1_01|_DFF_P0|I_1|MID  2e-12
I_PG1_01|_DFF_P0|I_1|B 0 _PG1_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_P0|I_3|B _PG1_01|_DFF_P0|A3 _PG1_01|_DFF_P0|I_3|MID  2e-12
I_PG1_01|_DFF_P0|I_3|B 0 _PG1_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_P0|I_T|B _PG1_01|_DFF_P0|T1 _PG1_01|_DFF_P0|I_T|MID  2e-12
I_PG1_01|_DFF_P0|I_T|B 0 _PG1_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_P0|I_6|B _PG1_01|_DFF_P0|Q1 _PG1_01|_DFF_P0|I_6|MID  2e-12
I_PG1_01|_DFF_P0|I_6|B 0 _PG1_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_P0|1|1 _PG1_01|_DFF_P0|A1 _PG1_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P0|1|P _PG1_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P0|1|B _PG1_01|_DFF_P0|A1 _PG1_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P0|1|RB _PG1_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P0|23|1 _PG1_01|_DFF_P0|A2 _PG1_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_P0|23|B _PG1_01|_DFF_P0|A2 _PG1_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_P0|23|RB _PG1_01|_DFF_P0|23|MID_SHUNT _PG1_01|_DFF_P0|A3  2.1704737578552e-12
B_PG1_01|_DFF_P0|3|1 _PG1_01|_DFF_P0|A3 _PG1_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P0|3|P _PG1_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P0|3|B _PG1_01|_DFF_P0|A3 _PG1_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P0|3|RB _PG1_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P0|4|1 _PG1_01|_DFF_P0|A4 _PG1_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P0|4|P _PG1_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P0|4|B _PG1_01|_DFF_P0|A4 _PG1_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P0|4|RB _PG1_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P0|T|1 _PG1_01|_DFF_P0|T1 _PG1_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P0|T|P _PG1_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P0|T|B _PG1_01|_DFF_P0|T1 _PG1_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P0|T|RB _PG1_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P0|45|1 _PG1_01|_DFF_P0|T2 _PG1_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_P0|45|B _PG1_01|_DFF_P0|T2 _PG1_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_P0|45|RB _PG1_01|_DFF_P0|45|MID_SHUNT _PG1_01|_DFF_P0|A4  2.1704737578552e-12
B_PG1_01|_DFF_P0|6|1 _PG1_01|_DFF_P0|Q1 _PG1_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P0|6|P _PG1_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P0|6|B _PG1_01|_DFF_P0|Q1 _PG1_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P0|6|RB _PG1_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_P1|I_1|B _PG1_01|_DFF_P1|A1 _PG1_01|_DFF_P1|I_1|MID  2e-12
I_PG1_01|_DFF_P1|I_1|B 0 _PG1_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_P1|I_3|B _PG1_01|_DFF_P1|A3 _PG1_01|_DFF_P1|I_3|MID  2e-12
I_PG1_01|_DFF_P1|I_3|B 0 _PG1_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_P1|I_T|B _PG1_01|_DFF_P1|T1 _PG1_01|_DFF_P1|I_T|MID  2e-12
I_PG1_01|_DFF_P1|I_T|B 0 _PG1_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_P1|I_6|B _PG1_01|_DFF_P1|Q1 _PG1_01|_DFF_P1|I_6|MID  2e-12
I_PG1_01|_DFF_P1|I_6|B 0 _PG1_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_P1|1|1 _PG1_01|_DFF_P1|A1 _PG1_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P1|1|P _PG1_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P1|1|B _PG1_01|_DFF_P1|A1 _PG1_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P1|1|RB _PG1_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P1|23|1 _PG1_01|_DFF_P1|A2 _PG1_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_P1|23|B _PG1_01|_DFF_P1|A2 _PG1_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_P1|23|RB _PG1_01|_DFF_P1|23|MID_SHUNT _PG1_01|_DFF_P1|A3  2.1704737578552e-12
B_PG1_01|_DFF_P1|3|1 _PG1_01|_DFF_P1|A3 _PG1_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P1|3|P _PG1_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P1|3|B _PG1_01|_DFF_P1|A3 _PG1_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P1|3|RB _PG1_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P1|4|1 _PG1_01|_DFF_P1|A4 _PG1_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P1|4|P _PG1_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P1|4|B _PG1_01|_DFF_P1|A4 _PG1_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P1|4|RB _PG1_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P1|T|1 _PG1_01|_DFF_P1|T1 _PG1_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P1|T|P _PG1_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P1|T|B _PG1_01|_DFF_P1|T1 _PG1_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P1|T|RB _PG1_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_P1|45|1 _PG1_01|_DFF_P1|T2 _PG1_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_P1|45|B _PG1_01|_DFF_P1|T2 _PG1_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_P1|45|RB _PG1_01|_DFF_P1|45|MID_SHUNT _PG1_01|_DFF_P1|A4  2.1704737578552e-12
B_PG1_01|_DFF_P1|6|1 _PG1_01|_DFF_P1|Q1 _PG1_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_P1|6|P _PG1_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_P1|6|B _PG1_01|_DFF_P1|Q1 _PG1_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_P1|6|RB _PG1_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_PG|I_1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|I_1|MID  2e-12
I_PG1_01|_DFF_PG|I_1|B 0 _PG1_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|I_3|MID  2e-12
I_PG1_01|_DFF_PG|I_3|B 0 _PG1_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_PG|I_T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|I_T|MID  2e-12
I_PG1_01|_DFF_PG|I_T|B 0 _PG1_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|I_6|MID  2e-12
I_PG1_01|_DFF_PG|I_6|B 0 _PG1_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_PG|1|1 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|1|P _PG1_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|1|RB _PG1_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|23|1 _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|23|B _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|23|RB _PG1_01|_DFF_PG|23|MID_SHUNT _PG1_01|_DFF_PG|A3  2.1704737578552e-12
B_PG1_01|_DFF_PG|3|1 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|3|P _PG1_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|3|RB _PG1_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|4|1 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|4|P _PG1_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|4|B _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|4|RB _PG1_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|T|1 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|T|P _PG1_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|T|RB _PG1_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|45|1 _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|45|B _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|45|RB _PG1_01|_DFF_PG|45|MID_SHUNT _PG1_01|_DFF_PG|A4  2.1704737578552e-12
B_PG1_01|_DFF_PG|6|1 _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|6|P _PG1_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|6|RB _PG1_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_GG|I_1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|I_1|MID  2e-12
I_PG1_01|_DFF_GG|I_1|B 0 _PG1_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|I_3|MID  2e-12
I_PG1_01|_DFF_GG|I_3|B 0 _PG1_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_GG|I_T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|I_T|MID  2e-12
I_PG1_01|_DFF_GG|I_T|B 0 _PG1_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|I_6|MID  2e-12
I_PG1_01|_DFF_GG|I_6|B 0 _PG1_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_GG|1|1 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|1|P _PG1_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|1|RB _PG1_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|23|1 _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|23|B _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|23|RB _PG1_01|_DFF_GG|23|MID_SHUNT _PG1_01|_DFF_GG|A3  2.1704737578552e-12
B_PG1_01|_DFF_GG|3|1 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|3|P _PG1_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|3|RB _PG1_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|4|1 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|4|P _PG1_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|4|B _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|4|RB _PG1_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|T|1 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|T|P _PG1_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|T|RB _PG1_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|45|1 _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|45|B _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|45|RB _PG1_01|_DFF_GG|45|MID_SHUNT _PG1_01|_DFF_GG|A4  2.1704737578552e-12
B_PG1_01|_DFF_GG|6|1 _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|6|P _PG1_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|6|RB _PG1_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_G|I_A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|I_A1|MID  2e-12
I_PG1_01|_AND_G|I_A1|B 0 _PG1_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|I_B1|MID  2e-12
I_PG1_01|_AND_G|I_B1|B 0 _PG1_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q3|B _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|I_Q3|MID  2e-12
I_PG1_01|_AND_G|I_Q3|B 0 _PG1_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_G|I_Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|I_Q2|MID  2e-12
I_PG1_01|_AND_G|I_Q2|B 0 _PG1_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|I_Q1|MID  2e-12
I_PG1_01|_AND_G|I_Q1|B 0 _PG1_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_G|A1|1 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A1|P _PG1_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A1|RB _PG1_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A2|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A2|P _PG1_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A2|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A2|RB _PG1_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A12|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|A12|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|A12|RB _PG1_01|_AND_G|A12|MID_SHUNT _PG1_01|_AND_G|A3  2.1704737578552e-12
B_PG1_01|_AND_G|B1|1 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B1|P _PG1_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B1|RB _PG1_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B2|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B2|P _PG1_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B2|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B2|RB _PG1_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B12|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|B12|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|B12|RB _PG1_01|_AND_G|B12|MID_SHUNT _PG1_01|_AND_G|B3  2.1704737578552e-12
B_PG1_01|_AND_G|Q2|1 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q2|P _PG1_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q2|RB _PG1_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|Q1|1 _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q1|P _PG1_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q1|RB _PG1_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_P|I_A1|B _PG1_01|_AND_P|A1 _PG1_01|_AND_P|I_A1|MID  2e-12
I_PG1_01|_AND_P|I_A1|B 0 _PG1_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_P|I_B1|B _PG1_01|_AND_P|B1 _PG1_01|_AND_P|I_B1|MID  2e-12
I_PG1_01|_AND_P|I_B1|B 0 _PG1_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_P|I_Q3|B _PG1_01|_AND_P|Q3 _PG1_01|_AND_P|I_Q3|MID  2e-12
I_PG1_01|_AND_P|I_Q3|B 0 _PG1_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_P|I_Q2|B _PG1_01|_AND_P|Q2 _PG1_01|_AND_P|I_Q2|MID  2e-12
I_PG1_01|_AND_P|I_Q2|B 0 _PG1_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_P|I_Q1|B _PG1_01|_AND_P|Q1 _PG1_01|_AND_P|I_Q1|MID  2e-12
I_PG1_01|_AND_P|I_Q1|B 0 _PG1_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_P|A1|1 _PG1_01|_AND_P|A1 _PG1_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_P|A1|P _PG1_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_P|A1|B _PG1_01|_AND_P|A1 _PG1_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_P|A1|RB _PG1_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_P|A2|1 _PG1_01|_AND_P|A2 _PG1_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_P|A2|P _PG1_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_P|A2|B _PG1_01|_AND_P|A2 _PG1_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_P|A2|RB _PG1_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_P|A12|1 _PG1_01|_AND_P|A2 _PG1_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_P|A12|B _PG1_01|_AND_P|A2 _PG1_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_P|A12|RB _PG1_01|_AND_P|A12|MID_SHUNT _PG1_01|_AND_P|A3  2.1704737578552e-12
B_PG1_01|_AND_P|B1|1 _PG1_01|_AND_P|B1 _PG1_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_P|B1|P _PG1_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_P|B1|B _PG1_01|_AND_P|B1 _PG1_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_P|B1|RB _PG1_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_P|B2|1 _PG1_01|_AND_P|B2 _PG1_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_P|B2|P _PG1_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_P|B2|B _PG1_01|_AND_P|B2 _PG1_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_P|B2|RB _PG1_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_P|B12|1 _PG1_01|_AND_P|B2 _PG1_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_P|B12|B _PG1_01|_AND_P|B2 _PG1_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_P|B12|RB _PG1_01|_AND_P|B12|MID_SHUNT _PG1_01|_AND_P|B3  2.1704737578552e-12
B_PG1_01|_AND_P|Q2|1 _PG1_01|_AND_P|Q2 _PG1_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_P|Q2|P _PG1_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_P|Q2|B _PG1_01|_AND_P|Q2 _PG1_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_P|Q2|RB _PG1_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_P|Q1|1 _PG1_01|_AND_P|Q1 _PG1_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_P|Q1|P _PG1_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_P|Q1|B _PG1_01|_AND_P|Q1 _PG1_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_P|Q1|RB _PG1_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|P|I_1|B _PG2_01|P|A1 _PG2_01|P|I_1|MID  2e-12
I_PG2_01|P|I_1|B 0 _PG2_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_3|B _PG2_01|P|A3 _PG2_01|P|I_3|MID  2e-12
I_PG2_01|P|I_3|B 0 _PG2_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|P|I_T|B _PG2_01|P|T1 _PG2_01|P|I_T|MID  2e-12
I_PG2_01|P|I_T|B 0 _PG2_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_6|B _PG2_01|P|Q1 _PG2_01|P|I_6|MID  2e-12
I_PG2_01|P|I_6|B 0 _PG2_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|P|1|1 _PG2_01|P|A1 _PG2_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|1|P _PG2_01|P|1|MID_SERIES 0  2e-13
R_PG2_01|P|1|B _PG2_01|P|A1 _PG2_01|P|1|MID_SHUNT  2.7439617672
L_PG2_01|P|1|RB _PG2_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|23|1 _PG2_01|P|A2 _PG2_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|P|23|B _PG2_01|P|A2 _PG2_01|P|23|MID_SHUNT  3.84154647408
L_PG2_01|P|23|RB _PG2_01|P|23|MID_SHUNT _PG2_01|P|A3  2.1704737578552e-12
B_PG2_01|P|3|1 _PG2_01|P|A3 _PG2_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|3|P _PG2_01|P|3|MID_SERIES 0  2e-13
R_PG2_01|P|3|B _PG2_01|P|A3 _PG2_01|P|3|MID_SHUNT  2.7439617672
L_PG2_01|P|3|RB _PG2_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|4|1 _PG2_01|P|A4 _PG2_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|4|P _PG2_01|P|4|MID_SERIES 0  2e-13
R_PG2_01|P|4|B _PG2_01|P|A4 _PG2_01|P|4|MID_SHUNT  2.7439617672
L_PG2_01|P|4|RB _PG2_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|T|1 _PG2_01|P|T1 _PG2_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|T|P _PG2_01|P|T|MID_SERIES 0  2e-13
R_PG2_01|P|T|B _PG2_01|P|T1 _PG2_01|P|T|MID_SHUNT  2.7439617672
L_PG2_01|P|T|RB _PG2_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|45|1 _PG2_01|P|T2 _PG2_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|P|45|B _PG2_01|P|T2 _PG2_01|P|45|MID_SHUNT  3.84154647408
L_PG2_01|P|45|RB _PG2_01|P|45|MID_SHUNT _PG2_01|P|A4  2.1704737578552e-12
B_PG2_01|P|6|1 _PG2_01|P|Q1 _PG2_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|6|P _PG2_01|P|6|MID_SERIES 0  2e-13
R_PG2_01|P|6|B _PG2_01|P|Q1 _PG2_01|P|6|MID_SHUNT  2.7439617672
L_PG2_01|P|6|RB _PG2_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|G|I_1|B _PG2_01|G|A1 _PG2_01|G|I_1|MID  2e-12
I_PG2_01|G|I_1|B 0 _PG2_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_3|B _PG2_01|G|A3 _PG2_01|G|I_3|MID  2e-12
I_PG2_01|G|I_3|B 0 _PG2_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|G|I_T|B _PG2_01|G|T1 _PG2_01|G|I_T|MID  2e-12
I_PG2_01|G|I_T|B 0 _PG2_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_6|B _PG2_01|G|Q1 _PG2_01|G|I_6|MID  2e-12
I_PG2_01|G|I_6|B 0 _PG2_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|G|1|1 _PG2_01|G|A1 _PG2_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|1|P _PG2_01|G|1|MID_SERIES 0  2e-13
R_PG2_01|G|1|B _PG2_01|G|A1 _PG2_01|G|1|MID_SHUNT  2.7439617672
L_PG2_01|G|1|RB _PG2_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|23|1 _PG2_01|G|A2 _PG2_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|G|23|B _PG2_01|G|A2 _PG2_01|G|23|MID_SHUNT  3.84154647408
L_PG2_01|G|23|RB _PG2_01|G|23|MID_SHUNT _PG2_01|G|A3  2.1704737578552e-12
B_PG2_01|G|3|1 _PG2_01|G|A3 _PG2_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|3|P _PG2_01|G|3|MID_SERIES 0  2e-13
R_PG2_01|G|3|B _PG2_01|G|A3 _PG2_01|G|3|MID_SHUNT  2.7439617672
L_PG2_01|G|3|RB _PG2_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|4|1 _PG2_01|G|A4 _PG2_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|4|P _PG2_01|G|4|MID_SERIES 0  2e-13
R_PG2_01|G|4|B _PG2_01|G|A4 _PG2_01|G|4|MID_SHUNT  2.7439617672
L_PG2_01|G|4|RB _PG2_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|T|1 _PG2_01|G|T1 _PG2_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|T|P _PG2_01|G|T|MID_SERIES 0  2e-13
R_PG2_01|G|T|B _PG2_01|G|T1 _PG2_01|G|T|MID_SHUNT  2.7439617672
L_PG2_01|G|T|RB _PG2_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|45|1 _PG2_01|G|T2 _PG2_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|G|45|B _PG2_01|G|T2 _PG2_01|G|45|MID_SHUNT  3.84154647408
L_PG2_01|G|45|RB _PG2_01|G|45|MID_SHUNT _PG2_01|G|A4  2.1704737578552e-12
B_PG2_01|G|6|1 _PG2_01|G|Q1 _PG2_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|6|P _PG2_01|G|6|MID_SERIES 0  2e-13
R_PG2_01|G|6|B _PG2_01|G|Q1 _PG2_01|G|6|MID_SHUNT  2.7439617672
L_PG2_01|G|6|RB _PG2_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_G1|I_D1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|I_D1|MID  2e-12
I_PG3_01|_SPL_G1|I_D1|B 0 _PG3_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_D2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|I_D2|MID  2e-12
I_PG3_01|_SPL_G1|I_D2|B 0 _PG3_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_G1|I_Q1|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|I_Q1|MID  2e-12
I_PG3_01|_SPL_G1|I_Q1|B 0 _PG3_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_Q2|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|I_Q2|MID  2e-12
I_PG3_01|_SPL_G1|I_Q2|B 0 _PG3_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_G1|1|1 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|1|P _PG3_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|1|RB _PG3_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|2|1 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|2|P _PG3_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|2|RB _PG3_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|A|1 _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|A|P _PG3_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|A|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|A|RB _PG3_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|B|1 _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|B|P _PG3_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|B|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|B|RB _PG3_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_P1|I_D1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|I_D1|MID  2e-12
I_PG3_01|_SPL_P1|I_D1|B 0 _PG3_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_D2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|I_D2|MID  2e-12
I_PG3_01|_SPL_P1|I_D2|B 0 _PG3_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_P1|I_Q1|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|I_Q1|MID  2e-12
I_PG3_01|_SPL_P1|I_Q1|B 0 _PG3_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_Q2|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|I_Q2|MID  2e-12
I_PG3_01|_SPL_P1|I_Q2|B 0 _PG3_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_P1|1|1 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|1|P _PG3_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|1|RB _PG3_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|2|1 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|2|P _PG3_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|2|RB _PG3_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|A|1 _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|A|P _PG3_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|A|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|A|RB _PG3_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|B|1 _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|B|P _PG3_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|B|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|B|RB _PG3_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_PG|I_A1|B _PG3_01|_PG|A1 _PG3_01|_PG|I_A1|MID  2e-12
I_PG3_01|_PG|I_A1|B 0 _PG3_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_B1|B _PG3_01|_PG|B1 _PG3_01|_PG|I_B1|MID  2e-12
I_PG3_01|_PG|I_B1|B 0 _PG3_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q3|B _PG3_01|_PG|Q3 _PG3_01|_PG|I_Q3|MID  2e-12
I_PG3_01|_PG|I_Q3|B 0 _PG3_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_PG|I_Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|I_Q2|MID  2e-12
I_PG3_01|_PG|I_Q2|B 0 _PG3_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|I_Q1|MID  2e-12
I_PG3_01|_PG|I_Q1|B 0 _PG3_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_PG|A1|1 _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A1|P _PG3_01|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01|_PG|A1|B _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A1|RB _PG3_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A2|1 _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A2|P _PG3_01|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01|_PG|A2|B _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A2|RB _PG3_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A12|1 _PG3_01|_PG|A2 _PG3_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|A12|B _PG3_01|_PG|A2 _PG3_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|A12|RB _PG3_01|_PG|A12|MID_SHUNT _PG3_01|_PG|A3  2.1704737578552e-12
B_PG3_01|_PG|B1|1 _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B1|P _PG3_01|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01|_PG|B1|B _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B1|RB _PG3_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B2|1 _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B2|P _PG3_01|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01|_PG|B2|B _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B2|RB _PG3_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B12|1 _PG3_01|_PG|B2 _PG3_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|B12|B _PG3_01|_PG|B2 _PG3_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|B12|RB _PG3_01|_PG|B12|MID_SHUNT _PG3_01|_PG|B3  2.1704737578552e-12
B_PG3_01|_PG|Q2|1 _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q2|P _PG3_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q2|RB _PG3_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|Q1|1 _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q1|P _PG3_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q1|RB _PG3_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_GG|I_A1|B _PG3_01|_GG|A1 _PG3_01|_GG|I_A1|MID  2e-12
I_PG3_01|_GG|I_A1|B 0 _PG3_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_B1|B _PG3_01|_GG|B1 _PG3_01|_GG|I_B1|MID  2e-12
I_PG3_01|_GG|I_B1|B 0 _PG3_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q3|B _PG3_01|_GG|Q3 _PG3_01|_GG|I_Q3|MID  2e-12
I_PG3_01|_GG|I_Q3|B 0 _PG3_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_GG|I_Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|I_Q2|MID  2e-12
I_PG3_01|_GG|I_Q2|B 0 _PG3_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|I_Q1|MID  2e-12
I_PG3_01|_GG|I_Q1|B 0 _PG3_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_GG|A1|1 _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A1|P _PG3_01|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01|_GG|A1|B _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A1|RB _PG3_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A2|1 _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A2|P _PG3_01|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01|_GG|A2|B _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A2|RB _PG3_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A12|1 _PG3_01|_GG|A2 _PG3_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|A12|B _PG3_01|_GG|A2 _PG3_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|A12|RB _PG3_01|_GG|A12|MID_SHUNT _PG3_01|_GG|A3  2.1704737578552e-12
B_PG3_01|_GG|B1|1 _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B1|P _PG3_01|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01|_GG|B1|B _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B1|RB _PG3_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B2|1 _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B2|P _PG3_01|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01|_GG|B2|B _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B2|RB _PG3_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B12|1 _PG3_01|_GG|B2 _PG3_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|B12|B _PG3_01|_GG|B2 _PG3_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|B12|RB _PG3_01|_GG|B12|MID_SHUNT _PG3_01|_GG|B3  2.1704737578552e-12
B_PG3_01|_GG|Q2|1 _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q2|P _PG3_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q2|RB _PG3_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|Q1|1 _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q1|P _PG3_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q1|RB _PG3_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P0|I_1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|I_1|MID  2e-12
I_PG3_01|_DFF_P0|I_1|B 0 _PG3_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|I_3|MID  2e-12
I_PG3_01|_DFF_P0|I_3|B 0 _PG3_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P0|I_T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|I_T|MID  2e-12
I_PG3_01|_DFF_P0|I_T|B 0 _PG3_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|I_6|MID  2e-12
I_PG3_01|_DFF_P0|I_6|B 0 _PG3_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P0|1|1 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|1|P _PG3_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|1|RB _PG3_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|23|1 _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|23|B _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|23|RB _PG3_01|_DFF_P0|23|MID_SHUNT _PG3_01|_DFF_P0|A3  2.1704737578552e-12
B_PG3_01|_DFF_P0|3|1 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|3|P _PG3_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|3|RB _PG3_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|4|1 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|4|P _PG3_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|4|B _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|4|RB _PG3_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|T|1 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|T|P _PG3_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|T|RB _PG3_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|45|1 _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|45|B _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|45|RB _PG3_01|_DFF_P0|45|MID_SHUNT _PG3_01|_DFF_P0|A4  2.1704737578552e-12
B_PG3_01|_DFF_P0|6|1 _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|6|P _PG3_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|6|RB _PG3_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P1|I_1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|I_1|MID  2e-12
I_PG3_01|_DFF_P1|I_1|B 0 _PG3_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|I_3|MID  2e-12
I_PG3_01|_DFF_P1|I_3|B 0 _PG3_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P1|I_T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|I_T|MID  2e-12
I_PG3_01|_DFF_P1|I_T|B 0 _PG3_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|I_6|MID  2e-12
I_PG3_01|_DFF_P1|I_6|B 0 _PG3_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P1|1|1 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|1|P _PG3_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|1|RB _PG3_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|23|1 _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|23|B _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|23|RB _PG3_01|_DFF_P1|23|MID_SHUNT _PG3_01|_DFF_P1|A3  2.1704737578552e-12
B_PG3_01|_DFF_P1|3|1 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|3|P _PG3_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|3|RB _PG3_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|4|1 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|4|P _PG3_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|4|B _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|4|RB _PG3_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|T|1 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|T|P _PG3_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|T|RB _PG3_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|45|1 _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|45|B _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|45|RB _PG3_01|_DFF_P1|45|MID_SHUNT _PG3_01|_DFF_P1|A4  2.1704737578552e-12
B_PG3_01|_DFF_P1|6|1 _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|6|P _PG3_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|6|RB _PG3_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_PG|I_1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|I_1|MID  2e-12
I_PG3_01|_DFF_PG|I_1|B 0 _PG3_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|I_3|MID  2e-12
I_PG3_01|_DFF_PG|I_3|B 0 _PG3_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_PG|I_T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|I_T|MID  2e-12
I_PG3_01|_DFF_PG|I_T|B 0 _PG3_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|I_6|MID  2e-12
I_PG3_01|_DFF_PG|I_6|B 0 _PG3_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_PG|1|1 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|1|P _PG3_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|1|RB _PG3_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|23|1 _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|23|B _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|23|RB _PG3_01|_DFF_PG|23|MID_SHUNT _PG3_01|_DFF_PG|A3  2.1704737578552e-12
B_PG3_01|_DFF_PG|3|1 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|3|P _PG3_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|3|RB _PG3_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|4|1 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|4|P _PG3_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|4|B _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|4|RB _PG3_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|T|1 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|T|P _PG3_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|T|RB _PG3_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|45|1 _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|45|B _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|45|RB _PG3_01|_DFF_PG|45|MID_SHUNT _PG3_01|_DFF_PG|A4  2.1704737578552e-12
B_PG3_01|_DFF_PG|6|1 _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|6|P _PG3_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|6|RB _PG3_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_GG|I_1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|I_1|MID  2e-12
I_PG3_01|_DFF_GG|I_1|B 0 _PG3_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|I_3|MID  2e-12
I_PG3_01|_DFF_GG|I_3|B 0 _PG3_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_GG|I_T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|I_T|MID  2e-12
I_PG3_01|_DFF_GG|I_T|B 0 _PG3_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|I_6|MID  2e-12
I_PG3_01|_DFF_GG|I_6|B 0 _PG3_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_GG|1|1 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|1|P _PG3_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|1|RB _PG3_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|23|1 _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|23|B _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|23|RB _PG3_01|_DFF_GG|23|MID_SHUNT _PG3_01|_DFF_GG|A3  2.1704737578552e-12
B_PG3_01|_DFF_GG|3|1 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|3|P _PG3_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|3|RB _PG3_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|4|1 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|4|P _PG3_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|4|B _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|4|RB _PG3_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|T|1 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|T|P _PG3_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|T|RB _PG3_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|45|1 _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|45|B _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|45|RB _PG3_01|_DFF_GG|45|MID_SHUNT _PG3_01|_DFF_GG|A4  2.1704737578552e-12
B_PG3_01|_DFF_GG|6|1 _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|6|P _PG3_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|6|RB _PG3_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_G|I_A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|I_A1|MID  2e-12
I_PG3_01|_AND_G|I_A1|B 0 _PG3_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|I_B1|MID  2e-12
I_PG3_01|_AND_G|I_B1|B 0 _PG3_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q3|B _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|I_Q3|MID  2e-12
I_PG3_01|_AND_G|I_Q3|B 0 _PG3_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_G|I_Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|I_Q2|MID  2e-12
I_PG3_01|_AND_G|I_Q2|B 0 _PG3_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|I_Q1|MID  2e-12
I_PG3_01|_AND_G|I_Q1|B 0 _PG3_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_G|A1|1 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A1|P _PG3_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A1|RB _PG3_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A2|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A2|P _PG3_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A2|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A2|RB _PG3_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A12|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|A12|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|A12|RB _PG3_01|_AND_G|A12|MID_SHUNT _PG3_01|_AND_G|A3  2.1704737578552e-12
B_PG3_01|_AND_G|B1|1 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B1|P _PG3_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B1|RB _PG3_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B2|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B2|P _PG3_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B2|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B2|RB _PG3_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B12|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|B12|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|B12|RB _PG3_01|_AND_G|B12|MID_SHUNT _PG3_01|_AND_G|B3  2.1704737578552e-12
B_PG3_01|_AND_G|Q2|1 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q2|P _PG3_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q2|RB _PG3_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|Q1|1 _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q1|P _PG3_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q1|RB _PG3_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_P|I_A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|I_A1|MID  2e-12
I_PG3_01|_AND_P|I_A1|B 0 _PG3_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|I_B1|MID  2e-12
I_PG3_01|_AND_P|I_B1|B 0 _PG3_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q3|B _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|I_Q3|MID  2e-12
I_PG3_01|_AND_P|I_Q3|B 0 _PG3_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_P|I_Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|I_Q2|MID  2e-12
I_PG3_01|_AND_P|I_Q2|B 0 _PG3_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|I_Q1|MID  2e-12
I_PG3_01|_AND_P|I_Q1|B 0 _PG3_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_P|A1|1 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A1|P _PG3_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A1|RB _PG3_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A2|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A2|P _PG3_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A2|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A2|RB _PG3_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A12|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|A12|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|A12|RB _PG3_01|_AND_P|A12|MID_SHUNT _PG3_01|_AND_P|A3  2.1704737578552e-12
B_PG3_01|_AND_P|B1|1 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B1|P _PG3_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B1|RB _PG3_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B2|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B2|P _PG3_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B2|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B2|RB _PG3_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B12|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|B12|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|B12|RB _PG3_01|_AND_P|B12|MID_SHUNT _PG3_01|_AND_P|B3  2.1704737578552e-12
B_PG3_01|_AND_P|Q2|1 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q2|P _PG3_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q2|RB _PG3_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|Q1|1 _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q1|P _PG3_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q1|RB _PG3_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG4_01|P|I_1|B _PG4_01|P|A1 _PG4_01|P|I_1|MID  2e-12
I_PG4_01|P|I_1|B 0 _PG4_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_01|P|I_3|B _PG4_01|P|A3 _PG4_01|P|I_3|MID  2e-12
I_PG4_01|P|I_3|B 0 _PG4_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_01|P|I_T|B _PG4_01|P|T1 _PG4_01|P|I_T|MID  2e-12
I_PG4_01|P|I_T|B 0 _PG4_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_01|P|I_6|B _PG4_01|P|Q1 _PG4_01|P|I_6|MID  2e-12
I_PG4_01|P|I_6|B 0 _PG4_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_01|P|1|1 _PG4_01|P|A1 _PG4_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG4_01|P|1|P _PG4_01|P|1|MID_SERIES 0  2e-13
R_PG4_01|P|1|B _PG4_01|P|A1 _PG4_01|P|1|MID_SHUNT  2.7439617672
L_PG4_01|P|1|RB _PG4_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|P|23|1 _PG4_01|P|A2 _PG4_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG4_01|P|23|B _PG4_01|P|A2 _PG4_01|P|23|MID_SHUNT  3.84154647408
L_PG4_01|P|23|RB _PG4_01|P|23|MID_SHUNT _PG4_01|P|A3  2.1704737578552e-12
B_PG4_01|P|3|1 _PG4_01|P|A3 _PG4_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG4_01|P|3|P _PG4_01|P|3|MID_SERIES 0  2e-13
R_PG4_01|P|3|B _PG4_01|P|A3 _PG4_01|P|3|MID_SHUNT  2.7439617672
L_PG4_01|P|3|RB _PG4_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|P|4|1 _PG4_01|P|A4 _PG4_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG4_01|P|4|P _PG4_01|P|4|MID_SERIES 0  2e-13
R_PG4_01|P|4|B _PG4_01|P|A4 _PG4_01|P|4|MID_SHUNT  2.7439617672
L_PG4_01|P|4|RB _PG4_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|P|T|1 _PG4_01|P|T1 _PG4_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG4_01|P|T|P _PG4_01|P|T|MID_SERIES 0  2e-13
R_PG4_01|P|T|B _PG4_01|P|T1 _PG4_01|P|T|MID_SHUNT  2.7439617672
L_PG4_01|P|T|RB _PG4_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|P|45|1 _PG4_01|P|T2 _PG4_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG4_01|P|45|B _PG4_01|P|T2 _PG4_01|P|45|MID_SHUNT  3.84154647408
L_PG4_01|P|45|RB _PG4_01|P|45|MID_SHUNT _PG4_01|P|A4  2.1704737578552e-12
B_PG4_01|P|6|1 _PG4_01|P|Q1 _PG4_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG4_01|P|6|P _PG4_01|P|6|MID_SERIES 0  2e-13
R_PG4_01|P|6|B _PG4_01|P|Q1 _PG4_01|P|6|MID_SHUNT  2.7439617672
L_PG4_01|P|6|RB _PG4_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_01|G|I_1|B _PG4_01|G|A1 _PG4_01|G|I_1|MID  2e-12
I_PG4_01|G|I_1|B 0 _PG4_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_01|G|I_3|B _PG4_01|G|A3 _PG4_01|G|I_3|MID  2e-12
I_PG4_01|G|I_3|B 0 _PG4_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_01|G|I_T|B _PG4_01|G|T1 _PG4_01|G|I_T|MID  2e-12
I_PG4_01|G|I_T|B 0 _PG4_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_01|G|I_6|B _PG4_01|G|Q1 _PG4_01|G|I_6|MID  2e-12
I_PG4_01|G|I_6|B 0 _PG4_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_01|G|1|1 _PG4_01|G|A1 _PG4_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG4_01|G|1|P _PG4_01|G|1|MID_SERIES 0  2e-13
R_PG4_01|G|1|B _PG4_01|G|A1 _PG4_01|G|1|MID_SHUNT  2.7439617672
L_PG4_01|G|1|RB _PG4_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|G|23|1 _PG4_01|G|A2 _PG4_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG4_01|G|23|B _PG4_01|G|A2 _PG4_01|G|23|MID_SHUNT  3.84154647408
L_PG4_01|G|23|RB _PG4_01|G|23|MID_SHUNT _PG4_01|G|A3  2.1704737578552e-12
B_PG4_01|G|3|1 _PG4_01|G|A3 _PG4_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG4_01|G|3|P _PG4_01|G|3|MID_SERIES 0  2e-13
R_PG4_01|G|3|B _PG4_01|G|A3 _PG4_01|G|3|MID_SHUNT  2.7439617672
L_PG4_01|G|3|RB _PG4_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|G|4|1 _PG4_01|G|A4 _PG4_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG4_01|G|4|P _PG4_01|G|4|MID_SERIES 0  2e-13
R_PG4_01|G|4|B _PG4_01|G|A4 _PG4_01|G|4|MID_SHUNT  2.7439617672
L_PG4_01|G|4|RB _PG4_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|G|T|1 _PG4_01|G|T1 _PG4_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG4_01|G|T|P _PG4_01|G|T|MID_SERIES 0  2e-13
R_PG4_01|G|T|B _PG4_01|G|T1 _PG4_01|G|T|MID_SHUNT  2.7439617672
L_PG4_01|G|T|RB _PG4_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_01|G|45|1 _PG4_01|G|T2 _PG4_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG4_01|G|45|B _PG4_01|G|T2 _PG4_01|G|45|MID_SHUNT  3.84154647408
L_PG4_01|G|45|RB _PG4_01|G|45|MID_SHUNT _PG4_01|G|A4  2.1704737578552e-12
B_PG4_01|G|6|1 _PG4_01|G|Q1 _PG4_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG4_01|G|6|P _PG4_01|G|6|MID_SERIES 0  2e-13
R_PG4_01|G|6|B _PG4_01|G|Q1 _PG4_01|G|6|MID_SHUNT  2.7439617672
L_PG4_01|G|6|RB _PG4_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_SPL_G1|I_D1|B _PG5_01|_SPL_G1|D1 _PG5_01|_SPL_G1|I_D1|MID  2e-12
I_PG5_01|_SPL_G1|I_D1|B 0 _PG5_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_01|_SPL_G1|I_D2|B _PG5_01|_SPL_G1|D2 _PG5_01|_SPL_G1|I_D2|MID  2e-12
I_PG5_01|_SPL_G1|I_D2|B 0 _PG5_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG5_01|_SPL_G1|I_Q1|B _PG5_01|_SPL_G1|QA1 _PG5_01|_SPL_G1|I_Q1|MID  2e-12
I_PG5_01|_SPL_G1|I_Q1|B 0 _PG5_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_01|_SPL_G1|I_Q2|B _PG5_01|_SPL_G1|QB1 _PG5_01|_SPL_G1|I_Q2|MID  2e-12
I_PG5_01|_SPL_G1|I_Q2|B 0 _PG5_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG5_01|_SPL_G1|1|1 _PG5_01|_SPL_G1|D1 _PG5_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_G1|1|P _PG5_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG5_01|_SPL_G1|1|B _PG5_01|_SPL_G1|D1 _PG5_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_G1|1|RB _PG5_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_SPL_G1|2|1 _PG5_01|_SPL_G1|D2 _PG5_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_G1|2|P _PG5_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG5_01|_SPL_G1|2|B _PG5_01|_SPL_G1|D2 _PG5_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_G1|2|RB _PG5_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_SPL_G1|A|1 _PG5_01|_SPL_G1|QA1 _PG5_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_G1|A|P _PG5_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG5_01|_SPL_G1|A|B _PG5_01|_SPL_G1|QA1 _PG5_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_G1|A|RB _PG5_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_SPL_G1|B|1 _PG5_01|_SPL_G1|QB1 _PG5_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_G1|B|P _PG5_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG5_01|_SPL_G1|B|B _PG5_01|_SPL_G1|QB1 _PG5_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_G1|B|RB _PG5_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_SPL_P1|I_D1|B _PG5_01|_SPL_P1|D1 _PG5_01|_SPL_P1|I_D1|MID  2e-12
I_PG5_01|_SPL_P1|I_D1|B 0 _PG5_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_01|_SPL_P1|I_D2|B _PG5_01|_SPL_P1|D2 _PG5_01|_SPL_P1|I_D2|MID  2e-12
I_PG5_01|_SPL_P1|I_D2|B 0 _PG5_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG5_01|_SPL_P1|I_Q1|B _PG5_01|_SPL_P1|QA1 _PG5_01|_SPL_P1|I_Q1|MID  2e-12
I_PG5_01|_SPL_P1|I_Q1|B 0 _PG5_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_01|_SPL_P1|I_Q2|B _PG5_01|_SPL_P1|QB1 _PG5_01|_SPL_P1|I_Q2|MID  2e-12
I_PG5_01|_SPL_P1|I_Q2|B 0 _PG5_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG5_01|_SPL_P1|1|1 _PG5_01|_SPL_P1|D1 _PG5_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_P1|1|P _PG5_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG5_01|_SPL_P1|1|B _PG5_01|_SPL_P1|D1 _PG5_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_P1|1|RB _PG5_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_SPL_P1|2|1 _PG5_01|_SPL_P1|D2 _PG5_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_P1|2|P _PG5_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG5_01|_SPL_P1|2|B _PG5_01|_SPL_P1|D2 _PG5_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_P1|2|RB _PG5_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_SPL_P1|A|1 _PG5_01|_SPL_P1|QA1 _PG5_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_P1|A|P _PG5_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG5_01|_SPL_P1|A|B _PG5_01|_SPL_P1|QA1 _PG5_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_P1|A|RB _PG5_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_SPL_P1|B|1 _PG5_01|_SPL_P1|QB1 _PG5_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_SPL_P1|B|P _PG5_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG5_01|_SPL_P1|B|B _PG5_01|_SPL_P1|QB1 _PG5_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG5_01|_SPL_P1|B|RB _PG5_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_PG|I_A1|B _PG5_01|_PG|A1 _PG5_01|_PG|I_A1|MID  2e-12
I_PG5_01|_PG|I_A1|B 0 _PG5_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_PG|I_B1|B _PG5_01|_PG|B1 _PG5_01|_PG|I_B1|MID  2e-12
I_PG5_01|_PG|I_B1|B 0 _PG5_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_PG|I_Q3|B _PG5_01|_PG|Q3 _PG5_01|_PG|I_Q3|MID  2e-12
I_PG5_01|_PG|I_Q3|B 0 _PG5_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_01|_PG|I_Q2|B _PG5_01|_PG|Q2 _PG5_01|_PG|I_Q2|MID  2e-12
I_PG5_01|_PG|I_Q2|B 0 _PG5_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_PG|I_Q1|B _PG5_01|_PG|Q1 _PG5_01|_PG|I_Q1|MID  2e-12
I_PG5_01|_PG|I_Q1|B 0 _PG5_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_PG|A1|1 _PG5_01|_PG|A1 _PG5_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_PG|A1|P _PG5_01|_PG|A1|MID_SERIES 0  2e-13
R_PG5_01|_PG|A1|B _PG5_01|_PG|A1 _PG5_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG5_01|_PG|A1|RB _PG5_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_PG|A2|1 _PG5_01|_PG|A2 _PG5_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_PG|A2|P _PG5_01|_PG|A2|MID_SERIES 0  2e-13
R_PG5_01|_PG|A2|B _PG5_01|_PG|A2 _PG5_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG5_01|_PG|A2|RB _PG5_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_PG|A12|1 _PG5_01|_PG|A2 _PG5_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_PG|A12|B _PG5_01|_PG|A2 _PG5_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG5_01|_PG|A12|RB _PG5_01|_PG|A12|MID_SHUNT _PG5_01|_PG|A3  2.1704737578552e-12
B_PG5_01|_PG|B1|1 _PG5_01|_PG|B1 _PG5_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_PG|B1|P _PG5_01|_PG|B1|MID_SERIES 0  2e-13
R_PG5_01|_PG|B1|B _PG5_01|_PG|B1 _PG5_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG5_01|_PG|B1|RB _PG5_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_PG|B2|1 _PG5_01|_PG|B2 _PG5_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_PG|B2|P _PG5_01|_PG|B2|MID_SERIES 0  2e-13
R_PG5_01|_PG|B2|B _PG5_01|_PG|B2 _PG5_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG5_01|_PG|B2|RB _PG5_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_PG|B12|1 _PG5_01|_PG|B2 _PG5_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG5_01|_PG|B12|B _PG5_01|_PG|B2 _PG5_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG5_01|_PG|B12|RB _PG5_01|_PG|B12|MID_SHUNT _PG5_01|_PG|B3  2.1704737578552e-12
B_PG5_01|_PG|Q2|1 _PG5_01|_PG|Q2 _PG5_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_PG|Q2|P _PG5_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG5_01|_PG|Q2|B _PG5_01|_PG|Q2 _PG5_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG5_01|_PG|Q2|RB _PG5_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_PG|Q1|1 _PG5_01|_PG|Q1 _PG5_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_PG|Q1|P _PG5_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG5_01|_PG|Q1|B _PG5_01|_PG|Q1 _PG5_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG5_01|_PG|Q1|RB _PG5_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_GG|I_A1|B _PG5_01|_GG|A1 _PG5_01|_GG|I_A1|MID  2e-12
I_PG5_01|_GG|I_A1|B 0 _PG5_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_GG|I_B1|B _PG5_01|_GG|B1 _PG5_01|_GG|I_B1|MID  2e-12
I_PG5_01|_GG|I_B1|B 0 _PG5_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_GG|I_Q3|B _PG5_01|_GG|Q3 _PG5_01|_GG|I_Q3|MID  2e-12
I_PG5_01|_GG|I_Q3|B 0 _PG5_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_01|_GG|I_Q2|B _PG5_01|_GG|Q2 _PG5_01|_GG|I_Q2|MID  2e-12
I_PG5_01|_GG|I_Q2|B 0 _PG5_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_GG|I_Q1|B _PG5_01|_GG|Q1 _PG5_01|_GG|I_Q1|MID  2e-12
I_PG5_01|_GG|I_Q1|B 0 _PG5_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_GG|A1|1 _PG5_01|_GG|A1 _PG5_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_GG|A1|P _PG5_01|_GG|A1|MID_SERIES 0  2e-13
R_PG5_01|_GG|A1|B _PG5_01|_GG|A1 _PG5_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG5_01|_GG|A1|RB _PG5_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_GG|A2|1 _PG5_01|_GG|A2 _PG5_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_GG|A2|P _PG5_01|_GG|A2|MID_SERIES 0  2e-13
R_PG5_01|_GG|A2|B _PG5_01|_GG|A2 _PG5_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG5_01|_GG|A2|RB _PG5_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_GG|A12|1 _PG5_01|_GG|A2 _PG5_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_GG|A12|B _PG5_01|_GG|A2 _PG5_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG5_01|_GG|A12|RB _PG5_01|_GG|A12|MID_SHUNT _PG5_01|_GG|A3  2.1704737578552e-12
B_PG5_01|_GG|B1|1 _PG5_01|_GG|B1 _PG5_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_GG|B1|P _PG5_01|_GG|B1|MID_SERIES 0  2e-13
R_PG5_01|_GG|B1|B _PG5_01|_GG|B1 _PG5_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG5_01|_GG|B1|RB _PG5_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_GG|B2|1 _PG5_01|_GG|B2 _PG5_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_GG|B2|P _PG5_01|_GG|B2|MID_SERIES 0  2e-13
R_PG5_01|_GG|B2|B _PG5_01|_GG|B2 _PG5_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG5_01|_GG|B2|RB _PG5_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_GG|B12|1 _PG5_01|_GG|B2 _PG5_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG5_01|_GG|B12|B _PG5_01|_GG|B2 _PG5_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG5_01|_GG|B12|RB _PG5_01|_GG|B12|MID_SHUNT _PG5_01|_GG|B3  2.1704737578552e-12
B_PG5_01|_GG|Q2|1 _PG5_01|_GG|Q2 _PG5_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_GG|Q2|P _PG5_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG5_01|_GG|Q2|B _PG5_01|_GG|Q2 _PG5_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG5_01|_GG|Q2|RB _PG5_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_GG|Q1|1 _PG5_01|_GG|Q1 _PG5_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_GG|Q1|P _PG5_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG5_01|_GG|Q1|B _PG5_01|_GG|Q1 _PG5_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG5_01|_GG|Q1|RB _PG5_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_DFF_P0|I_1|B _PG5_01|_DFF_P0|A1 _PG5_01|_DFF_P0|I_1|MID  2e-12
I_PG5_01|_DFF_P0|I_1|B 0 _PG5_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_P0|I_3|B _PG5_01|_DFF_P0|A3 _PG5_01|_DFF_P0|I_3|MID  2e-12
I_PG5_01|_DFF_P0|I_3|B 0 _PG5_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_01|_DFF_P0|I_T|B _PG5_01|_DFF_P0|T1 _PG5_01|_DFF_P0|I_T|MID  2e-12
I_PG5_01|_DFF_P0|I_T|B 0 _PG5_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_P0|I_6|B _PG5_01|_DFF_P0|Q1 _PG5_01|_DFF_P0|I_6|MID  2e-12
I_PG5_01|_DFF_P0|I_6|B 0 _PG5_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_DFF_P0|1|1 _PG5_01|_DFF_P0|A1 _PG5_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P0|1|P _PG5_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P0|1|B _PG5_01|_DFF_P0|A1 _PG5_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P0|1|RB _PG5_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P0|23|1 _PG5_01|_DFF_P0|A2 _PG5_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_P0|23|B _PG5_01|_DFF_P0|A2 _PG5_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_P0|23|RB _PG5_01|_DFF_P0|23|MID_SHUNT _PG5_01|_DFF_P0|A3  2.1704737578552e-12
B_PG5_01|_DFF_P0|3|1 _PG5_01|_DFF_P0|A3 _PG5_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P0|3|P _PG5_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P0|3|B _PG5_01|_DFF_P0|A3 _PG5_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P0|3|RB _PG5_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P0|4|1 _PG5_01|_DFF_P0|A4 _PG5_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P0|4|P _PG5_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P0|4|B _PG5_01|_DFF_P0|A4 _PG5_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P0|4|RB _PG5_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P0|T|1 _PG5_01|_DFF_P0|T1 _PG5_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P0|T|P _PG5_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P0|T|B _PG5_01|_DFF_P0|T1 _PG5_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P0|T|RB _PG5_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P0|45|1 _PG5_01|_DFF_P0|T2 _PG5_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_P0|45|B _PG5_01|_DFF_P0|T2 _PG5_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_P0|45|RB _PG5_01|_DFF_P0|45|MID_SHUNT _PG5_01|_DFF_P0|A4  2.1704737578552e-12
B_PG5_01|_DFF_P0|6|1 _PG5_01|_DFF_P0|Q1 _PG5_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P0|6|P _PG5_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P0|6|B _PG5_01|_DFF_P0|Q1 _PG5_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P0|6|RB _PG5_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_DFF_P1|I_1|B _PG5_01|_DFF_P1|A1 _PG5_01|_DFF_P1|I_1|MID  2e-12
I_PG5_01|_DFF_P1|I_1|B 0 _PG5_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_P1|I_3|B _PG5_01|_DFF_P1|A3 _PG5_01|_DFF_P1|I_3|MID  2e-12
I_PG5_01|_DFF_P1|I_3|B 0 _PG5_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_01|_DFF_P1|I_T|B _PG5_01|_DFF_P1|T1 _PG5_01|_DFF_P1|I_T|MID  2e-12
I_PG5_01|_DFF_P1|I_T|B 0 _PG5_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_P1|I_6|B _PG5_01|_DFF_P1|Q1 _PG5_01|_DFF_P1|I_6|MID  2e-12
I_PG5_01|_DFF_P1|I_6|B 0 _PG5_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_DFF_P1|1|1 _PG5_01|_DFF_P1|A1 _PG5_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P1|1|P _PG5_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P1|1|B _PG5_01|_DFF_P1|A1 _PG5_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P1|1|RB _PG5_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P1|23|1 _PG5_01|_DFF_P1|A2 _PG5_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_P1|23|B _PG5_01|_DFF_P1|A2 _PG5_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_P1|23|RB _PG5_01|_DFF_P1|23|MID_SHUNT _PG5_01|_DFF_P1|A3  2.1704737578552e-12
B_PG5_01|_DFF_P1|3|1 _PG5_01|_DFF_P1|A3 _PG5_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P1|3|P _PG5_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P1|3|B _PG5_01|_DFF_P1|A3 _PG5_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P1|3|RB _PG5_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P1|4|1 _PG5_01|_DFF_P1|A4 _PG5_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P1|4|P _PG5_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P1|4|B _PG5_01|_DFF_P1|A4 _PG5_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P1|4|RB _PG5_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P1|T|1 _PG5_01|_DFF_P1|T1 _PG5_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P1|T|P _PG5_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P1|T|B _PG5_01|_DFF_P1|T1 _PG5_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P1|T|RB _PG5_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_P1|45|1 _PG5_01|_DFF_P1|T2 _PG5_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_P1|45|B _PG5_01|_DFF_P1|T2 _PG5_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_P1|45|RB _PG5_01|_DFF_P1|45|MID_SHUNT _PG5_01|_DFF_P1|A4  2.1704737578552e-12
B_PG5_01|_DFF_P1|6|1 _PG5_01|_DFF_P1|Q1 _PG5_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_P1|6|P _PG5_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG5_01|_DFF_P1|6|B _PG5_01|_DFF_P1|Q1 _PG5_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_P1|6|RB _PG5_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_DFF_PG|I_1|B _PG5_01|_DFF_PG|A1 _PG5_01|_DFF_PG|I_1|MID  2e-12
I_PG5_01|_DFF_PG|I_1|B 0 _PG5_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_PG|I_3|B _PG5_01|_DFF_PG|A3 _PG5_01|_DFF_PG|I_3|MID  2e-12
I_PG5_01|_DFF_PG|I_3|B 0 _PG5_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_01|_DFF_PG|I_T|B _PG5_01|_DFF_PG|T1 _PG5_01|_DFF_PG|I_T|MID  2e-12
I_PG5_01|_DFF_PG|I_T|B 0 _PG5_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_PG|I_6|B _PG5_01|_DFF_PG|Q1 _PG5_01|_DFF_PG|I_6|MID  2e-12
I_PG5_01|_DFF_PG|I_6|B 0 _PG5_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_DFF_PG|1|1 _PG5_01|_DFF_PG|A1 _PG5_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_PG|1|P _PG5_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG5_01|_DFF_PG|1|B _PG5_01|_DFF_PG|A1 _PG5_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_PG|1|RB _PG5_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_PG|23|1 _PG5_01|_DFF_PG|A2 _PG5_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_PG|23|B _PG5_01|_DFF_PG|A2 _PG5_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_PG|23|RB _PG5_01|_DFF_PG|23|MID_SHUNT _PG5_01|_DFF_PG|A3  2.1704737578552e-12
B_PG5_01|_DFF_PG|3|1 _PG5_01|_DFF_PG|A3 _PG5_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_PG|3|P _PG5_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG5_01|_DFF_PG|3|B _PG5_01|_DFF_PG|A3 _PG5_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_PG|3|RB _PG5_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_PG|4|1 _PG5_01|_DFF_PG|A4 _PG5_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_PG|4|P _PG5_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG5_01|_DFF_PG|4|B _PG5_01|_DFF_PG|A4 _PG5_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_PG|4|RB _PG5_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_PG|T|1 _PG5_01|_DFF_PG|T1 _PG5_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_PG|T|P _PG5_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG5_01|_DFF_PG|T|B _PG5_01|_DFF_PG|T1 _PG5_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_PG|T|RB _PG5_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_PG|45|1 _PG5_01|_DFF_PG|T2 _PG5_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_PG|45|B _PG5_01|_DFF_PG|T2 _PG5_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_PG|45|RB _PG5_01|_DFF_PG|45|MID_SHUNT _PG5_01|_DFF_PG|A4  2.1704737578552e-12
B_PG5_01|_DFF_PG|6|1 _PG5_01|_DFF_PG|Q1 _PG5_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_PG|6|P _PG5_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG5_01|_DFF_PG|6|B _PG5_01|_DFF_PG|Q1 _PG5_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_PG|6|RB _PG5_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_DFF_GG|I_1|B _PG5_01|_DFF_GG|A1 _PG5_01|_DFF_GG|I_1|MID  2e-12
I_PG5_01|_DFF_GG|I_1|B 0 _PG5_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_GG|I_3|B _PG5_01|_DFF_GG|A3 _PG5_01|_DFF_GG|I_3|MID  2e-12
I_PG5_01|_DFF_GG|I_3|B 0 _PG5_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_01|_DFF_GG|I_T|B _PG5_01|_DFF_GG|T1 _PG5_01|_DFF_GG|I_T|MID  2e-12
I_PG5_01|_DFF_GG|I_T|B 0 _PG5_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_DFF_GG|I_6|B _PG5_01|_DFF_GG|Q1 _PG5_01|_DFF_GG|I_6|MID  2e-12
I_PG5_01|_DFF_GG|I_6|B 0 _PG5_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_DFF_GG|1|1 _PG5_01|_DFF_GG|A1 _PG5_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_GG|1|P _PG5_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG5_01|_DFF_GG|1|B _PG5_01|_DFF_GG|A1 _PG5_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_GG|1|RB _PG5_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_GG|23|1 _PG5_01|_DFF_GG|A2 _PG5_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_GG|23|B _PG5_01|_DFF_GG|A2 _PG5_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_GG|23|RB _PG5_01|_DFF_GG|23|MID_SHUNT _PG5_01|_DFF_GG|A3  2.1704737578552e-12
B_PG5_01|_DFF_GG|3|1 _PG5_01|_DFF_GG|A3 _PG5_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_GG|3|P _PG5_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG5_01|_DFF_GG|3|B _PG5_01|_DFF_GG|A3 _PG5_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_GG|3|RB _PG5_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_GG|4|1 _PG5_01|_DFF_GG|A4 _PG5_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_GG|4|P _PG5_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG5_01|_DFF_GG|4|B _PG5_01|_DFF_GG|A4 _PG5_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_GG|4|RB _PG5_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_GG|T|1 _PG5_01|_DFF_GG|T1 _PG5_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_GG|T|P _PG5_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG5_01|_DFF_GG|T|B _PG5_01|_DFF_GG|T1 _PG5_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_GG|T|RB _PG5_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_DFF_GG|45|1 _PG5_01|_DFF_GG|T2 _PG5_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG5_01|_DFF_GG|45|B _PG5_01|_DFF_GG|T2 _PG5_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG5_01|_DFF_GG|45|RB _PG5_01|_DFF_GG|45|MID_SHUNT _PG5_01|_DFF_GG|A4  2.1704737578552e-12
B_PG5_01|_DFF_GG|6|1 _PG5_01|_DFF_GG|Q1 _PG5_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_DFF_GG|6|P _PG5_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG5_01|_DFF_GG|6|B _PG5_01|_DFF_GG|Q1 _PG5_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG5_01|_DFF_GG|6|RB _PG5_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_AND_G|I_A1|B _PG5_01|_AND_G|A1 _PG5_01|_AND_G|I_A1|MID  2e-12
I_PG5_01|_AND_G|I_A1|B 0 _PG5_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_AND_G|I_B1|B _PG5_01|_AND_G|B1 _PG5_01|_AND_G|I_B1|MID  2e-12
I_PG5_01|_AND_G|I_B1|B 0 _PG5_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_AND_G|I_Q3|B _PG5_01|_AND_G|Q3 _PG5_01|_AND_G|I_Q3|MID  2e-12
I_PG5_01|_AND_G|I_Q3|B 0 _PG5_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG5_01|_AND_G|I_Q2|B _PG5_01|_AND_G|Q2 _PG5_01|_AND_G|I_Q2|MID  2e-12
I_PG5_01|_AND_G|I_Q2|B 0 _PG5_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_AND_G|I_Q1|B _PG5_01|_AND_G|Q1 _PG5_01|_AND_G|I_Q1|MID  2e-12
I_PG5_01|_AND_G|I_Q1|B 0 _PG5_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_AND_G|A1|1 _PG5_01|_AND_G|A1 _PG5_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_G|A1|P _PG5_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG5_01|_AND_G|A1|B _PG5_01|_AND_G|A1 _PG5_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG5_01|_AND_G|A1|RB _PG5_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_G|A2|1 _PG5_01|_AND_G|A2 _PG5_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_G|A2|P _PG5_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG5_01|_AND_G|A2|B _PG5_01|_AND_G|A2 _PG5_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG5_01|_AND_G|A2|RB _PG5_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_G|A12|1 _PG5_01|_AND_G|A2 _PG5_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_AND_G|A12|B _PG5_01|_AND_G|A2 _PG5_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG5_01|_AND_G|A12|RB _PG5_01|_AND_G|A12|MID_SHUNT _PG5_01|_AND_G|A3  2.1704737578552e-12
B_PG5_01|_AND_G|B1|1 _PG5_01|_AND_G|B1 _PG5_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_G|B1|P _PG5_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG5_01|_AND_G|B1|B _PG5_01|_AND_G|B1 _PG5_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG5_01|_AND_G|B1|RB _PG5_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_G|B2|1 _PG5_01|_AND_G|B2 _PG5_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_G|B2|P _PG5_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG5_01|_AND_G|B2|B _PG5_01|_AND_G|B2 _PG5_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG5_01|_AND_G|B2|RB _PG5_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_G|B12|1 _PG5_01|_AND_G|B2 _PG5_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG5_01|_AND_G|B12|B _PG5_01|_AND_G|B2 _PG5_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG5_01|_AND_G|B12|RB _PG5_01|_AND_G|B12|MID_SHUNT _PG5_01|_AND_G|B3  2.1704737578552e-12
B_PG5_01|_AND_G|Q2|1 _PG5_01|_AND_G|Q2 _PG5_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_G|Q2|P _PG5_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG5_01|_AND_G|Q2|B _PG5_01|_AND_G|Q2 _PG5_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG5_01|_AND_G|Q2|RB _PG5_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_G|Q1|1 _PG5_01|_AND_G|Q1 _PG5_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_G|Q1|P _PG5_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG5_01|_AND_G|Q1|B _PG5_01|_AND_G|Q1 _PG5_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG5_01|_AND_G|Q1|RB _PG5_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_01|_AND_P|I_A1|B _PG5_01|_AND_P|A1 _PG5_01|_AND_P|I_A1|MID  2e-12
I_PG5_01|_AND_P|I_A1|B 0 _PG5_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_AND_P|I_B1|B _PG5_01|_AND_P|B1 _PG5_01|_AND_P|I_B1|MID  2e-12
I_PG5_01|_AND_P|I_B1|B 0 _PG5_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_AND_P|I_Q3|B _PG5_01|_AND_P|Q3 _PG5_01|_AND_P|I_Q3|MID  2e-12
I_PG5_01|_AND_P|I_Q3|B 0 _PG5_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG5_01|_AND_P|I_Q2|B _PG5_01|_AND_P|Q2 _PG5_01|_AND_P|I_Q2|MID  2e-12
I_PG5_01|_AND_P|I_Q2|B 0 _PG5_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_01|_AND_P|I_Q1|B _PG5_01|_AND_P|Q1 _PG5_01|_AND_P|I_Q1|MID  2e-12
I_PG5_01|_AND_P|I_Q1|B 0 _PG5_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_01|_AND_P|A1|1 _PG5_01|_AND_P|A1 _PG5_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_P|A1|P _PG5_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG5_01|_AND_P|A1|B _PG5_01|_AND_P|A1 _PG5_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG5_01|_AND_P|A1|RB _PG5_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_P|A2|1 _PG5_01|_AND_P|A2 _PG5_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_P|A2|P _PG5_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG5_01|_AND_P|A2|B _PG5_01|_AND_P|A2 _PG5_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG5_01|_AND_P|A2|RB _PG5_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_P|A12|1 _PG5_01|_AND_P|A2 _PG5_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG5_01|_AND_P|A12|B _PG5_01|_AND_P|A2 _PG5_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG5_01|_AND_P|A12|RB _PG5_01|_AND_P|A12|MID_SHUNT _PG5_01|_AND_P|A3  2.1704737578552e-12
B_PG5_01|_AND_P|B1|1 _PG5_01|_AND_P|B1 _PG5_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_P|B1|P _PG5_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG5_01|_AND_P|B1|B _PG5_01|_AND_P|B1 _PG5_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG5_01|_AND_P|B1|RB _PG5_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_P|B2|1 _PG5_01|_AND_P|B2 _PG5_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_P|B2|P _PG5_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG5_01|_AND_P|B2|B _PG5_01|_AND_P|B2 _PG5_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG5_01|_AND_P|B2|RB _PG5_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_P|B12|1 _PG5_01|_AND_P|B2 _PG5_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG5_01|_AND_P|B12|B _PG5_01|_AND_P|B2 _PG5_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG5_01|_AND_P|B12|RB _PG5_01|_AND_P|B12|MID_SHUNT _PG5_01|_AND_P|B3  2.1704737578552e-12
B_PG5_01|_AND_P|Q2|1 _PG5_01|_AND_P|Q2 _PG5_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_P|Q2|P _PG5_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG5_01|_AND_P|Q2|B _PG5_01|_AND_P|Q2 _PG5_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG5_01|_AND_P|Q2|RB _PG5_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_01|_AND_P|Q1|1 _PG5_01|_AND_P|Q1 _PG5_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_01|_AND_P|Q1|P _PG5_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG5_01|_AND_P|Q1|B _PG5_01|_AND_P|Q1 _PG5_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG5_01|_AND_P|Q1|RB _PG5_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG6_01|P|I_1|B _PG6_01|P|A1 _PG6_01|P|I_1|MID  2e-12
I_PG6_01|P|I_1|B 0 _PG6_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_01|P|I_3|B _PG6_01|P|A3 _PG6_01|P|I_3|MID  2e-12
I_PG6_01|P|I_3|B 0 _PG6_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_01|P|I_T|B _PG6_01|P|T1 _PG6_01|P|I_T|MID  2e-12
I_PG6_01|P|I_T|B 0 _PG6_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_01|P|I_6|B _PG6_01|P|Q1 _PG6_01|P|I_6|MID  2e-12
I_PG6_01|P|I_6|B 0 _PG6_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_01|P|1|1 _PG6_01|P|A1 _PG6_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG6_01|P|1|P _PG6_01|P|1|MID_SERIES 0  2e-13
R_PG6_01|P|1|B _PG6_01|P|A1 _PG6_01|P|1|MID_SHUNT  2.7439617672
L_PG6_01|P|1|RB _PG6_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|P|23|1 _PG6_01|P|A2 _PG6_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG6_01|P|23|B _PG6_01|P|A2 _PG6_01|P|23|MID_SHUNT  3.84154647408
L_PG6_01|P|23|RB _PG6_01|P|23|MID_SHUNT _PG6_01|P|A3  2.1704737578552e-12
B_PG6_01|P|3|1 _PG6_01|P|A3 _PG6_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG6_01|P|3|P _PG6_01|P|3|MID_SERIES 0  2e-13
R_PG6_01|P|3|B _PG6_01|P|A3 _PG6_01|P|3|MID_SHUNT  2.7439617672
L_PG6_01|P|3|RB _PG6_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|P|4|1 _PG6_01|P|A4 _PG6_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG6_01|P|4|P _PG6_01|P|4|MID_SERIES 0  2e-13
R_PG6_01|P|4|B _PG6_01|P|A4 _PG6_01|P|4|MID_SHUNT  2.7439617672
L_PG6_01|P|4|RB _PG6_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|P|T|1 _PG6_01|P|T1 _PG6_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG6_01|P|T|P _PG6_01|P|T|MID_SERIES 0  2e-13
R_PG6_01|P|T|B _PG6_01|P|T1 _PG6_01|P|T|MID_SHUNT  2.7439617672
L_PG6_01|P|T|RB _PG6_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|P|45|1 _PG6_01|P|T2 _PG6_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG6_01|P|45|B _PG6_01|P|T2 _PG6_01|P|45|MID_SHUNT  3.84154647408
L_PG6_01|P|45|RB _PG6_01|P|45|MID_SHUNT _PG6_01|P|A4  2.1704737578552e-12
B_PG6_01|P|6|1 _PG6_01|P|Q1 _PG6_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG6_01|P|6|P _PG6_01|P|6|MID_SERIES 0  2e-13
R_PG6_01|P|6|B _PG6_01|P|Q1 _PG6_01|P|6|MID_SHUNT  2.7439617672
L_PG6_01|P|6|RB _PG6_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_01|G|I_1|B _PG6_01|G|A1 _PG6_01|G|I_1|MID  2e-12
I_PG6_01|G|I_1|B 0 _PG6_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_01|G|I_3|B _PG6_01|G|A3 _PG6_01|G|I_3|MID  2e-12
I_PG6_01|G|I_3|B 0 _PG6_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_01|G|I_T|B _PG6_01|G|T1 _PG6_01|G|I_T|MID  2e-12
I_PG6_01|G|I_T|B 0 _PG6_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_01|G|I_6|B _PG6_01|G|Q1 _PG6_01|G|I_6|MID  2e-12
I_PG6_01|G|I_6|B 0 _PG6_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_01|G|1|1 _PG6_01|G|A1 _PG6_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG6_01|G|1|P _PG6_01|G|1|MID_SERIES 0  2e-13
R_PG6_01|G|1|B _PG6_01|G|A1 _PG6_01|G|1|MID_SHUNT  2.7439617672
L_PG6_01|G|1|RB _PG6_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|G|23|1 _PG6_01|G|A2 _PG6_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG6_01|G|23|B _PG6_01|G|A2 _PG6_01|G|23|MID_SHUNT  3.84154647408
L_PG6_01|G|23|RB _PG6_01|G|23|MID_SHUNT _PG6_01|G|A3  2.1704737578552e-12
B_PG6_01|G|3|1 _PG6_01|G|A3 _PG6_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG6_01|G|3|P _PG6_01|G|3|MID_SERIES 0  2e-13
R_PG6_01|G|3|B _PG6_01|G|A3 _PG6_01|G|3|MID_SHUNT  2.7439617672
L_PG6_01|G|3|RB _PG6_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|G|4|1 _PG6_01|G|A4 _PG6_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG6_01|G|4|P _PG6_01|G|4|MID_SERIES 0  2e-13
R_PG6_01|G|4|B _PG6_01|G|A4 _PG6_01|G|4|MID_SHUNT  2.7439617672
L_PG6_01|G|4|RB _PG6_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|G|T|1 _PG6_01|G|T1 _PG6_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG6_01|G|T|P _PG6_01|G|T|MID_SERIES 0  2e-13
R_PG6_01|G|T|B _PG6_01|G|T1 _PG6_01|G|T|MID_SHUNT  2.7439617672
L_PG6_01|G|T|RB _PG6_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_01|G|45|1 _PG6_01|G|T2 _PG6_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG6_01|G|45|B _PG6_01|G|T2 _PG6_01|G|45|MID_SHUNT  3.84154647408
L_PG6_01|G|45|RB _PG6_01|G|45|MID_SHUNT _PG6_01|G|A4  2.1704737578552e-12
B_PG6_01|G|6|1 _PG6_01|G|Q1 _PG6_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG6_01|G|6|P _PG6_01|G|6|MID_SERIES 0  2e-13
R_PG6_01|G|6|B _PG6_01|G|Q1 _PG6_01|G|6|MID_SHUNT  2.7439617672
L_PG6_01|G|6|RB _PG6_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_SPL_G1|I_D1|B _PG7_01|_SPL_G1|D1 _PG7_01|_SPL_G1|I_D1|MID  2e-12
I_PG7_01|_SPL_G1|I_D1|B 0 _PG7_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_01|_SPL_G1|I_D2|B _PG7_01|_SPL_G1|D2 _PG7_01|_SPL_G1|I_D2|MID  2e-12
I_PG7_01|_SPL_G1|I_D2|B 0 _PG7_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG7_01|_SPL_G1|I_Q1|B _PG7_01|_SPL_G1|QA1 _PG7_01|_SPL_G1|I_Q1|MID  2e-12
I_PG7_01|_SPL_G1|I_Q1|B 0 _PG7_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_01|_SPL_G1|I_Q2|B _PG7_01|_SPL_G1|QB1 _PG7_01|_SPL_G1|I_Q2|MID  2e-12
I_PG7_01|_SPL_G1|I_Q2|B 0 _PG7_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG7_01|_SPL_G1|1|1 _PG7_01|_SPL_G1|D1 _PG7_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_G1|1|P _PG7_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG7_01|_SPL_G1|1|B _PG7_01|_SPL_G1|D1 _PG7_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_G1|1|RB _PG7_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_SPL_G1|2|1 _PG7_01|_SPL_G1|D2 _PG7_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_G1|2|P _PG7_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG7_01|_SPL_G1|2|B _PG7_01|_SPL_G1|D2 _PG7_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_G1|2|RB _PG7_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_SPL_G1|A|1 _PG7_01|_SPL_G1|QA1 _PG7_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_G1|A|P _PG7_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG7_01|_SPL_G1|A|B _PG7_01|_SPL_G1|QA1 _PG7_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_G1|A|RB _PG7_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_SPL_G1|B|1 _PG7_01|_SPL_G1|QB1 _PG7_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_G1|B|P _PG7_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG7_01|_SPL_G1|B|B _PG7_01|_SPL_G1|QB1 _PG7_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_G1|B|RB _PG7_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_SPL_P1|I_D1|B _PG7_01|_SPL_P1|D1 _PG7_01|_SPL_P1|I_D1|MID  2e-12
I_PG7_01|_SPL_P1|I_D1|B 0 _PG7_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_01|_SPL_P1|I_D2|B _PG7_01|_SPL_P1|D2 _PG7_01|_SPL_P1|I_D2|MID  2e-12
I_PG7_01|_SPL_P1|I_D2|B 0 _PG7_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG7_01|_SPL_P1|I_Q1|B _PG7_01|_SPL_P1|QA1 _PG7_01|_SPL_P1|I_Q1|MID  2e-12
I_PG7_01|_SPL_P1|I_Q1|B 0 _PG7_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_01|_SPL_P1|I_Q2|B _PG7_01|_SPL_P1|QB1 _PG7_01|_SPL_P1|I_Q2|MID  2e-12
I_PG7_01|_SPL_P1|I_Q2|B 0 _PG7_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG7_01|_SPL_P1|1|1 _PG7_01|_SPL_P1|D1 _PG7_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_P1|1|P _PG7_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG7_01|_SPL_P1|1|B _PG7_01|_SPL_P1|D1 _PG7_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_P1|1|RB _PG7_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_SPL_P1|2|1 _PG7_01|_SPL_P1|D2 _PG7_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_P1|2|P _PG7_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG7_01|_SPL_P1|2|B _PG7_01|_SPL_P1|D2 _PG7_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_P1|2|RB _PG7_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_SPL_P1|A|1 _PG7_01|_SPL_P1|QA1 _PG7_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_P1|A|P _PG7_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG7_01|_SPL_P1|A|B _PG7_01|_SPL_P1|QA1 _PG7_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_P1|A|RB _PG7_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_SPL_P1|B|1 _PG7_01|_SPL_P1|QB1 _PG7_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_SPL_P1|B|P _PG7_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG7_01|_SPL_P1|B|B _PG7_01|_SPL_P1|QB1 _PG7_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG7_01|_SPL_P1|B|RB _PG7_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_PG|I_A1|B _PG7_01|_PG|A1 _PG7_01|_PG|I_A1|MID  2e-12
I_PG7_01|_PG|I_A1|B 0 _PG7_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_PG|I_B1|B _PG7_01|_PG|B1 _PG7_01|_PG|I_B1|MID  2e-12
I_PG7_01|_PG|I_B1|B 0 _PG7_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_PG|I_Q3|B _PG7_01|_PG|Q3 _PG7_01|_PG|I_Q3|MID  2e-12
I_PG7_01|_PG|I_Q3|B 0 _PG7_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_01|_PG|I_Q2|B _PG7_01|_PG|Q2 _PG7_01|_PG|I_Q2|MID  2e-12
I_PG7_01|_PG|I_Q2|B 0 _PG7_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_PG|I_Q1|B _PG7_01|_PG|Q1 _PG7_01|_PG|I_Q1|MID  2e-12
I_PG7_01|_PG|I_Q1|B 0 _PG7_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_PG|A1|1 _PG7_01|_PG|A1 _PG7_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_PG|A1|P _PG7_01|_PG|A1|MID_SERIES 0  2e-13
R_PG7_01|_PG|A1|B _PG7_01|_PG|A1 _PG7_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG7_01|_PG|A1|RB _PG7_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_PG|A2|1 _PG7_01|_PG|A2 _PG7_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_PG|A2|P _PG7_01|_PG|A2|MID_SERIES 0  2e-13
R_PG7_01|_PG|A2|B _PG7_01|_PG|A2 _PG7_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG7_01|_PG|A2|RB _PG7_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_PG|A12|1 _PG7_01|_PG|A2 _PG7_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_PG|A12|B _PG7_01|_PG|A2 _PG7_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG7_01|_PG|A12|RB _PG7_01|_PG|A12|MID_SHUNT _PG7_01|_PG|A3  2.1704737578552e-12
B_PG7_01|_PG|B1|1 _PG7_01|_PG|B1 _PG7_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_PG|B1|P _PG7_01|_PG|B1|MID_SERIES 0  2e-13
R_PG7_01|_PG|B1|B _PG7_01|_PG|B1 _PG7_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG7_01|_PG|B1|RB _PG7_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_PG|B2|1 _PG7_01|_PG|B2 _PG7_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_PG|B2|P _PG7_01|_PG|B2|MID_SERIES 0  2e-13
R_PG7_01|_PG|B2|B _PG7_01|_PG|B2 _PG7_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG7_01|_PG|B2|RB _PG7_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_PG|B12|1 _PG7_01|_PG|B2 _PG7_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG7_01|_PG|B12|B _PG7_01|_PG|B2 _PG7_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG7_01|_PG|B12|RB _PG7_01|_PG|B12|MID_SHUNT _PG7_01|_PG|B3  2.1704737578552e-12
B_PG7_01|_PG|Q2|1 _PG7_01|_PG|Q2 _PG7_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_PG|Q2|P _PG7_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG7_01|_PG|Q2|B _PG7_01|_PG|Q2 _PG7_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG7_01|_PG|Q2|RB _PG7_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_PG|Q1|1 _PG7_01|_PG|Q1 _PG7_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_PG|Q1|P _PG7_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG7_01|_PG|Q1|B _PG7_01|_PG|Q1 _PG7_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG7_01|_PG|Q1|RB _PG7_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_GG|I_A1|B _PG7_01|_GG|A1 _PG7_01|_GG|I_A1|MID  2e-12
I_PG7_01|_GG|I_A1|B 0 _PG7_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_GG|I_B1|B _PG7_01|_GG|B1 _PG7_01|_GG|I_B1|MID  2e-12
I_PG7_01|_GG|I_B1|B 0 _PG7_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_GG|I_Q3|B _PG7_01|_GG|Q3 _PG7_01|_GG|I_Q3|MID  2e-12
I_PG7_01|_GG|I_Q3|B 0 _PG7_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_01|_GG|I_Q2|B _PG7_01|_GG|Q2 _PG7_01|_GG|I_Q2|MID  2e-12
I_PG7_01|_GG|I_Q2|B 0 _PG7_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_GG|I_Q1|B _PG7_01|_GG|Q1 _PG7_01|_GG|I_Q1|MID  2e-12
I_PG7_01|_GG|I_Q1|B 0 _PG7_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_GG|A1|1 _PG7_01|_GG|A1 _PG7_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_GG|A1|P _PG7_01|_GG|A1|MID_SERIES 0  2e-13
R_PG7_01|_GG|A1|B _PG7_01|_GG|A1 _PG7_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG7_01|_GG|A1|RB _PG7_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_GG|A2|1 _PG7_01|_GG|A2 _PG7_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_GG|A2|P _PG7_01|_GG|A2|MID_SERIES 0  2e-13
R_PG7_01|_GG|A2|B _PG7_01|_GG|A2 _PG7_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG7_01|_GG|A2|RB _PG7_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_GG|A12|1 _PG7_01|_GG|A2 _PG7_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_GG|A12|B _PG7_01|_GG|A2 _PG7_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG7_01|_GG|A12|RB _PG7_01|_GG|A12|MID_SHUNT _PG7_01|_GG|A3  2.1704737578552e-12
B_PG7_01|_GG|B1|1 _PG7_01|_GG|B1 _PG7_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_GG|B1|P _PG7_01|_GG|B1|MID_SERIES 0  2e-13
R_PG7_01|_GG|B1|B _PG7_01|_GG|B1 _PG7_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG7_01|_GG|B1|RB _PG7_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_GG|B2|1 _PG7_01|_GG|B2 _PG7_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_GG|B2|P _PG7_01|_GG|B2|MID_SERIES 0  2e-13
R_PG7_01|_GG|B2|B _PG7_01|_GG|B2 _PG7_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG7_01|_GG|B2|RB _PG7_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_GG|B12|1 _PG7_01|_GG|B2 _PG7_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG7_01|_GG|B12|B _PG7_01|_GG|B2 _PG7_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG7_01|_GG|B12|RB _PG7_01|_GG|B12|MID_SHUNT _PG7_01|_GG|B3  2.1704737578552e-12
B_PG7_01|_GG|Q2|1 _PG7_01|_GG|Q2 _PG7_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_GG|Q2|P _PG7_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG7_01|_GG|Q2|B _PG7_01|_GG|Q2 _PG7_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG7_01|_GG|Q2|RB _PG7_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_GG|Q1|1 _PG7_01|_GG|Q1 _PG7_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_GG|Q1|P _PG7_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG7_01|_GG|Q1|B _PG7_01|_GG|Q1 _PG7_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG7_01|_GG|Q1|RB _PG7_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_DFF_P0|I_1|B _PG7_01|_DFF_P0|A1 _PG7_01|_DFF_P0|I_1|MID  2e-12
I_PG7_01|_DFF_P0|I_1|B 0 _PG7_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_P0|I_3|B _PG7_01|_DFF_P0|A3 _PG7_01|_DFF_P0|I_3|MID  2e-12
I_PG7_01|_DFF_P0|I_3|B 0 _PG7_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_01|_DFF_P0|I_T|B _PG7_01|_DFF_P0|T1 _PG7_01|_DFF_P0|I_T|MID  2e-12
I_PG7_01|_DFF_P0|I_T|B 0 _PG7_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_P0|I_6|B _PG7_01|_DFF_P0|Q1 _PG7_01|_DFF_P0|I_6|MID  2e-12
I_PG7_01|_DFF_P0|I_6|B 0 _PG7_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_DFF_P0|1|1 _PG7_01|_DFF_P0|A1 _PG7_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P0|1|P _PG7_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P0|1|B _PG7_01|_DFF_P0|A1 _PG7_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P0|1|RB _PG7_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P0|23|1 _PG7_01|_DFF_P0|A2 _PG7_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_P0|23|B _PG7_01|_DFF_P0|A2 _PG7_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_P0|23|RB _PG7_01|_DFF_P0|23|MID_SHUNT _PG7_01|_DFF_P0|A3  2.1704737578552e-12
B_PG7_01|_DFF_P0|3|1 _PG7_01|_DFF_P0|A3 _PG7_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P0|3|P _PG7_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P0|3|B _PG7_01|_DFF_P0|A3 _PG7_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P0|3|RB _PG7_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P0|4|1 _PG7_01|_DFF_P0|A4 _PG7_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P0|4|P _PG7_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P0|4|B _PG7_01|_DFF_P0|A4 _PG7_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P0|4|RB _PG7_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P0|T|1 _PG7_01|_DFF_P0|T1 _PG7_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P0|T|P _PG7_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P0|T|B _PG7_01|_DFF_P0|T1 _PG7_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P0|T|RB _PG7_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P0|45|1 _PG7_01|_DFF_P0|T2 _PG7_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_P0|45|B _PG7_01|_DFF_P0|T2 _PG7_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_P0|45|RB _PG7_01|_DFF_P0|45|MID_SHUNT _PG7_01|_DFF_P0|A4  2.1704737578552e-12
B_PG7_01|_DFF_P0|6|1 _PG7_01|_DFF_P0|Q1 _PG7_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P0|6|P _PG7_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P0|6|B _PG7_01|_DFF_P0|Q1 _PG7_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P0|6|RB _PG7_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_DFF_P1|I_1|B _PG7_01|_DFF_P1|A1 _PG7_01|_DFF_P1|I_1|MID  2e-12
I_PG7_01|_DFF_P1|I_1|B 0 _PG7_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_P1|I_3|B _PG7_01|_DFF_P1|A3 _PG7_01|_DFF_P1|I_3|MID  2e-12
I_PG7_01|_DFF_P1|I_3|B 0 _PG7_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_01|_DFF_P1|I_T|B _PG7_01|_DFF_P1|T1 _PG7_01|_DFF_P1|I_T|MID  2e-12
I_PG7_01|_DFF_P1|I_T|B 0 _PG7_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_P1|I_6|B _PG7_01|_DFF_P1|Q1 _PG7_01|_DFF_P1|I_6|MID  2e-12
I_PG7_01|_DFF_P1|I_6|B 0 _PG7_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_DFF_P1|1|1 _PG7_01|_DFF_P1|A1 _PG7_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P1|1|P _PG7_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P1|1|B _PG7_01|_DFF_P1|A1 _PG7_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P1|1|RB _PG7_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P1|23|1 _PG7_01|_DFF_P1|A2 _PG7_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_P1|23|B _PG7_01|_DFF_P1|A2 _PG7_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_P1|23|RB _PG7_01|_DFF_P1|23|MID_SHUNT _PG7_01|_DFF_P1|A3  2.1704737578552e-12
B_PG7_01|_DFF_P1|3|1 _PG7_01|_DFF_P1|A3 _PG7_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P1|3|P _PG7_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P1|3|B _PG7_01|_DFF_P1|A3 _PG7_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P1|3|RB _PG7_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P1|4|1 _PG7_01|_DFF_P1|A4 _PG7_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P1|4|P _PG7_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P1|4|B _PG7_01|_DFF_P1|A4 _PG7_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P1|4|RB _PG7_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P1|T|1 _PG7_01|_DFF_P1|T1 _PG7_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P1|T|P _PG7_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P1|T|B _PG7_01|_DFF_P1|T1 _PG7_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P1|T|RB _PG7_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_P1|45|1 _PG7_01|_DFF_P1|T2 _PG7_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_P1|45|B _PG7_01|_DFF_P1|T2 _PG7_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_P1|45|RB _PG7_01|_DFF_P1|45|MID_SHUNT _PG7_01|_DFF_P1|A4  2.1704737578552e-12
B_PG7_01|_DFF_P1|6|1 _PG7_01|_DFF_P1|Q1 _PG7_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_P1|6|P _PG7_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG7_01|_DFF_P1|6|B _PG7_01|_DFF_P1|Q1 _PG7_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_P1|6|RB _PG7_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_DFF_PG|I_1|B _PG7_01|_DFF_PG|A1 _PG7_01|_DFF_PG|I_1|MID  2e-12
I_PG7_01|_DFF_PG|I_1|B 0 _PG7_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_PG|I_3|B _PG7_01|_DFF_PG|A3 _PG7_01|_DFF_PG|I_3|MID  2e-12
I_PG7_01|_DFF_PG|I_3|B 0 _PG7_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_01|_DFF_PG|I_T|B _PG7_01|_DFF_PG|T1 _PG7_01|_DFF_PG|I_T|MID  2e-12
I_PG7_01|_DFF_PG|I_T|B 0 _PG7_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_PG|I_6|B _PG7_01|_DFF_PG|Q1 _PG7_01|_DFF_PG|I_6|MID  2e-12
I_PG7_01|_DFF_PG|I_6|B 0 _PG7_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_DFF_PG|1|1 _PG7_01|_DFF_PG|A1 _PG7_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_PG|1|P _PG7_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG7_01|_DFF_PG|1|B _PG7_01|_DFF_PG|A1 _PG7_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_PG|1|RB _PG7_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_PG|23|1 _PG7_01|_DFF_PG|A2 _PG7_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_PG|23|B _PG7_01|_DFF_PG|A2 _PG7_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_PG|23|RB _PG7_01|_DFF_PG|23|MID_SHUNT _PG7_01|_DFF_PG|A3  2.1704737578552e-12
B_PG7_01|_DFF_PG|3|1 _PG7_01|_DFF_PG|A3 _PG7_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_PG|3|P _PG7_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG7_01|_DFF_PG|3|B _PG7_01|_DFF_PG|A3 _PG7_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_PG|3|RB _PG7_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_PG|4|1 _PG7_01|_DFF_PG|A4 _PG7_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_PG|4|P _PG7_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG7_01|_DFF_PG|4|B _PG7_01|_DFF_PG|A4 _PG7_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_PG|4|RB _PG7_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_PG|T|1 _PG7_01|_DFF_PG|T1 _PG7_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_PG|T|P _PG7_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG7_01|_DFF_PG|T|B _PG7_01|_DFF_PG|T1 _PG7_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_PG|T|RB _PG7_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_PG|45|1 _PG7_01|_DFF_PG|T2 _PG7_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_PG|45|B _PG7_01|_DFF_PG|T2 _PG7_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_PG|45|RB _PG7_01|_DFF_PG|45|MID_SHUNT _PG7_01|_DFF_PG|A4  2.1704737578552e-12
B_PG7_01|_DFF_PG|6|1 _PG7_01|_DFF_PG|Q1 _PG7_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_PG|6|P _PG7_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG7_01|_DFF_PG|6|B _PG7_01|_DFF_PG|Q1 _PG7_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_PG|6|RB _PG7_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_DFF_GG|I_1|B _PG7_01|_DFF_GG|A1 _PG7_01|_DFF_GG|I_1|MID  2e-12
I_PG7_01|_DFF_GG|I_1|B 0 _PG7_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_GG|I_3|B _PG7_01|_DFF_GG|A3 _PG7_01|_DFF_GG|I_3|MID  2e-12
I_PG7_01|_DFF_GG|I_3|B 0 _PG7_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_01|_DFF_GG|I_T|B _PG7_01|_DFF_GG|T1 _PG7_01|_DFF_GG|I_T|MID  2e-12
I_PG7_01|_DFF_GG|I_T|B 0 _PG7_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_DFF_GG|I_6|B _PG7_01|_DFF_GG|Q1 _PG7_01|_DFF_GG|I_6|MID  2e-12
I_PG7_01|_DFF_GG|I_6|B 0 _PG7_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_DFF_GG|1|1 _PG7_01|_DFF_GG|A1 _PG7_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_GG|1|P _PG7_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG7_01|_DFF_GG|1|B _PG7_01|_DFF_GG|A1 _PG7_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_GG|1|RB _PG7_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_GG|23|1 _PG7_01|_DFF_GG|A2 _PG7_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_GG|23|B _PG7_01|_DFF_GG|A2 _PG7_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_GG|23|RB _PG7_01|_DFF_GG|23|MID_SHUNT _PG7_01|_DFF_GG|A3  2.1704737578552e-12
B_PG7_01|_DFF_GG|3|1 _PG7_01|_DFF_GG|A3 _PG7_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_GG|3|P _PG7_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG7_01|_DFF_GG|3|B _PG7_01|_DFF_GG|A3 _PG7_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_GG|3|RB _PG7_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_GG|4|1 _PG7_01|_DFF_GG|A4 _PG7_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_GG|4|P _PG7_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG7_01|_DFF_GG|4|B _PG7_01|_DFF_GG|A4 _PG7_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_GG|4|RB _PG7_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_GG|T|1 _PG7_01|_DFF_GG|T1 _PG7_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_GG|T|P _PG7_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG7_01|_DFF_GG|T|B _PG7_01|_DFF_GG|T1 _PG7_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_GG|T|RB _PG7_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_DFF_GG|45|1 _PG7_01|_DFF_GG|T2 _PG7_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG7_01|_DFF_GG|45|B _PG7_01|_DFF_GG|T2 _PG7_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG7_01|_DFF_GG|45|RB _PG7_01|_DFF_GG|45|MID_SHUNT _PG7_01|_DFF_GG|A4  2.1704737578552e-12
B_PG7_01|_DFF_GG|6|1 _PG7_01|_DFF_GG|Q1 _PG7_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_DFF_GG|6|P _PG7_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG7_01|_DFF_GG|6|B _PG7_01|_DFF_GG|Q1 _PG7_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG7_01|_DFF_GG|6|RB _PG7_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_AND_G|I_A1|B _PG7_01|_AND_G|A1 _PG7_01|_AND_G|I_A1|MID  2e-12
I_PG7_01|_AND_G|I_A1|B 0 _PG7_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_AND_G|I_B1|B _PG7_01|_AND_G|B1 _PG7_01|_AND_G|I_B1|MID  2e-12
I_PG7_01|_AND_G|I_B1|B 0 _PG7_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_AND_G|I_Q3|B _PG7_01|_AND_G|Q3 _PG7_01|_AND_G|I_Q3|MID  2e-12
I_PG7_01|_AND_G|I_Q3|B 0 _PG7_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG7_01|_AND_G|I_Q2|B _PG7_01|_AND_G|Q2 _PG7_01|_AND_G|I_Q2|MID  2e-12
I_PG7_01|_AND_G|I_Q2|B 0 _PG7_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_AND_G|I_Q1|B _PG7_01|_AND_G|Q1 _PG7_01|_AND_G|I_Q1|MID  2e-12
I_PG7_01|_AND_G|I_Q1|B 0 _PG7_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_AND_G|A1|1 _PG7_01|_AND_G|A1 _PG7_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_G|A1|P _PG7_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG7_01|_AND_G|A1|B _PG7_01|_AND_G|A1 _PG7_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG7_01|_AND_G|A1|RB _PG7_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_G|A2|1 _PG7_01|_AND_G|A2 _PG7_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_G|A2|P _PG7_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG7_01|_AND_G|A2|B _PG7_01|_AND_G|A2 _PG7_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG7_01|_AND_G|A2|RB _PG7_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_G|A12|1 _PG7_01|_AND_G|A2 _PG7_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_AND_G|A12|B _PG7_01|_AND_G|A2 _PG7_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG7_01|_AND_G|A12|RB _PG7_01|_AND_G|A12|MID_SHUNT _PG7_01|_AND_G|A3  2.1704737578552e-12
B_PG7_01|_AND_G|B1|1 _PG7_01|_AND_G|B1 _PG7_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_G|B1|P _PG7_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG7_01|_AND_G|B1|B _PG7_01|_AND_G|B1 _PG7_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG7_01|_AND_G|B1|RB _PG7_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_G|B2|1 _PG7_01|_AND_G|B2 _PG7_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_G|B2|P _PG7_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG7_01|_AND_G|B2|B _PG7_01|_AND_G|B2 _PG7_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG7_01|_AND_G|B2|RB _PG7_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_G|B12|1 _PG7_01|_AND_G|B2 _PG7_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG7_01|_AND_G|B12|B _PG7_01|_AND_G|B2 _PG7_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG7_01|_AND_G|B12|RB _PG7_01|_AND_G|B12|MID_SHUNT _PG7_01|_AND_G|B3  2.1704737578552e-12
B_PG7_01|_AND_G|Q2|1 _PG7_01|_AND_G|Q2 _PG7_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_G|Q2|P _PG7_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG7_01|_AND_G|Q2|B _PG7_01|_AND_G|Q2 _PG7_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG7_01|_AND_G|Q2|RB _PG7_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_G|Q1|1 _PG7_01|_AND_G|Q1 _PG7_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_G|Q1|P _PG7_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG7_01|_AND_G|Q1|B _PG7_01|_AND_G|Q1 _PG7_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG7_01|_AND_G|Q1|RB _PG7_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_01|_AND_P|I_A1|B _PG7_01|_AND_P|A1 _PG7_01|_AND_P|I_A1|MID  2e-12
I_PG7_01|_AND_P|I_A1|B 0 _PG7_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_AND_P|I_B1|B _PG7_01|_AND_P|B1 _PG7_01|_AND_P|I_B1|MID  2e-12
I_PG7_01|_AND_P|I_B1|B 0 _PG7_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_AND_P|I_Q3|B _PG7_01|_AND_P|Q3 _PG7_01|_AND_P|I_Q3|MID  2e-12
I_PG7_01|_AND_P|I_Q3|B 0 _PG7_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG7_01|_AND_P|I_Q2|B _PG7_01|_AND_P|Q2 _PG7_01|_AND_P|I_Q2|MID  2e-12
I_PG7_01|_AND_P|I_Q2|B 0 _PG7_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_01|_AND_P|I_Q1|B _PG7_01|_AND_P|Q1 _PG7_01|_AND_P|I_Q1|MID  2e-12
I_PG7_01|_AND_P|I_Q1|B 0 _PG7_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_01|_AND_P|A1|1 _PG7_01|_AND_P|A1 _PG7_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_P|A1|P _PG7_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG7_01|_AND_P|A1|B _PG7_01|_AND_P|A1 _PG7_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG7_01|_AND_P|A1|RB _PG7_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_P|A2|1 _PG7_01|_AND_P|A2 _PG7_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_P|A2|P _PG7_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG7_01|_AND_P|A2|B _PG7_01|_AND_P|A2 _PG7_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG7_01|_AND_P|A2|RB _PG7_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_P|A12|1 _PG7_01|_AND_P|A2 _PG7_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG7_01|_AND_P|A12|B _PG7_01|_AND_P|A2 _PG7_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG7_01|_AND_P|A12|RB _PG7_01|_AND_P|A12|MID_SHUNT _PG7_01|_AND_P|A3  2.1704737578552e-12
B_PG7_01|_AND_P|B1|1 _PG7_01|_AND_P|B1 _PG7_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_P|B1|P _PG7_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG7_01|_AND_P|B1|B _PG7_01|_AND_P|B1 _PG7_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG7_01|_AND_P|B1|RB _PG7_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_P|B2|1 _PG7_01|_AND_P|B2 _PG7_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_P|B2|P _PG7_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG7_01|_AND_P|B2|B _PG7_01|_AND_P|B2 _PG7_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG7_01|_AND_P|B2|RB _PG7_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_P|B12|1 _PG7_01|_AND_P|B2 _PG7_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG7_01|_AND_P|B12|B _PG7_01|_AND_P|B2 _PG7_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG7_01|_AND_P|B12|RB _PG7_01|_AND_P|B12|MID_SHUNT _PG7_01|_AND_P|B3  2.1704737578552e-12
B_PG7_01|_AND_P|Q2|1 _PG7_01|_AND_P|Q2 _PG7_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_P|Q2|P _PG7_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG7_01|_AND_P|Q2|B _PG7_01|_AND_P|Q2 _PG7_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG7_01|_AND_P|Q2|RB _PG7_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_01|_AND_P|Q1|1 _PG7_01|_AND_P|Q1 _PG7_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_01|_AND_P|Q1|P _PG7_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG7_01|_AND_P|Q1|B _PG7_01|_AND_P|Q1 _PG7_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG7_01|_AND_P|Q1|RB _PG7_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PTL_P1_1|_SPL|I_D1|B _PTL_P1_1|_SPL|D1 _PTL_P1_1|_SPL|I_D1|MID  2e-12
I_PTL_P1_1|_SPL|I_D1|B 0 _PTL_P1_1|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P1_1|_SPL|I_D2|B _PTL_P1_1|_SPL|D2 _PTL_P1_1|_SPL|I_D2|MID  2e-12
I_PTL_P1_1|_SPL|I_D2|B 0 _PTL_P1_1|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P1_1|_SPL|I_Q1|B _PTL_P1_1|_SPL|QA1 _PTL_P1_1|_SPL|I_Q1|MID  2e-12
I_PTL_P1_1|_SPL|I_Q1|B 0 _PTL_P1_1|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P1_1|_SPL|I_Q2|B _PTL_P1_1|_SPL|QB1 _PTL_P1_1|_SPL|I_Q2|MID  2e-12
I_PTL_P1_1|_SPL|I_Q2|B 0 _PTL_P1_1|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P1_1|_SPL|1|1 _PTL_P1_1|_SPL|D1 _PTL_P1_1|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P1_1|_SPL|1|P _PTL_P1_1|_SPL|1|MID_SERIES 0  2e-13
R_PTL_P1_1|_SPL|1|B _PTL_P1_1|_SPL|D1 _PTL_P1_1|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_P1_1|_SPL|1|RB _PTL_P1_1|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P1_1|_SPL|2|1 _PTL_P1_1|_SPL|D2 _PTL_P1_1|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P1_1|_SPL|2|P _PTL_P1_1|_SPL|2|MID_SERIES 0  2e-13
R_PTL_P1_1|_SPL|2|B _PTL_P1_1|_SPL|D2 _PTL_P1_1|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_P1_1|_SPL|2|RB _PTL_P1_1|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P1_1|_SPL|A|1 _PTL_P1_1|_SPL|QA1 _PTL_P1_1|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P1_1|_SPL|A|P _PTL_P1_1|_SPL|A|MID_SERIES 0  2e-13
R_PTL_P1_1|_SPL|A|B _PTL_P1_1|_SPL|QA1 _PTL_P1_1|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_P1_1|_SPL|A|RB _PTL_P1_1|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P1_1|_SPL|B|1 _PTL_P1_1|_SPL|QB1 _PTL_P1_1|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P1_1|_SPL|B|P _PTL_P1_1|_SPL|B|MID_SERIES 0  2e-13
R_PTL_P1_1|_SPL|B|B _PTL_P1_1|_SPL|QB1 _PTL_P1_1|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_P1_1|_SPL|B|RB _PTL_P1_1|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_G1_1|_SPL|SPL1|1 _PTL_G1_1|D _PTL_G1_1|_SPL|SPL1|D1  2e-12
L_PTL_G1_1|_SPL|SPL1|2 _PTL_G1_1|_SPL|SPL1|D1 _PTL_G1_1|_SPL|SPL1|D2  4.135667696e-12
L_PTL_G1_1|_SPL|SPL1|3 _PTL_G1_1|_SPL|SPL1|D2 _PTL_G1_1|_SPL|SPL1|JCT  9.84682784761905e-13
L_PTL_G1_1|_SPL|SPL1|4 _PTL_G1_1|_SPL|SPL1|JCT _PTL_G1_1|_SPL|SPL1|QA1  9.84682784761905e-13
L_PTL_G1_1|_SPL|SPL1|5 _PTL_G1_1|_SPL|SPL1|QA1 G1_1_TO2  2e-12
L_PTL_G1_1|_SPL|SPL1|6 _PTL_G1_1|_SPL|SPL1|JCT _PTL_G1_1|_SPL|SPL1|QB1  9.84682784761905e-13
L_PTL_G1_1|_SPL|SPL1|7 _PTL_G1_1|_SPL|SPL1|QB1 _PTL_G1_1|_SPL|QTMP  2e-12
L_PTL_G1_1|_SPL|SPL2|1 _PTL_G1_1|_SPL|QTMP _PTL_G1_1|_SPL|SPL2|D1  2e-12
L_PTL_G1_1|_SPL|SPL2|2 _PTL_G1_1|_SPL|SPL2|D1 _PTL_G1_1|_SPL|SPL2|D2  4.135667696e-12
L_PTL_G1_1|_SPL|SPL2|3 _PTL_G1_1|_SPL|SPL2|D2 _PTL_G1_1|_SPL|SPL2|JCT  9.84682784761905e-13
L_PTL_G1_1|_SPL|SPL2|4 _PTL_G1_1|_SPL|SPL2|JCT _PTL_G1_1|_SPL|SPL2|QA1  9.84682784761905e-13
L_PTL_G1_1|_SPL|SPL2|5 _PTL_G1_1|_SPL|SPL2|QA1 G1_1_TO3  2e-12
L_PTL_G1_1|_SPL|SPL2|6 _PTL_G1_1|_SPL|SPL2|JCT _PTL_G1_1|_SPL|SPL2|QB1  9.84682784761905e-13
L_PTL_G1_1|_SPL|SPL2|7 _PTL_G1_1|_SPL|SPL2|QB1 G1_1_OUT  2e-12
L_PTL_P2_1|_SPL|I_D1|B _PTL_P2_1|_SPL|D1 _PTL_P2_1|_SPL|I_D1|MID  2e-12
I_PTL_P2_1|_SPL|I_D1|B 0 _PTL_P2_1|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_SPL|I_D2|B _PTL_P2_1|_SPL|D2 _PTL_P2_1|_SPL|I_D2|MID  2e-12
I_PTL_P2_1|_SPL|I_D2|B 0 _PTL_P2_1|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P2_1|_SPL|I_Q1|B _PTL_P2_1|_SPL|QA1 _PTL_P2_1|_SPL|I_Q1|MID  2e-12
I_PTL_P2_1|_SPL|I_Q1|B 0 _PTL_P2_1|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P2_1|_SPL|I_Q2|B _PTL_P2_1|_SPL|QB1 _PTL_P2_1|_SPL|I_Q2|MID  2e-12
I_PTL_P2_1|_SPL|I_Q2|B 0 _PTL_P2_1|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P2_1|_SPL|1|1 _PTL_P2_1|_SPL|D1 _PTL_P2_1|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P2_1|_SPL|1|P _PTL_P2_1|_SPL|1|MID_SERIES 0  2e-13
R_PTL_P2_1|_SPL|1|B _PTL_P2_1|_SPL|D1 _PTL_P2_1|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_P2_1|_SPL|1|RB _PTL_P2_1|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P2_1|_SPL|2|1 _PTL_P2_1|_SPL|D2 _PTL_P2_1|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P2_1|_SPL|2|P _PTL_P2_1|_SPL|2|MID_SERIES 0  2e-13
R_PTL_P2_1|_SPL|2|B _PTL_P2_1|_SPL|D2 _PTL_P2_1|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_P2_1|_SPL|2|RB _PTL_P2_1|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P2_1|_SPL|A|1 _PTL_P2_1|_SPL|QA1 _PTL_P2_1|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P2_1|_SPL|A|P _PTL_P2_1|_SPL|A|MID_SERIES 0  2e-13
R_PTL_P2_1|_SPL|A|B _PTL_P2_1|_SPL|QA1 _PTL_P2_1|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_P2_1|_SPL|A|RB _PTL_P2_1|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P2_1|_SPL|B|1 _PTL_P2_1|_SPL|QB1 _PTL_P2_1|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P2_1|_SPL|B|P _PTL_P2_1|_SPL|B|MID_SERIES 0  2e-13
R_PTL_P2_1|_SPL|B|B _PTL_P2_1|_SPL|QB1 _PTL_P2_1|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_P2_1|_SPL|B|RB _PTL_P2_1|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_P5_1|_SPL|I_D1|B _PTL_P5_1|_SPL|D1 _PTL_P5_1|_SPL|I_D1|MID  2e-12
I_PTL_P5_1|_SPL|I_D1|B 0 _PTL_P5_1|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P5_1|_SPL|I_D2|B _PTL_P5_1|_SPL|D2 _PTL_P5_1|_SPL|I_D2|MID  2e-12
I_PTL_P5_1|_SPL|I_D2|B 0 _PTL_P5_1|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P5_1|_SPL|I_Q1|B _PTL_P5_1|_SPL|QA1 _PTL_P5_1|_SPL|I_Q1|MID  2e-12
I_PTL_P5_1|_SPL|I_Q1|B 0 _PTL_P5_1|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P5_1|_SPL|I_Q2|B _PTL_P5_1|_SPL|QB1 _PTL_P5_1|_SPL|I_Q2|MID  2e-12
I_PTL_P5_1|_SPL|I_Q2|B 0 _PTL_P5_1|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P5_1|_SPL|1|1 _PTL_P5_1|_SPL|D1 _PTL_P5_1|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P5_1|_SPL|1|P _PTL_P5_1|_SPL|1|MID_SERIES 0  2e-13
R_PTL_P5_1|_SPL|1|B _PTL_P5_1|_SPL|D1 _PTL_P5_1|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_P5_1|_SPL|1|RB _PTL_P5_1|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P5_1|_SPL|2|1 _PTL_P5_1|_SPL|D2 _PTL_P5_1|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P5_1|_SPL|2|P _PTL_P5_1|_SPL|2|MID_SERIES 0  2e-13
R_PTL_P5_1|_SPL|2|B _PTL_P5_1|_SPL|D2 _PTL_P5_1|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_P5_1|_SPL|2|RB _PTL_P5_1|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P5_1|_SPL|A|1 _PTL_P5_1|_SPL|QA1 _PTL_P5_1|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P5_1|_SPL|A|P _PTL_P5_1|_SPL|A|MID_SERIES 0  2e-13
R_PTL_P5_1|_SPL|A|B _PTL_P5_1|_SPL|QA1 _PTL_P5_1|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_P5_1|_SPL|A|RB _PTL_P5_1|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P5_1|_SPL|B|1 _PTL_P5_1|_SPL|QB1 _PTL_P5_1|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P5_1|_SPL|B|P _PTL_P5_1|_SPL|B|MID_SERIES 0  2e-13
R_PTL_P5_1|_SPL|B|B _PTL_P5_1|_SPL|QB1 _PTL_P5_1|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_P5_1|_SPL|B|RB _PTL_P5_1|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_G5_1|_SPL|I_D1|B _PTL_G5_1|_SPL|D1 _PTL_G5_1|_SPL|I_D1|MID  2e-12
I_PTL_G5_1|_SPL|I_D1|B 0 _PTL_G5_1|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G5_1|_SPL|I_D2|B _PTL_G5_1|_SPL|D2 _PTL_G5_1|_SPL|I_D2|MID  2e-12
I_PTL_G5_1|_SPL|I_D2|B 0 _PTL_G5_1|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G5_1|_SPL|I_Q1|B _PTL_G5_1|_SPL|QA1 _PTL_G5_1|_SPL|I_Q1|MID  2e-12
I_PTL_G5_1|_SPL|I_Q1|B 0 _PTL_G5_1|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G5_1|_SPL|I_Q2|B _PTL_G5_1|_SPL|QB1 _PTL_G5_1|_SPL|I_Q2|MID  2e-12
I_PTL_G5_1|_SPL|I_Q2|B 0 _PTL_G5_1|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G5_1|_SPL|1|1 _PTL_G5_1|_SPL|D1 _PTL_G5_1|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_1|_SPL|1|P _PTL_G5_1|_SPL|1|MID_SERIES 0  2e-13
R_PTL_G5_1|_SPL|1|B _PTL_G5_1|_SPL|D1 _PTL_G5_1|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_G5_1|_SPL|1|RB _PTL_G5_1|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G5_1|_SPL|2|1 _PTL_G5_1|_SPL|D2 _PTL_G5_1|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_1|_SPL|2|P _PTL_G5_1|_SPL|2|MID_SERIES 0  2e-13
R_PTL_G5_1|_SPL|2|B _PTL_G5_1|_SPL|D2 _PTL_G5_1|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_G5_1|_SPL|2|RB _PTL_G5_1|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G5_1|_SPL|A|1 _PTL_G5_1|_SPL|QA1 _PTL_G5_1|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_1|_SPL|A|P _PTL_G5_1|_SPL|A|MID_SERIES 0  2e-13
R_PTL_G5_1|_SPL|A|B _PTL_G5_1|_SPL|QA1 _PTL_G5_1|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_G5_1|_SPL|A|RB _PTL_G5_1|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G5_1|_SPL|B|1 _PTL_G5_1|_SPL|QB1 _PTL_G5_1|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_1|_SPL|B|P _PTL_G5_1|_SPL|B|MID_SERIES 0  2e-13
R_PTL_G5_1|_SPL|B|B _PTL_G5_1|_SPL|QB1 _PTL_G5_1|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_G5_1|_SPL|B|RB _PTL_G5_1|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|I_D1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|I_D1|MID  2e-12
I_PG2_12|_SPL_G1|I_D1|B 0 _PG2_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_D2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|I_D2|MID  2e-12
I_PG2_12|_SPL_G1|I_D2|B 0 _PG2_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG2_12|_SPL_G1|I_Q1|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|I_Q1|MID  2e-12
I_PG2_12|_SPL_G1|I_Q1|B 0 _PG2_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_Q2|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|I_Q2|MID  2e-12
I_PG2_12|_SPL_G1|I_Q2|B 0 _PG2_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG2_12|_SPL_G1|1|1 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|1|P _PG2_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|1|RB _PG2_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|2|1 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|2|P _PG2_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|2|RB _PG2_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|A|1 _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|A|P _PG2_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|A|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|A|RB _PG2_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|B|1 _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|B|P _PG2_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|B|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|B|RB _PG2_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_P1|I_D1|B _PG2_12|_SPL_P1|D1 _PG2_12|_SPL_P1|I_D1|MID  2e-12
I_PG2_12|_SPL_P1|I_D1|B 0 _PG2_12|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_P1|I_D2|B _PG2_12|_SPL_P1|D2 _PG2_12|_SPL_P1|I_D2|MID  2e-12
I_PG2_12|_SPL_P1|I_D2|B 0 _PG2_12|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG2_12|_SPL_P1|I_Q1|B _PG2_12|_SPL_P1|QA1 _PG2_12|_SPL_P1|I_Q1|MID  2e-12
I_PG2_12|_SPL_P1|I_Q1|B 0 _PG2_12|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_P1|I_Q2|B _PG2_12|_SPL_P1|QB1 _PG2_12|_SPL_P1|I_Q2|MID  2e-12
I_PG2_12|_SPL_P1|I_Q2|B 0 _PG2_12|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG2_12|_SPL_P1|1|1 _PG2_12|_SPL_P1|D1 _PG2_12|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_P1|1|P _PG2_12|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG2_12|_SPL_P1|1|B _PG2_12|_SPL_P1|D1 _PG2_12|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_P1|1|RB _PG2_12|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_P1|2|1 _PG2_12|_SPL_P1|D2 _PG2_12|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_P1|2|P _PG2_12|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG2_12|_SPL_P1|2|B _PG2_12|_SPL_P1|D2 _PG2_12|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_P1|2|RB _PG2_12|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_P1|A|1 _PG2_12|_SPL_P1|QA1 _PG2_12|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_P1|A|P _PG2_12|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG2_12|_SPL_P1|A|B _PG2_12|_SPL_P1|QA1 _PG2_12|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_P1|A|RB _PG2_12|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_P1|B|1 _PG2_12|_SPL_P1|QB1 _PG2_12|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_P1|B|P _PG2_12|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG2_12|_SPL_P1|B|B _PG2_12|_SPL_P1|QB1 _PG2_12|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_P1|B|RB _PG2_12|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_PG|I_A1|B _PG2_12|_PG|A1 _PG2_12|_PG|I_A1|MID  2e-12
I_PG2_12|_PG|I_A1|B 0 _PG2_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_B1|B _PG2_12|_PG|B1 _PG2_12|_PG|I_B1|MID  2e-12
I_PG2_12|_PG|I_B1|B 0 _PG2_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q3|B _PG2_12|_PG|Q3 _PG2_12|_PG|I_Q3|MID  2e-12
I_PG2_12|_PG|I_Q3|B 0 _PG2_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_PG|I_Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|I_Q2|MID  2e-12
I_PG2_12|_PG|I_Q2|B 0 _PG2_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|I_Q1|MID  2e-12
I_PG2_12|_PG|I_Q1|B 0 _PG2_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_PG|A1|1 _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A1|P _PG2_12|_PG|A1|MID_SERIES 0  2e-13
R_PG2_12|_PG|A1|B _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A1|RB _PG2_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A2|1 _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A2|P _PG2_12|_PG|A2|MID_SERIES 0  2e-13
R_PG2_12|_PG|A2|B _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A2|RB _PG2_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A12|1 _PG2_12|_PG|A2 _PG2_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|A12|B _PG2_12|_PG|A2 _PG2_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|A12|RB _PG2_12|_PG|A12|MID_SHUNT _PG2_12|_PG|A3  2.1704737578552e-12
B_PG2_12|_PG|B1|1 _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B1|P _PG2_12|_PG|B1|MID_SERIES 0  2e-13
R_PG2_12|_PG|B1|B _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B1|RB _PG2_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B2|1 _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B2|P _PG2_12|_PG|B2|MID_SERIES 0  2e-13
R_PG2_12|_PG|B2|B _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B2|RB _PG2_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B12|1 _PG2_12|_PG|B2 _PG2_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|B12|B _PG2_12|_PG|B2 _PG2_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|B12|RB _PG2_12|_PG|B12|MID_SHUNT _PG2_12|_PG|B3  2.1704737578552e-12
B_PG2_12|_PG|Q2|1 _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q2|P _PG2_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q2|RB _PG2_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|Q1|1 _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q1|P _PG2_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q1|RB _PG2_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_GG|I_A1|B _PG2_12|_GG|A1 _PG2_12|_GG|I_A1|MID  2e-12
I_PG2_12|_GG|I_A1|B 0 _PG2_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_B1|B _PG2_12|_GG|B1 _PG2_12|_GG|I_B1|MID  2e-12
I_PG2_12|_GG|I_B1|B 0 _PG2_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q3|B _PG2_12|_GG|Q3 _PG2_12|_GG|I_Q3|MID  2e-12
I_PG2_12|_GG|I_Q3|B 0 _PG2_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_GG|I_Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|I_Q2|MID  2e-12
I_PG2_12|_GG|I_Q2|B 0 _PG2_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|I_Q1|MID  2e-12
I_PG2_12|_GG|I_Q1|B 0 _PG2_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_GG|A1|1 _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A1|P _PG2_12|_GG|A1|MID_SERIES 0  2e-13
R_PG2_12|_GG|A1|B _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A1|RB _PG2_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A2|1 _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A2|P _PG2_12|_GG|A2|MID_SERIES 0  2e-13
R_PG2_12|_GG|A2|B _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A2|RB _PG2_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A12|1 _PG2_12|_GG|A2 _PG2_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|A12|B _PG2_12|_GG|A2 _PG2_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|A12|RB _PG2_12|_GG|A12|MID_SHUNT _PG2_12|_GG|A3  2.1704737578552e-12
B_PG2_12|_GG|B1|1 _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B1|P _PG2_12|_GG|B1|MID_SERIES 0  2e-13
R_PG2_12|_GG|B1|B _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B1|RB _PG2_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B2|1 _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B2|P _PG2_12|_GG|B2|MID_SERIES 0  2e-13
R_PG2_12|_GG|B2|B _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B2|RB _PG2_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B12|1 _PG2_12|_GG|B2 _PG2_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|B12|B _PG2_12|_GG|B2 _PG2_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|B12|RB _PG2_12|_GG|B12|MID_SHUNT _PG2_12|_GG|B3  2.1704737578552e-12
B_PG2_12|_GG|Q2|1 _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q2|P _PG2_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q2|RB _PG2_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|Q1|1 _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q1|P _PG2_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q1|RB _PG2_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_P0|I_1|B _PG2_12|_DFF_P0|A1 _PG2_12|_DFF_P0|I_1|MID  2e-12
I_PG2_12|_DFF_P0|I_1|B 0 _PG2_12|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_P0|I_3|B _PG2_12|_DFF_P0|A3 _PG2_12|_DFF_P0|I_3|MID  2e-12
I_PG2_12|_DFF_P0|I_3|B 0 _PG2_12|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_P0|I_T|B _PG2_12|_DFF_P0|T1 _PG2_12|_DFF_P0|I_T|MID  2e-12
I_PG2_12|_DFF_P0|I_T|B 0 _PG2_12|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_P0|I_6|B _PG2_12|_DFF_P0|Q1 _PG2_12|_DFF_P0|I_6|MID  2e-12
I_PG2_12|_DFF_P0|I_6|B 0 _PG2_12|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_P0|1|1 _PG2_12|_DFF_P0|A1 _PG2_12|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P0|1|P _PG2_12|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P0|1|B _PG2_12|_DFF_P0|A1 _PG2_12|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P0|1|RB _PG2_12|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P0|23|1 _PG2_12|_DFF_P0|A2 _PG2_12|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_P0|23|B _PG2_12|_DFF_P0|A2 _PG2_12|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_P0|23|RB _PG2_12|_DFF_P0|23|MID_SHUNT _PG2_12|_DFF_P0|A3  2.1704737578552e-12
B_PG2_12|_DFF_P0|3|1 _PG2_12|_DFF_P0|A3 _PG2_12|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P0|3|P _PG2_12|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P0|3|B _PG2_12|_DFF_P0|A3 _PG2_12|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P0|3|RB _PG2_12|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P0|4|1 _PG2_12|_DFF_P0|A4 _PG2_12|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P0|4|P _PG2_12|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P0|4|B _PG2_12|_DFF_P0|A4 _PG2_12|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P0|4|RB _PG2_12|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P0|T|1 _PG2_12|_DFF_P0|T1 _PG2_12|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P0|T|P _PG2_12|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P0|T|B _PG2_12|_DFF_P0|T1 _PG2_12|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P0|T|RB _PG2_12|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P0|45|1 _PG2_12|_DFF_P0|T2 _PG2_12|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_P0|45|B _PG2_12|_DFF_P0|T2 _PG2_12|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_P0|45|RB _PG2_12|_DFF_P0|45|MID_SHUNT _PG2_12|_DFF_P0|A4  2.1704737578552e-12
B_PG2_12|_DFF_P0|6|1 _PG2_12|_DFF_P0|Q1 _PG2_12|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P0|6|P _PG2_12|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P0|6|B _PG2_12|_DFF_P0|Q1 _PG2_12|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P0|6|RB _PG2_12|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_P1|I_1|B _PG2_12|_DFF_P1|A1 _PG2_12|_DFF_P1|I_1|MID  2e-12
I_PG2_12|_DFF_P1|I_1|B 0 _PG2_12|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_P1|I_3|B _PG2_12|_DFF_P1|A3 _PG2_12|_DFF_P1|I_3|MID  2e-12
I_PG2_12|_DFF_P1|I_3|B 0 _PG2_12|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_P1|I_T|B _PG2_12|_DFF_P1|T1 _PG2_12|_DFF_P1|I_T|MID  2e-12
I_PG2_12|_DFF_P1|I_T|B 0 _PG2_12|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_P1|I_6|B _PG2_12|_DFF_P1|Q1 _PG2_12|_DFF_P1|I_6|MID  2e-12
I_PG2_12|_DFF_P1|I_6|B 0 _PG2_12|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_P1|1|1 _PG2_12|_DFF_P1|A1 _PG2_12|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P1|1|P _PG2_12|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P1|1|B _PG2_12|_DFF_P1|A1 _PG2_12|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P1|1|RB _PG2_12|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P1|23|1 _PG2_12|_DFF_P1|A2 _PG2_12|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_P1|23|B _PG2_12|_DFF_P1|A2 _PG2_12|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_P1|23|RB _PG2_12|_DFF_P1|23|MID_SHUNT _PG2_12|_DFF_P1|A3  2.1704737578552e-12
B_PG2_12|_DFF_P1|3|1 _PG2_12|_DFF_P1|A3 _PG2_12|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P1|3|P _PG2_12|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P1|3|B _PG2_12|_DFF_P1|A3 _PG2_12|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P1|3|RB _PG2_12|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P1|4|1 _PG2_12|_DFF_P1|A4 _PG2_12|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P1|4|P _PG2_12|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P1|4|B _PG2_12|_DFF_P1|A4 _PG2_12|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P1|4|RB _PG2_12|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P1|T|1 _PG2_12|_DFF_P1|T1 _PG2_12|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P1|T|P _PG2_12|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P1|T|B _PG2_12|_DFF_P1|T1 _PG2_12|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P1|T|RB _PG2_12|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_P1|45|1 _PG2_12|_DFF_P1|T2 _PG2_12|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_P1|45|B _PG2_12|_DFF_P1|T2 _PG2_12|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_P1|45|RB _PG2_12|_DFF_P1|45|MID_SHUNT _PG2_12|_DFF_P1|A4  2.1704737578552e-12
B_PG2_12|_DFF_P1|6|1 _PG2_12|_DFF_P1|Q1 _PG2_12|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_P1|6|P _PG2_12|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_P1|6|B _PG2_12|_DFF_P1|Q1 _PG2_12|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_P1|6|RB _PG2_12|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_PG|I_1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|I_1|MID  2e-12
I_PG2_12|_DFF_PG|I_1|B 0 _PG2_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|I_3|MID  2e-12
I_PG2_12|_DFF_PG|I_3|B 0 _PG2_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_PG|I_T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|I_T|MID  2e-12
I_PG2_12|_DFF_PG|I_T|B 0 _PG2_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|I_6|MID  2e-12
I_PG2_12|_DFF_PG|I_6|B 0 _PG2_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_PG|1|1 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|1|P _PG2_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|1|RB _PG2_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|23|1 _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|23|B _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|23|RB _PG2_12|_DFF_PG|23|MID_SHUNT _PG2_12|_DFF_PG|A3  2.1704737578552e-12
B_PG2_12|_DFF_PG|3|1 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|3|P _PG2_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|3|RB _PG2_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|4|1 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|4|P _PG2_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|4|B _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|4|RB _PG2_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|T|1 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|T|P _PG2_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|T|RB _PG2_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|45|1 _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|45|B _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|45|RB _PG2_12|_DFF_PG|45|MID_SHUNT _PG2_12|_DFF_PG|A4  2.1704737578552e-12
B_PG2_12|_DFF_PG|6|1 _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|6|P _PG2_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|6|RB _PG2_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_GG|I_1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|I_1|MID  2e-12
I_PG2_12|_DFF_GG|I_1|B 0 _PG2_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|I_3|MID  2e-12
I_PG2_12|_DFF_GG|I_3|B 0 _PG2_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_GG|I_T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|I_T|MID  2e-12
I_PG2_12|_DFF_GG|I_T|B 0 _PG2_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|I_6|MID  2e-12
I_PG2_12|_DFF_GG|I_6|B 0 _PG2_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_GG|1|1 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|1|P _PG2_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|1|RB _PG2_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|23|1 _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|23|B _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|23|RB _PG2_12|_DFF_GG|23|MID_SHUNT _PG2_12|_DFF_GG|A3  2.1704737578552e-12
B_PG2_12|_DFF_GG|3|1 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|3|P _PG2_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|3|RB _PG2_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|4|1 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|4|P _PG2_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|4|B _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|4|RB _PG2_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|T|1 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|T|P _PG2_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|T|RB _PG2_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|45|1 _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|45|B _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|45|RB _PG2_12|_DFF_GG|45|MID_SHUNT _PG2_12|_DFF_GG|A4  2.1704737578552e-12
B_PG2_12|_DFF_GG|6|1 _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|6|P _PG2_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|6|RB _PG2_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_G|I_A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|I_A1|MID  2e-12
I_PG2_12|_AND_G|I_A1|B 0 _PG2_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|I_B1|MID  2e-12
I_PG2_12|_AND_G|I_B1|B 0 _PG2_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q3|B _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|I_Q3|MID  2e-12
I_PG2_12|_AND_G|I_Q3|B 0 _PG2_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_G|I_Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|I_Q2|MID  2e-12
I_PG2_12|_AND_G|I_Q2|B 0 _PG2_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|I_Q1|MID  2e-12
I_PG2_12|_AND_G|I_Q1|B 0 _PG2_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_G|A1|1 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A1|P _PG2_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A1|RB _PG2_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A2|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A2|P _PG2_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A2|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A2|RB _PG2_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A12|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|A12|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|A12|RB _PG2_12|_AND_G|A12|MID_SHUNT _PG2_12|_AND_G|A3  2.1704737578552e-12
B_PG2_12|_AND_G|B1|1 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B1|P _PG2_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B1|RB _PG2_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B2|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B2|P _PG2_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B2|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B2|RB _PG2_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B12|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|B12|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|B12|RB _PG2_12|_AND_G|B12|MID_SHUNT _PG2_12|_AND_G|B3  2.1704737578552e-12
B_PG2_12|_AND_G|Q2|1 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q2|P _PG2_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q2|RB _PG2_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|Q1|1 _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q1|P _PG2_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q1|RB _PG2_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_P|I_A1|B _PG2_12|_AND_P|A1 _PG2_12|_AND_P|I_A1|MID  2e-12
I_PG2_12|_AND_P|I_A1|B 0 _PG2_12|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_P|I_B1|B _PG2_12|_AND_P|B1 _PG2_12|_AND_P|I_B1|MID  2e-12
I_PG2_12|_AND_P|I_B1|B 0 _PG2_12|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_P|I_Q3|B _PG2_12|_AND_P|Q3 _PG2_12|_AND_P|I_Q3|MID  2e-12
I_PG2_12|_AND_P|I_Q3|B 0 _PG2_12|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_P|I_Q2|B _PG2_12|_AND_P|Q2 _PG2_12|_AND_P|I_Q2|MID  2e-12
I_PG2_12|_AND_P|I_Q2|B 0 _PG2_12|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_P|I_Q1|B _PG2_12|_AND_P|Q1 _PG2_12|_AND_P|I_Q1|MID  2e-12
I_PG2_12|_AND_P|I_Q1|B 0 _PG2_12|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_P|A1|1 _PG2_12|_AND_P|A1 _PG2_12|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_P|A1|P _PG2_12|_AND_P|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_P|A1|B _PG2_12|_AND_P|A1 _PG2_12|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_P|A1|RB _PG2_12|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_P|A2|1 _PG2_12|_AND_P|A2 _PG2_12|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_P|A2|P _PG2_12|_AND_P|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_P|A2|B _PG2_12|_AND_P|A2 _PG2_12|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_P|A2|RB _PG2_12|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_P|A12|1 _PG2_12|_AND_P|A2 _PG2_12|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_P|A12|B _PG2_12|_AND_P|A2 _PG2_12|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_P|A12|RB _PG2_12|_AND_P|A12|MID_SHUNT _PG2_12|_AND_P|A3  2.1704737578552e-12
B_PG2_12|_AND_P|B1|1 _PG2_12|_AND_P|B1 _PG2_12|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_P|B1|P _PG2_12|_AND_P|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_P|B1|B _PG2_12|_AND_P|B1 _PG2_12|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_P|B1|RB _PG2_12|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_P|B2|1 _PG2_12|_AND_P|B2 _PG2_12|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_P|B2|P _PG2_12|_AND_P|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_P|B2|B _PG2_12|_AND_P|B2 _PG2_12|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_P|B2|RB _PG2_12|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_P|B12|1 _PG2_12|_AND_P|B2 _PG2_12|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_P|B12|B _PG2_12|_AND_P|B2 _PG2_12|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_P|B12|RB _PG2_12|_AND_P|B12|MID_SHUNT _PG2_12|_AND_P|B3  2.1704737578552e-12
B_PG2_12|_AND_P|Q2|1 _PG2_12|_AND_P|Q2 _PG2_12|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_P|Q2|P _PG2_12|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_P|Q2|B _PG2_12|_AND_P|Q2 _PG2_12|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_P|Q2|RB _PG2_12|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_P|Q1|1 _PG2_12|_AND_P|Q1 _PG2_12|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_P|Q1|P _PG2_12|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_P|Q1|B _PG2_12|_AND_P|Q1 _PG2_12|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_P|Q1|RB _PG2_12|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_SPL_G1|I_D1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|I_D1|MID  2e-12
I_PG3_12|_SPL_G1|I_D1|B 0 _PG3_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_D2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|I_D2|MID  2e-12
I_PG3_12|_SPL_G1|I_D2|B 0 _PG3_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_12|_SPL_G1|I_Q1|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|I_Q1|MID  2e-12
I_PG3_12|_SPL_G1|I_Q1|B 0 _PG3_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_Q2|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|I_Q2|MID  2e-12
I_PG3_12|_SPL_G1|I_Q2|B 0 _PG3_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_12|_SPL_G1|1|1 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|1|P _PG3_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|1|RB _PG3_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|2|1 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|2|P _PG3_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|2|RB _PG3_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|A|1 _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|A|P _PG3_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|A|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|A|RB _PG3_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|B|1 _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|B|P _PG3_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|B|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|B|RB _PG3_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_SPL_P1|I_D1|B _PG3_12|_SPL_P1|D1 _PG3_12|_SPL_P1|I_D1|MID  2e-12
I_PG3_12|_SPL_P1|I_D1|B 0 _PG3_12|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_P1|I_D2|B _PG3_12|_SPL_P1|D2 _PG3_12|_SPL_P1|I_D2|MID  2e-12
I_PG3_12|_SPL_P1|I_D2|B 0 _PG3_12|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_12|_SPL_P1|I_Q1|B _PG3_12|_SPL_P1|QA1 _PG3_12|_SPL_P1|I_Q1|MID  2e-12
I_PG3_12|_SPL_P1|I_Q1|B 0 _PG3_12|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_P1|I_Q2|B _PG3_12|_SPL_P1|QB1 _PG3_12|_SPL_P1|I_Q2|MID  2e-12
I_PG3_12|_SPL_P1|I_Q2|B 0 _PG3_12|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_12|_SPL_P1|1|1 _PG3_12|_SPL_P1|D1 _PG3_12|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_P1|1|P _PG3_12|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_12|_SPL_P1|1|B _PG3_12|_SPL_P1|D1 _PG3_12|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_P1|1|RB _PG3_12|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_P1|2|1 _PG3_12|_SPL_P1|D2 _PG3_12|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_P1|2|P _PG3_12|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_12|_SPL_P1|2|B _PG3_12|_SPL_P1|D2 _PG3_12|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_P1|2|RB _PG3_12|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_P1|A|1 _PG3_12|_SPL_P1|QA1 _PG3_12|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_P1|A|P _PG3_12|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_12|_SPL_P1|A|B _PG3_12|_SPL_P1|QA1 _PG3_12|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_P1|A|RB _PG3_12|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_P1|B|1 _PG3_12|_SPL_P1|QB1 _PG3_12|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_P1|B|P _PG3_12|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_12|_SPL_P1|B|B _PG3_12|_SPL_P1|QB1 _PG3_12|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_P1|B|RB _PG3_12|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_PG|I_A1|B _PG3_12|_PG|A1 _PG3_12|_PG|I_A1|MID  2e-12
I_PG3_12|_PG|I_A1|B 0 _PG3_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_B1|B _PG3_12|_PG|B1 _PG3_12|_PG|I_B1|MID  2e-12
I_PG3_12|_PG|I_B1|B 0 _PG3_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q3|B _PG3_12|_PG|Q3 _PG3_12|_PG|I_Q3|MID  2e-12
I_PG3_12|_PG|I_Q3|B 0 _PG3_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_PG|I_Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|I_Q2|MID  2e-12
I_PG3_12|_PG|I_Q2|B 0 _PG3_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|I_Q1|MID  2e-12
I_PG3_12|_PG|I_Q1|B 0 _PG3_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_PG|A1|1 _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A1|P _PG3_12|_PG|A1|MID_SERIES 0  2e-13
R_PG3_12|_PG|A1|B _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A1|RB _PG3_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A2|1 _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A2|P _PG3_12|_PG|A2|MID_SERIES 0  2e-13
R_PG3_12|_PG|A2|B _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A2|RB _PG3_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A12|1 _PG3_12|_PG|A2 _PG3_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|A12|B _PG3_12|_PG|A2 _PG3_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|A12|RB _PG3_12|_PG|A12|MID_SHUNT _PG3_12|_PG|A3  2.1704737578552e-12
B_PG3_12|_PG|B1|1 _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B1|P _PG3_12|_PG|B1|MID_SERIES 0  2e-13
R_PG3_12|_PG|B1|B _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B1|RB _PG3_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B2|1 _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B2|P _PG3_12|_PG|B2|MID_SERIES 0  2e-13
R_PG3_12|_PG|B2|B _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B2|RB _PG3_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B12|1 _PG3_12|_PG|B2 _PG3_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|B12|B _PG3_12|_PG|B2 _PG3_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|B12|RB _PG3_12|_PG|B12|MID_SHUNT _PG3_12|_PG|B3  2.1704737578552e-12
B_PG3_12|_PG|Q2|1 _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q2|P _PG3_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q2|RB _PG3_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|Q1|1 _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q1|P _PG3_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q1|RB _PG3_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_GG|I_A1|B _PG3_12|_GG|A1 _PG3_12|_GG|I_A1|MID  2e-12
I_PG3_12|_GG|I_A1|B 0 _PG3_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_B1|B _PG3_12|_GG|B1 _PG3_12|_GG|I_B1|MID  2e-12
I_PG3_12|_GG|I_B1|B 0 _PG3_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q3|B _PG3_12|_GG|Q3 _PG3_12|_GG|I_Q3|MID  2e-12
I_PG3_12|_GG|I_Q3|B 0 _PG3_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_GG|I_Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|I_Q2|MID  2e-12
I_PG3_12|_GG|I_Q2|B 0 _PG3_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|I_Q1|MID  2e-12
I_PG3_12|_GG|I_Q1|B 0 _PG3_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_GG|A1|1 _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A1|P _PG3_12|_GG|A1|MID_SERIES 0  2e-13
R_PG3_12|_GG|A1|B _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A1|RB _PG3_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A2|1 _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A2|P _PG3_12|_GG|A2|MID_SERIES 0  2e-13
R_PG3_12|_GG|A2|B _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A2|RB _PG3_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A12|1 _PG3_12|_GG|A2 _PG3_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|A12|B _PG3_12|_GG|A2 _PG3_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|A12|RB _PG3_12|_GG|A12|MID_SHUNT _PG3_12|_GG|A3  2.1704737578552e-12
B_PG3_12|_GG|B1|1 _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B1|P _PG3_12|_GG|B1|MID_SERIES 0  2e-13
R_PG3_12|_GG|B1|B _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B1|RB _PG3_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B2|1 _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B2|P _PG3_12|_GG|B2|MID_SERIES 0  2e-13
R_PG3_12|_GG|B2|B _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B2|RB _PG3_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B12|1 _PG3_12|_GG|B2 _PG3_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|B12|B _PG3_12|_GG|B2 _PG3_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|B12|RB _PG3_12|_GG|B12|MID_SHUNT _PG3_12|_GG|B3  2.1704737578552e-12
B_PG3_12|_GG|Q2|1 _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q2|P _PG3_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q2|RB _PG3_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|Q1|1 _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q1|P _PG3_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q1|RB _PG3_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_P0|I_1|B _PG3_12|_DFF_P0|A1 _PG3_12|_DFF_P0|I_1|MID  2e-12
I_PG3_12|_DFF_P0|I_1|B 0 _PG3_12|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_P0|I_3|B _PG3_12|_DFF_P0|A3 _PG3_12|_DFF_P0|I_3|MID  2e-12
I_PG3_12|_DFF_P0|I_3|B 0 _PG3_12|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_P0|I_T|B _PG3_12|_DFF_P0|T1 _PG3_12|_DFF_P0|I_T|MID  2e-12
I_PG3_12|_DFF_P0|I_T|B 0 _PG3_12|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_P0|I_6|B _PG3_12|_DFF_P0|Q1 _PG3_12|_DFF_P0|I_6|MID  2e-12
I_PG3_12|_DFF_P0|I_6|B 0 _PG3_12|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_P0|1|1 _PG3_12|_DFF_P0|A1 _PG3_12|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P0|1|P _PG3_12|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P0|1|B _PG3_12|_DFF_P0|A1 _PG3_12|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P0|1|RB _PG3_12|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P0|23|1 _PG3_12|_DFF_P0|A2 _PG3_12|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_P0|23|B _PG3_12|_DFF_P0|A2 _PG3_12|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_P0|23|RB _PG3_12|_DFF_P0|23|MID_SHUNT _PG3_12|_DFF_P0|A3  2.1704737578552e-12
B_PG3_12|_DFF_P0|3|1 _PG3_12|_DFF_P0|A3 _PG3_12|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P0|3|P _PG3_12|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P0|3|B _PG3_12|_DFF_P0|A3 _PG3_12|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P0|3|RB _PG3_12|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P0|4|1 _PG3_12|_DFF_P0|A4 _PG3_12|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P0|4|P _PG3_12|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P0|4|B _PG3_12|_DFF_P0|A4 _PG3_12|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P0|4|RB _PG3_12|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P0|T|1 _PG3_12|_DFF_P0|T1 _PG3_12|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P0|T|P _PG3_12|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P0|T|B _PG3_12|_DFF_P0|T1 _PG3_12|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P0|T|RB _PG3_12|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P0|45|1 _PG3_12|_DFF_P0|T2 _PG3_12|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_P0|45|B _PG3_12|_DFF_P0|T2 _PG3_12|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_P0|45|RB _PG3_12|_DFF_P0|45|MID_SHUNT _PG3_12|_DFF_P0|A4  2.1704737578552e-12
B_PG3_12|_DFF_P0|6|1 _PG3_12|_DFF_P0|Q1 _PG3_12|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P0|6|P _PG3_12|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P0|6|B _PG3_12|_DFF_P0|Q1 _PG3_12|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P0|6|RB _PG3_12|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_P1|I_1|B _PG3_12|_DFF_P1|A1 _PG3_12|_DFF_P1|I_1|MID  2e-12
I_PG3_12|_DFF_P1|I_1|B 0 _PG3_12|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_P1|I_3|B _PG3_12|_DFF_P1|A3 _PG3_12|_DFF_P1|I_3|MID  2e-12
I_PG3_12|_DFF_P1|I_3|B 0 _PG3_12|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_P1|I_T|B _PG3_12|_DFF_P1|T1 _PG3_12|_DFF_P1|I_T|MID  2e-12
I_PG3_12|_DFF_P1|I_T|B 0 _PG3_12|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_P1|I_6|B _PG3_12|_DFF_P1|Q1 _PG3_12|_DFF_P1|I_6|MID  2e-12
I_PG3_12|_DFF_P1|I_6|B 0 _PG3_12|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_P1|1|1 _PG3_12|_DFF_P1|A1 _PG3_12|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P1|1|P _PG3_12|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P1|1|B _PG3_12|_DFF_P1|A1 _PG3_12|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P1|1|RB _PG3_12|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P1|23|1 _PG3_12|_DFF_P1|A2 _PG3_12|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_P1|23|B _PG3_12|_DFF_P1|A2 _PG3_12|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_P1|23|RB _PG3_12|_DFF_P1|23|MID_SHUNT _PG3_12|_DFF_P1|A3  2.1704737578552e-12
B_PG3_12|_DFF_P1|3|1 _PG3_12|_DFF_P1|A3 _PG3_12|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P1|3|P _PG3_12|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P1|3|B _PG3_12|_DFF_P1|A3 _PG3_12|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P1|3|RB _PG3_12|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P1|4|1 _PG3_12|_DFF_P1|A4 _PG3_12|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P1|4|P _PG3_12|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P1|4|B _PG3_12|_DFF_P1|A4 _PG3_12|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P1|4|RB _PG3_12|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P1|T|1 _PG3_12|_DFF_P1|T1 _PG3_12|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P1|T|P _PG3_12|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P1|T|B _PG3_12|_DFF_P1|T1 _PG3_12|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P1|T|RB _PG3_12|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_P1|45|1 _PG3_12|_DFF_P1|T2 _PG3_12|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_P1|45|B _PG3_12|_DFF_P1|T2 _PG3_12|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_P1|45|RB _PG3_12|_DFF_P1|45|MID_SHUNT _PG3_12|_DFF_P1|A4  2.1704737578552e-12
B_PG3_12|_DFF_P1|6|1 _PG3_12|_DFF_P1|Q1 _PG3_12|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_P1|6|P _PG3_12|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_P1|6|B _PG3_12|_DFF_P1|Q1 _PG3_12|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_P1|6|RB _PG3_12|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_PG|I_1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|I_1|MID  2e-12
I_PG3_12|_DFF_PG|I_1|B 0 _PG3_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|I_3|MID  2e-12
I_PG3_12|_DFF_PG|I_3|B 0 _PG3_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_PG|I_T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|I_T|MID  2e-12
I_PG3_12|_DFF_PG|I_T|B 0 _PG3_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|I_6|MID  2e-12
I_PG3_12|_DFF_PG|I_6|B 0 _PG3_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_PG|1|1 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|1|P _PG3_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|1|RB _PG3_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|23|1 _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|23|B _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|23|RB _PG3_12|_DFF_PG|23|MID_SHUNT _PG3_12|_DFF_PG|A3  2.1704737578552e-12
B_PG3_12|_DFF_PG|3|1 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|3|P _PG3_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|3|RB _PG3_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|4|1 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|4|P _PG3_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|4|B _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|4|RB _PG3_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|T|1 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|T|P _PG3_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|T|RB _PG3_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|45|1 _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|45|B _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|45|RB _PG3_12|_DFF_PG|45|MID_SHUNT _PG3_12|_DFF_PG|A4  2.1704737578552e-12
B_PG3_12|_DFF_PG|6|1 _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|6|P _PG3_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|6|RB _PG3_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_GG|I_1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|I_1|MID  2e-12
I_PG3_12|_DFF_GG|I_1|B 0 _PG3_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|I_3|MID  2e-12
I_PG3_12|_DFF_GG|I_3|B 0 _PG3_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_GG|I_T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|I_T|MID  2e-12
I_PG3_12|_DFF_GG|I_T|B 0 _PG3_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|I_6|MID  2e-12
I_PG3_12|_DFF_GG|I_6|B 0 _PG3_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_GG|1|1 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|1|P _PG3_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|1|RB _PG3_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|23|1 _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|23|B _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|23|RB _PG3_12|_DFF_GG|23|MID_SHUNT _PG3_12|_DFF_GG|A3  2.1704737578552e-12
B_PG3_12|_DFF_GG|3|1 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|3|P _PG3_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|3|RB _PG3_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|4|1 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|4|P _PG3_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|4|B _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|4|RB _PG3_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|T|1 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|T|P _PG3_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|T|RB _PG3_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|45|1 _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|45|B _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|45|RB _PG3_12|_DFF_GG|45|MID_SHUNT _PG3_12|_DFF_GG|A4  2.1704737578552e-12
B_PG3_12|_DFF_GG|6|1 _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|6|P _PG3_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|6|RB _PG3_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_G|I_A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|I_A1|MID  2e-12
I_PG3_12|_AND_G|I_A1|B 0 _PG3_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|I_B1|MID  2e-12
I_PG3_12|_AND_G|I_B1|B 0 _PG3_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q3|B _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|I_Q3|MID  2e-12
I_PG3_12|_AND_G|I_Q3|B 0 _PG3_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_G|I_Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|I_Q2|MID  2e-12
I_PG3_12|_AND_G|I_Q2|B 0 _PG3_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|I_Q1|MID  2e-12
I_PG3_12|_AND_G|I_Q1|B 0 _PG3_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_G|A1|1 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A1|P _PG3_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A1|RB _PG3_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A2|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A2|P _PG3_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A2|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A2|RB _PG3_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A12|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|A12|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|A12|RB _PG3_12|_AND_G|A12|MID_SHUNT _PG3_12|_AND_G|A3  2.1704737578552e-12
B_PG3_12|_AND_G|B1|1 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B1|P _PG3_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B1|RB _PG3_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B2|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B2|P _PG3_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B2|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B2|RB _PG3_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B12|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|B12|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|B12|RB _PG3_12|_AND_G|B12|MID_SHUNT _PG3_12|_AND_G|B3  2.1704737578552e-12
B_PG3_12|_AND_G|Q2|1 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q2|P _PG3_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q2|RB _PG3_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|Q1|1 _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q1|P _PG3_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q1|RB _PG3_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_P|I_A1|B _PG3_12|_AND_P|A1 _PG3_12|_AND_P|I_A1|MID  2e-12
I_PG3_12|_AND_P|I_A1|B 0 _PG3_12|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_P|I_B1|B _PG3_12|_AND_P|B1 _PG3_12|_AND_P|I_B1|MID  2e-12
I_PG3_12|_AND_P|I_B1|B 0 _PG3_12|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_P|I_Q3|B _PG3_12|_AND_P|Q3 _PG3_12|_AND_P|I_Q3|MID  2e-12
I_PG3_12|_AND_P|I_Q3|B 0 _PG3_12|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_P|I_Q2|B _PG3_12|_AND_P|Q2 _PG3_12|_AND_P|I_Q2|MID  2e-12
I_PG3_12|_AND_P|I_Q2|B 0 _PG3_12|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_P|I_Q1|B _PG3_12|_AND_P|Q1 _PG3_12|_AND_P|I_Q1|MID  2e-12
I_PG3_12|_AND_P|I_Q1|B 0 _PG3_12|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_P|A1|1 _PG3_12|_AND_P|A1 _PG3_12|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_P|A1|P _PG3_12|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_P|A1|B _PG3_12|_AND_P|A1 _PG3_12|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_P|A1|RB _PG3_12|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_P|A2|1 _PG3_12|_AND_P|A2 _PG3_12|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_P|A2|P _PG3_12|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_P|A2|B _PG3_12|_AND_P|A2 _PG3_12|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_P|A2|RB _PG3_12|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_P|A12|1 _PG3_12|_AND_P|A2 _PG3_12|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_P|A12|B _PG3_12|_AND_P|A2 _PG3_12|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_P|A12|RB _PG3_12|_AND_P|A12|MID_SHUNT _PG3_12|_AND_P|A3  2.1704737578552e-12
B_PG3_12|_AND_P|B1|1 _PG3_12|_AND_P|B1 _PG3_12|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_P|B1|P _PG3_12|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_P|B1|B _PG3_12|_AND_P|B1 _PG3_12|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_P|B1|RB _PG3_12|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_P|B2|1 _PG3_12|_AND_P|B2 _PG3_12|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_P|B2|P _PG3_12|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_P|B2|B _PG3_12|_AND_P|B2 _PG3_12|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_P|B2|RB _PG3_12|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_P|B12|1 _PG3_12|_AND_P|B2 _PG3_12|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_P|B12|B _PG3_12|_AND_P|B2 _PG3_12|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_P|B12|RB _PG3_12|_AND_P|B12|MID_SHUNT _PG3_12|_AND_P|B3  2.1704737578552e-12
B_PG3_12|_AND_P|Q2|1 _PG3_12|_AND_P|Q2 _PG3_12|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_P|Q2|P _PG3_12|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_P|Q2|B _PG3_12|_AND_P|Q2 _PG3_12|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_P|Q2|RB _PG3_12|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_P|Q1|1 _PG3_12|_AND_P|Q1 _PG3_12|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_P|Q1|P _PG3_12|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_P|Q1|B _PG3_12|_AND_P|Q1 _PG3_12|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_P|Q1|RB _PG3_12|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG4_12|P|I_1|B _PG4_12|P|A1 _PG4_12|P|I_1|MID  2e-12
I_PG4_12|P|I_1|B 0 _PG4_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_12|P|I_3|B _PG4_12|P|A3 _PG4_12|P|I_3|MID  2e-12
I_PG4_12|P|I_3|B 0 _PG4_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_12|P|I_T|B _PG4_12|P|T1 _PG4_12|P|I_T|MID  2e-12
I_PG4_12|P|I_T|B 0 _PG4_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_12|P|I_6|B _PG4_12|P|Q1 _PG4_12|P|I_6|MID  2e-12
I_PG4_12|P|I_6|B 0 _PG4_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_12|P|1|1 _PG4_12|P|A1 _PG4_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG4_12|P|1|P _PG4_12|P|1|MID_SERIES 0  2e-13
R_PG4_12|P|1|B _PG4_12|P|A1 _PG4_12|P|1|MID_SHUNT  2.7439617672
L_PG4_12|P|1|RB _PG4_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|P|23|1 _PG4_12|P|A2 _PG4_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG4_12|P|23|B _PG4_12|P|A2 _PG4_12|P|23|MID_SHUNT  3.84154647408
L_PG4_12|P|23|RB _PG4_12|P|23|MID_SHUNT _PG4_12|P|A3  2.1704737578552e-12
B_PG4_12|P|3|1 _PG4_12|P|A3 _PG4_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG4_12|P|3|P _PG4_12|P|3|MID_SERIES 0  2e-13
R_PG4_12|P|3|B _PG4_12|P|A3 _PG4_12|P|3|MID_SHUNT  2.7439617672
L_PG4_12|P|3|RB _PG4_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|P|4|1 _PG4_12|P|A4 _PG4_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG4_12|P|4|P _PG4_12|P|4|MID_SERIES 0  2e-13
R_PG4_12|P|4|B _PG4_12|P|A4 _PG4_12|P|4|MID_SHUNT  2.7439617672
L_PG4_12|P|4|RB _PG4_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|P|T|1 _PG4_12|P|T1 _PG4_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG4_12|P|T|P _PG4_12|P|T|MID_SERIES 0  2e-13
R_PG4_12|P|T|B _PG4_12|P|T1 _PG4_12|P|T|MID_SHUNT  2.7439617672
L_PG4_12|P|T|RB _PG4_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|P|45|1 _PG4_12|P|T2 _PG4_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG4_12|P|45|B _PG4_12|P|T2 _PG4_12|P|45|MID_SHUNT  3.84154647408
L_PG4_12|P|45|RB _PG4_12|P|45|MID_SHUNT _PG4_12|P|A4  2.1704737578552e-12
B_PG4_12|P|6|1 _PG4_12|P|Q1 _PG4_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG4_12|P|6|P _PG4_12|P|6|MID_SERIES 0  2e-13
R_PG4_12|P|6|B _PG4_12|P|Q1 _PG4_12|P|6|MID_SHUNT  2.7439617672
L_PG4_12|P|6|RB _PG4_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_12|G|I_1|B _PG4_12|G|A1 _PG4_12|G|I_1|MID  2e-12
I_PG4_12|G|I_1|B 0 _PG4_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_12|G|I_3|B _PG4_12|G|A3 _PG4_12|G|I_3|MID  2e-12
I_PG4_12|G|I_3|B 0 _PG4_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_12|G|I_T|B _PG4_12|G|T1 _PG4_12|G|I_T|MID  2e-12
I_PG4_12|G|I_T|B 0 _PG4_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_12|G|I_6|B _PG4_12|G|Q1 _PG4_12|G|I_6|MID  2e-12
I_PG4_12|G|I_6|B 0 _PG4_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_12|G|1|1 _PG4_12|G|A1 _PG4_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG4_12|G|1|P _PG4_12|G|1|MID_SERIES 0  2e-13
R_PG4_12|G|1|B _PG4_12|G|A1 _PG4_12|G|1|MID_SHUNT  2.7439617672
L_PG4_12|G|1|RB _PG4_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|G|23|1 _PG4_12|G|A2 _PG4_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG4_12|G|23|B _PG4_12|G|A2 _PG4_12|G|23|MID_SHUNT  3.84154647408
L_PG4_12|G|23|RB _PG4_12|G|23|MID_SHUNT _PG4_12|G|A3  2.1704737578552e-12
B_PG4_12|G|3|1 _PG4_12|G|A3 _PG4_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG4_12|G|3|P _PG4_12|G|3|MID_SERIES 0  2e-13
R_PG4_12|G|3|B _PG4_12|G|A3 _PG4_12|G|3|MID_SHUNT  2.7439617672
L_PG4_12|G|3|RB _PG4_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|G|4|1 _PG4_12|G|A4 _PG4_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG4_12|G|4|P _PG4_12|G|4|MID_SERIES 0  2e-13
R_PG4_12|G|4|B _PG4_12|G|A4 _PG4_12|G|4|MID_SHUNT  2.7439617672
L_PG4_12|G|4|RB _PG4_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|G|T|1 _PG4_12|G|T1 _PG4_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG4_12|G|T|P _PG4_12|G|T|MID_SERIES 0  2e-13
R_PG4_12|G|T|B _PG4_12|G|T1 _PG4_12|G|T|MID_SHUNT  2.7439617672
L_PG4_12|G|T|RB _PG4_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_12|G|45|1 _PG4_12|G|T2 _PG4_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG4_12|G|45|B _PG4_12|G|T2 _PG4_12|G|45|MID_SHUNT  3.84154647408
L_PG4_12|G|45|RB _PG4_12|G|45|MID_SHUNT _PG4_12|G|A4  2.1704737578552e-12
B_PG4_12|G|6|1 _PG4_12|G|Q1 _PG4_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG4_12|G|6|P _PG4_12|G|6|MID_SERIES 0  2e-13
R_PG4_12|G|6|B _PG4_12|G|Q1 _PG4_12|G|6|MID_SHUNT  2.7439617672
L_PG4_12|G|6|RB _PG4_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_12|P|I_1|B _PG5_12|P|A1 _PG5_12|P|I_1|MID  2e-12
I_PG5_12|P|I_1|B 0 _PG5_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_12|P|I_3|B _PG5_12|P|A3 _PG5_12|P|I_3|MID  2e-12
I_PG5_12|P|I_3|B 0 _PG5_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_12|P|I_T|B _PG5_12|P|T1 _PG5_12|P|I_T|MID  2e-12
I_PG5_12|P|I_T|B 0 _PG5_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_12|P|I_6|B _PG5_12|P|Q1 _PG5_12|P|I_6|MID  2e-12
I_PG5_12|P|I_6|B 0 _PG5_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_12|P|1|1 _PG5_12|P|A1 _PG5_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG5_12|P|1|P _PG5_12|P|1|MID_SERIES 0  2e-13
R_PG5_12|P|1|B _PG5_12|P|A1 _PG5_12|P|1|MID_SHUNT  2.7439617672
L_PG5_12|P|1|RB _PG5_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|P|23|1 _PG5_12|P|A2 _PG5_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG5_12|P|23|B _PG5_12|P|A2 _PG5_12|P|23|MID_SHUNT  3.84154647408
L_PG5_12|P|23|RB _PG5_12|P|23|MID_SHUNT _PG5_12|P|A3  2.1704737578552e-12
B_PG5_12|P|3|1 _PG5_12|P|A3 _PG5_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG5_12|P|3|P _PG5_12|P|3|MID_SERIES 0  2e-13
R_PG5_12|P|3|B _PG5_12|P|A3 _PG5_12|P|3|MID_SHUNT  2.7439617672
L_PG5_12|P|3|RB _PG5_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|P|4|1 _PG5_12|P|A4 _PG5_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG5_12|P|4|P _PG5_12|P|4|MID_SERIES 0  2e-13
R_PG5_12|P|4|B _PG5_12|P|A4 _PG5_12|P|4|MID_SHUNT  2.7439617672
L_PG5_12|P|4|RB _PG5_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|P|T|1 _PG5_12|P|T1 _PG5_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG5_12|P|T|P _PG5_12|P|T|MID_SERIES 0  2e-13
R_PG5_12|P|T|B _PG5_12|P|T1 _PG5_12|P|T|MID_SHUNT  2.7439617672
L_PG5_12|P|T|RB _PG5_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|P|45|1 _PG5_12|P|T2 _PG5_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG5_12|P|45|B _PG5_12|P|T2 _PG5_12|P|45|MID_SHUNT  3.84154647408
L_PG5_12|P|45|RB _PG5_12|P|45|MID_SHUNT _PG5_12|P|A4  2.1704737578552e-12
B_PG5_12|P|6|1 _PG5_12|P|Q1 _PG5_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG5_12|P|6|P _PG5_12|P|6|MID_SERIES 0  2e-13
R_PG5_12|P|6|B _PG5_12|P|Q1 _PG5_12|P|6|MID_SHUNT  2.7439617672
L_PG5_12|P|6|RB _PG5_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_12|G|I_1|B _PG5_12|G|A1 _PG5_12|G|I_1|MID  2e-12
I_PG5_12|G|I_1|B 0 _PG5_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_12|G|I_3|B _PG5_12|G|A3 _PG5_12|G|I_3|MID  2e-12
I_PG5_12|G|I_3|B 0 _PG5_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_12|G|I_T|B _PG5_12|G|T1 _PG5_12|G|I_T|MID  2e-12
I_PG5_12|G|I_T|B 0 _PG5_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_12|G|I_6|B _PG5_12|G|Q1 _PG5_12|G|I_6|MID  2e-12
I_PG5_12|G|I_6|B 0 _PG5_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_12|G|1|1 _PG5_12|G|A1 _PG5_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG5_12|G|1|P _PG5_12|G|1|MID_SERIES 0  2e-13
R_PG5_12|G|1|B _PG5_12|G|A1 _PG5_12|G|1|MID_SHUNT  2.7439617672
L_PG5_12|G|1|RB _PG5_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|G|23|1 _PG5_12|G|A2 _PG5_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG5_12|G|23|B _PG5_12|G|A2 _PG5_12|G|23|MID_SHUNT  3.84154647408
L_PG5_12|G|23|RB _PG5_12|G|23|MID_SHUNT _PG5_12|G|A3  2.1704737578552e-12
B_PG5_12|G|3|1 _PG5_12|G|A3 _PG5_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG5_12|G|3|P _PG5_12|G|3|MID_SERIES 0  2e-13
R_PG5_12|G|3|B _PG5_12|G|A3 _PG5_12|G|3|MID_SHUNT  2.7439617672
L_PG5_12|G|3|RB _PG5_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|G|4|1 _PG5_12|G|A4 _PG5_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG5_12|G|4|P _PG5_12|G|4|MID_SERIES 0  2e-13
R_PG5_12|G|4|B _PG5_12|G|A4 _PG5_12|G|4|MID_SHUNT  2.7439617672
L_PG5_12|G|4|RB _PG5_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|G|T|1 _PG5_12|G|T1 _PG5_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG5_12|G|T|P _PG5_12|G|T|MID_SERIES 0  2e-13
R_PG5_12|G|T|B _PG5_12|G|T1 _PG5_12|G|T|MID_SHUNT  2.7439617672
L_PG5_12|G|T|RB _PG5_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_12|G|45|1 _PG5_12|G|T2 _PG5_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG5_12|G|45|B _PG5_12|G|T2 _PG5_12|G|45|MID_SHUNT  3.84154647408
L_PG5_12|G|45|RB _PG5_12|G|45|MID_SHUNT _PG5_12|G|A4  2.1704737578552e-12
B_PG5_12|G|6|1 _PG5_12|G|Q1 _PG5_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG5_12|G|6|P _PG5_12|G|6|MID_SERIES 0  2e-13
R_PG5_12|G|6|B _PG5_12|G|Q1 _PG5_12|G|6|MID_SHUNT  2.7439617672
L_PG5_12|G|6|RB _PG5_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_12|P|I_1|B _PG6_12|P|A1 _PG6_12|P|I_1|MID  2e-12
I_PG6_12|P|I_1|B 0 _PG6_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_12|P|I_3|B _PG6_12|P|A3 _PG6_12|P|I_3|MID  2e-12
I_PG6_12|P|I_3|B 0 _PG6_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_12|P|I_T|B _PG6_12|P|T1 _PG6_12|P|I_T|MID  2e-12
I_PG6_12|P|I_T|B 0 _PG6_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_12|P|I_6|B _PG6_12|P|Q1 _PG6_12|P|I_6|MID  2e-12
I_PG6_12|P|I_6|B 0 _PG6_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_12|P|1|1 _PG6_12|P|A1 _PG6_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG6_12|P|1|P _PG6_12|P|1|MID_SERIES 0  2e-13
R_PG6_12|P|1|B _PG6_12|P|A1 _PG6_12|P|1|MID_SHUNT  2.7439617672
L_PG6_12|P|1|RB _PG6_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|P|23|1 _PG6_12|P|A2 _PG6_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG6_12|P|23|B _PG6_12|P|A2 _PG6_12|P|23|MID_SHUNT  3.84154647408
L_PG6_12|P|23|RB _PG6_12|P|23|MID_SHUNT _PG6_12|P|A3  2.1704737578552e-12
B_PG6_12|P|3|1 _PG6_12|P|A3 _PG6_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG6_12|P|3|P _PG6_12|P|3|MID_SERIES 0  2e-13
R_PG6_12|P|3|B _PG6_12|P|A3 _PG6_12|P|3|MID_SHUNT  2.7439617672
L_PG6_12|P|3|RB _PG6_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|P|4|1 _PG6_12|P|A4 _PG6_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG6_12|P|4|P _PG6_12|P|4|MID_SERIES 0  2e-13
R_PG6_12|P|4|B _PG6_12|P|A4 _PG6_12|P|4|MID_SHUNT  2.7439617672
L_PG6_12|P|4|RB _PG6_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|P|T|1 _PG6_12|P|T1 _PG6_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG6_12|P|T|P _PG6_12|P|T|MID_SERIES 0  2e-13
R_PG6_12|P|T|B _PG6_12|P|T1 _PG6_12|P|T|MID_SHUNT  2.7439617672
L_PG6_12|P|T|RB _PG6_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|P|45|1 _PG6_12|P|T2 _PG6_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG6_12|P|45|B _PG6_12|P|T2 _PG6_12|P|45|MID_SHUNT  3.84154647408
L_PG6_12|P|45|RB _PG6_12|P|45|MID_SHUNT _PG6_12|P|A4  2.1704737578552e-12
B_PG6_12|P|6|1 _PG6_12|P|Q1 _PG6_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG6_12|P|6|P _PG6_12|P|6|MID_SERIES 0  2e-13
R_PG6_12|P|6|B _PG6_12|P|Q1 _PG6_12|P|6|MID_SHUNT  2.7439617672
L_PG6_12|P|6|RB _PG6_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_12|G|I_1|B _PG6_12|G|A1 _PG6_12|G|I_1|MID  2e-12
I_PG6_12|G|I_1|B 0 _PG6_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_12|G|I_3|B _PG6_12|G|A3 _PG6_12|G|I_3|MID  2e-12
I_PG6_12|G|I_3|B 0 _PG6_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_12|G|I_T|B _PG6_12|G|T1 _PG6_12|G|I_T|MID  2e-12
I_PG6_12|G|I_T|B 0 _PG6_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_12|G|I_6|B _PG6_12|G|Q1 _PG6_12|G|I_6|MID  2e-12
I_PG6_12|G|I_6|B 0 _PG6_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_12|G|1|1 _PG6_12|G|A1 _PG6_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG6_12|G|1|P _PG6_12|G|1|MID_SERIES 0  2e-13
R_PG6_12|G|1|B _PG6_12|G|A1 _PG6_12|G|1|MID_SHUNT  2.7439617672
L_PG6_12|G|1|RB _PG6_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|G|23|1 _PG6_12|G|A2 _PG6_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG6_12|G|23|B _PG6_12|G|A2 _PG6_12|G|23|MID_SHUNT  3.84154647408
L_PG6_12|G|23|RB _PG6_12|G|23|MID_SHUNT _PG6_12|G|A3  2.1704737578552e-12
B_PG6_12|G|3|1 _PG6_12|G|A3 _PG6_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG6_12|G|3|P _PG6_12|G|3|MID_SERIES 0  2e-13
R_PG6_12|G|3|B _PG6_12|G|A3 _PG6_12|G|3|MID_SHUNT  2.7439617672
L_PG6_12|G|3|RB _PG6_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|G|4|1 _PG6_12|G|A4 _PG6_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG6_12|G|4|P _PG6_12|G|4|MID_SERIES 0  2e-13
R_PG6_12|G|4|B _PG6_12|G|A4 _PG6_12|G|4|MID_SHUNT  2.7439617672
L_PG6_12|G|4|RB _PG6_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|G|T|1 _PG6_12|G|T1 _PG6_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG6_12|G|T|P _PG6_12|G|T|MID_SERIES 0  2e-13
R_PG6_12|G|T|B _PG6_12|G|T1 _PG6_12|G|T|MID_SHUNT  2.7439617672
L_PG6_12|G|T|RB _PG6_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_12|G|45|1 _PG6_12|G|T2 _PG6_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG6_12|G|45|B _PG6_12|G|T2 _PG6_12|G|45|MID_SHUNT  3.84154647408
L_PG6_12|G|45|RB _PG6_12|G|45|MID_SHUNT _PG6_12|G|A4  2.1704737578552e-12
B_PG6_12|G|6|1 _PG6_12|G|Q1 _PG6_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG6_12|G|6|P _PG6_12|G|6|MID_SERIES 0  2e-13
R_PG6_12|G|6|B _PG6_12|G|Q1 _PG6_12|G|6|MID_SHUNT  2.7439617672
L_PG6_12|G|6|RB _PG6_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_SPL_G1|I_D1|B _PG7_12|_SPL_G1|D1 _PG7_12|_SPL_G1|I_D1|MID  2e-12
I_PG7_12|_SPL_G1|I_D1|B 0 _PG7_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_12|_SPL_G1|I_D2|B _PG7_12|_SPL_G1|D2 _PG7_12|_SPL_G1|I_D2|MID  2e-12
I_PG7_12|_SPL_G1|I_D2|B 0 _PG7_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG7_12|_SPL_G1|I_Q1|B _PG7_12|_SPL_G1|QA1 _PG7_12|_SPL_G1|I_Q1|MID  2e-12
I_PG7_12|_SPL_G1|I_Q1|B 0 _PG7_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_12|_SPL_G1|I_Q2|B _PG7_12|_SPL_G1|QB1 _PG7_12|_SPL_G1|I_Q2|MID  2e-12
I_PG7_12|_SPL_G1|I_Q2|B 0 _PG7_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG7_12|_SPL_G1|1|1 _PG7_12|_SPL_G1|D1 _PG7_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_G1|1|P _PG7_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG7_12|_SPL_G1|1|B _PG7_12|_SPL_G1|D1 _PG7_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_G1|1|RB _PG7_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_SPL_G1|2|1 _PG7_12|_SPL_G1|D2 _PG7_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_G1|2|P _PG7_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG7_12|_SPL_G1|2|B _PG7_12|_SPL_G1|D2 _PG7_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_G1|2|RB _PG7_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_SPL_G1|A|1 _PG7_12|_SPL_G1|QA1 _PG7_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_G1|A|P _PG7_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG7_12|_SPL_G1|A|B _PG7_12|_SPL_G1|QA1 _PG7_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_G1|A|RB _PG7_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_SPL_G1|B|1 _PG7_12|_SPL_G1|QB1 _PG7_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_G1|B|P _PG7_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG7_12|_SPL_G1|B|B _PG7_12|_SPL_G1|QB1 _PG7_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_G1|B|RB _PG7_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_SPL_P1|I_D1|B _PG7_12|_SPL_P1|D1 _PG7_12|_SPL_P1|I_D1|MID  2e-12
I_PG7_12|_SPL_P1|I_D1|B 0 _PG7_12|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_12|_SPL_P1|I_D2|B _PG7_12|_SPL_P1|D2 _PG7_12|_SPL_P1|I_D2|MID  2e-12
I_PG7_12|_SPL_P1|I_D2|B 0 _PG7_12|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG7_12|_SPL_P1|I_Q1|B _PG7_12|_SPL_P1|QA1 _PG7_12|_SPL_P1|I_Q1|MID  2e-12
I_PG7_12|_SPL_P1|I_Q1|B 0 _PG7_12|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_12|_SPL_P1|I_Q2|B _PG7_12|_SPL_P1|QB1 _PG7_12|_SPL_P1|I_Q2|MID  2e-12
I_PG7_12|_SPL_P1|I_Q2|B 0 _PG7_12|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG7_12|_SPL_P1|1|1 _PG7_12|_SPL_P1|D1 _PG7_12|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_P1|1|P _PG7_12|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG7_12|_SPL_P1|1|B _PG7_12|_SPL_P1|D1 _PG7_12|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_P1|1|RB _PG7_12|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_SPL_P1|2|1 _PG7_12|_SPL_P1|D2 _PG7_12|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_P1|2|P _PG7_12|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG7_12|_SPL_P1|2|B _PG7_12|_SPL_P1|D2 _PG7_12|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_P1|2|RB _PG7_12|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_SPL_P1|A|1 _PG7_12|_SPL_P1|QA1 _PG7_12|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_P1|A|P _PG7_12|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG7_12|_SPL_P1|A|B _PG7_12|_SPL_P1|QA1 _PG7_12|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_P1|A|RB _PG7_12|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_SPL_P1|B|1 _PG7_12|_SPL_P1|QB1 _PG7_12|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_SPL_P1|B|P _PG7_12|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG7_12|_SPL_P1|B|B _PG7_12|_SPL_P1|QB1 _PG7_12|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG7_12|_SPL_P1|B|RB _PG7_12|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_PG|I_A1|B _PG7_12|_PG|A1 _PG7_12|_PG|I_A1|MID  2e-12
I_PG7_12|_PG|I_A1|B 0 _PG7_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_PG|I_B1|B _PG7_12|_PG|B1 _PG7_12|_PG|I_B1|MID  2e-12
I_PG7_12|_PG|I_B1|B 0 _PG7_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_PG|I_Q3|B _PG7_12|_PG|Q3 _PG7_12|_PG|I_Q3|MID  2e-12
I_PG7_12|_PG|I_Q3|B 0 _PG7_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_12|_PG|I_Q2|B _PG7_12|_PG|Q2 _PG7_12|_PG|I_Q2|MID  2e-12
I_PG7_12|_PG|I_Q2|B 0 _PG7_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_PG|I_Q1|B _PG7_12|_PG|Q1 _PG7_12|_PG|I_Q1|MID  2e-12
I_PG7_12|_PG|I_Q1|B 0 _PG7_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_PG|A1|1 _PG7_12|_PG|A1 _PG7_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_PG|A1|P _PG7_12|_PG|A1|MID_SERIES 0  2e-13
R_PG7_12|_PG|A1|B _PG7_12|_PG|A1 _PG7_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG7_12|_PG|A1|RB _PG7_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_PG|A2|1 _PG7_12|_PG|A2 _PG7_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_PG|A2|P _PG7_12|_PG|A2|MID_SERIES 0  2e-13
R_PG7_12|_PG|A2|B _PG7_12|_PG|A2 _PG7_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG7_12|_PG|A2|RB _PG7_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_PG|A12|1 _PG7_12|_PG|A2 _PG7_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_PG|A12|B _PG7_12|_PG|A2 _PG7_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG7_12|_PG|A12|RB _PG7_12|_PG|A12|MID_SHUNT _PG7_12|_PG|A3  2.1704737578552e-12
B_PG7_12|_PG|B1|1 _PG7_12|_PG|B1 _PG7_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_PG|B1|P _PG7_12|_PG|B1|MID_SERIES 0  2e-13
R_PG7_12|_PG|B1|B _PG7_12|_PG|B1 _PG7_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG7_12|_PG|B1|RB _PG7_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_PG|B2|1 _PG7_12|_PG|B2 _PG7_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_PG|B2|P _PG7_12|_PG|B2|MID_SERIES 0  2e-13
R_PG7_12|_PG|B2|B _PG7_12|_PG|B2 _PG7_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG7_12|_PG|B2|RB _PG7_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_PG|B12|1 _PG7_12|_PG|B2 _PG7_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG7_12|_PG|B12|B _PG7_12|_PG|B2 _PG7_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG7_12|_PG|B12|RB _PG7_12|_PG|B12|MID_SHUNT _PG7_12|_PG|B3  2.1704737578552e-12
B_PG7_12|_PG|Q2|1 _PG7_12|_PG|Q2 _PG7_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_PG|Q2|P _PG7_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG7_12|_PG|Q2|B _PG7_12|_PG|Q2 _PG7_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG7_12|_PG|Q2|RB _PG7_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_PG|Q1|1 _PG7_12|_PG|Q1 _PG7_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_PG|Q1|P _PG7_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG7_12|_PG|Q1|B _PG7_12|_PG|Q1 _PG7_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG7_12|_PG|Q1|RB _PG7_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_GG|I_A1|B _PG7_12|_GG|A1 _PG7_12|_GG|I_A1|MID  2e-12
I_PG7_12|_GG|I_A1|B 0 _PG7_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_GG|I_B1|B _PG7_12|_GG|B1 _PG7_12|_GG|I_B1|MID  2e-12
I_PG7_12|_GG|I_B1|B 0 _PG7_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_GG|I_Q3|B _PG7_12|_GG|Q3 _PG7_12|_GG|I_Q3|MID  2e-12
I_PG7_12|_GG|I_Q3|B 0 _PG7_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_12|_GG|I_Q2|B _PG7_12|_GG|Q2 _PG7_12|_GG|I_Q2|MID  2e-12
I_PG7_12|_GG|I_Q2|B 0 _PG7_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_GG|I_Q1|B _PG7_12|_GG|Q1 _PG7_12|_GG|I_Q1|MID  2e-12
I_PG7_12|_GG|I_Q1|B 0 _PG7_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_GG|A1|1 _PG7_12|_GG|A1 _PG7_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_GG|A1|P _PG7_12|_GG|A1|MID_SERIES 0  2e-13
R_PG7_12|_GG|A1|B _PG7_12|_GG|A1 _PG7_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG7_12|_GG|A1|RB _PG7_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_GG|A2|1 _PG7_12|_GG|A2 _PG7_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_GG|A2|P _PG7_12|_GG|A2|MID_SERIES 0  2e-13
R_PG7_12|_GG|A2|B _PG7_12|_GG|A2 _PG7_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG7_12|_GG|A2|RB _PG7_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_GG|A12|1 _PG7_12|_GG|A2 _PG7_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_GG|A12|B _PG7_12|_GG|A2 _PG7_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG7_12|_GG|A12|RB _PG7_12|_GG|A12|MID_SHUNT _PG7_12|_GG|A3  2.1704737578552e-12
B_PG7_12|_GG|B1|1 _PG7_12|_GG|B1 _PG7_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_GG|B1|P _PG7_12|_GG|B1|MID_SERIES 0  2e-13
R_PG7_12|_GG|B1|B _PG7_12|_GG|B1 _PG7_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG7_12|_GG|B1|RB _PG7_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_GG|B2|1 _PG7_12|_GG|B2 _PG7_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_GG|B2|P _PG7_12|_GG|B2|MID_SERIES 0  2e-13
R_PG7_12|_GG|B2|B _PG7_12|_GG|B2 _PG7_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG7_12|_GG|B2|RB _PG7_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_GG|B12|1 _PG7_12|_GG|B2 _PG7_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG7_12|_GG|B12|B _PG7_12|_GG|B2 _PG7_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG7_12|_GG|B12|RB _PG7_12|_GG|B12|MID_SHUNT _PG7_12|_GG|B3  2.1704737578552e-12
B_PG7_12|_GG|Q2|1 _PG7_12|_GG|Q2 _PG7_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_GG|Q2|P _PG7_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG7_12|_GG|Q2|B _PG7_12|_GG|Q2 _PG7_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG7_12|_GG|Q2|RB _PG7_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_GG|Q1|1 _PG7_12|_GG|Q1 _PG7_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_GG|Q1|P _PG7_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG7_12|_GG|Q1|B _PG7_12|_GG|Q1 _PG7_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG7_12|_GG|Q1|RB _PG7_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_DFF_P0|I_1|B _PG7_12|_DFF_P0|A1 _PG7_12|_DFF_P0|I_1|MID  2e-12
I_PG7_12|_DFF_P0|I_1|B 0 _PG7_12|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_P0|I_3|B _PG7_12|_DFF_P0|A3 _PG7_12|_DFF_P0|I_3|MID  2e-12
I_PG7_12|_DFF_P0|I_3|B 0 _PG7_12|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_12|_DFF_P0|I_T|B _PG7_12|_DFF_P0|T1 _PG7_12|_DFF_P0|I_T|MID  2e-12
I_PG7_12|_DFF_P0|I_T|B 0 _PG7_12|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_P0|I_6|B _PG7_12|_DFF_P0|Q1 _PG7_12|_DFF_P0|I_6|MID  2e-12
I_PG7_12|_DFF_P0|I_6|B 0 _PG7_12|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_DFF_P0|1|1 _PG7_12|_DFF_P0|A1 _PG7_12|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P0|1|P _PG7_12|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P0|1|B _PG7_12|_DFF_P0|A1 _PG7_12|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P0|1|RB _PG7_12|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P0|23|1 _PG7_12|_DFF_P0|A2 _PG7_12|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_P0|23|B _PG7_12|_DFF_P0|A2 _PG7_12|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_P0|23|RB _PG7_12|_DFF_P0|23|MID_SHUNT _PG7_12|_DFF_P0|A3  2.1704737578552e-12
B_PG7_12|_DFF_P0|3|1 _PG7_12|_DFF_P0|A3 _PG7_12|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P0|3|P _PG7_12|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P0|3|B _PG7_12|_DFF_P0|A3 _PG7_12|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P0|3|RB _PG7_12|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P0|4|1 _PG7_12|_DFF_P0|A4 _PG7_12|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P0|4|P _PG7_12|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P0|4|B _PG7_12|_DFF_P0|A4 _PG7_12|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P0|4|RB _PG7_12|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P0|T|1 _PG7_12|_DFF_P0|T1 _PG7_12|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P0|T|P _PG7_12|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P0|T|B _PG7_12|_DFF_P0|T1 _PG7_12|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P0|T|RB _PG7_12|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P0|45|1 _PG7_12|_DFF_P0|T2 _PG7_12|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_P0|45|B _PG7_12|_DFF_P0|T2 _PG7_12|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_P0|45|RB _PG7_12|_DFF_P0|45|MID_SHUNT _PG7_12|_DFF_P0|A4  2.1704737578552e-12
B_PG7_12|_DFF_P0|6|1 _PG7_12|_DFF_P0|Q1 _PG7_12|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P0|6|P _PG7_12|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P0|6|B _PG7_12|_DFF_P0|Q1 _PG7_12|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P0|6|RB _PG7_12|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_DFF_P1|I_1|B _PG7_12|_DFF_P1|A1 _PG7_12|_DFF_P1|I_1|MID  2e-12
I_PG7_12|_DFF_P1|I_1|B 0 _PG7_12|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_P1|I_3|B _PG7_12|_DFF_P1|A3 _PG7_12|_DFF_P1|I_3|MID  2e-12
I_PG7_12|_DFF_P1|I_3|B 0 _PG7_12|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_12|_DFF_P1|I_T|B _PG7_12|_DFF_P1|T1 _PG7_12|_DFF_P1|I_T|MID  2e-12
I_PG7_12|_DFF_P1|I_T|B 0 _PG7_12|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_P1|I_6|B _PG7_12|_DFF_P1|Q1 _PG7_12|_DFF_P1|I_6|MID  2e-12
I_PG7_12|_DFF_P1|I_6|B 0 _PG7_12|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_DFF_P1|1|1 _PG7_12|_DFF_P1|A1 _PG7_12|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P1|1|P _PG7_12|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P1|1|B _PG7_12|_DFF_P1|A1 _PG7_12|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P1|1|RB _PG7_12|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P1|23|1 _PG7_12|_DFF_P1|A2 _PG7_12|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_P1|23|B _PG7_12|_DFF_P1|A2 _PG7_12|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_P1|23|RB _PG7_12|_DFF_P1|23|MID_SHUNT _PG7_12|_DFF_P1|A3  2.1704737578552e-12
B_PG7_12|_DFF_P1|3|1 _PG7_12|_DFF_P1|A3 _PG7_12|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P1|3|P _PG7_12|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P1|3|B _PG7_12|_DFF_P1|A3 _PG7_12|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P1|3|RB _PG7_12|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P1|4|1 _PG7_12|_DFF_P1|A4 _PG7_12|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P1|4|P _PG7_12|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P1|4|B _PG7_12|_DFF_P1|A4 _PG7_12|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P1|4|RB _PG7_12|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P1|T|1 _PG7_12|_DFF_P1|T1 _PG7_12|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P1|T|P _PG7_12|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P1|T|B _PG7_12|_DFF_P1|T1 _PG7_12|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P1|T|RB _PG7_12|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_P1|45|1 _PG7_12|_DFF_P1|T2 _PG7_12|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_P1|45|B _PG7_12|_DFF_P1|T2 _PG7_12|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_P1|45|RB _PG7_12|_DFF_P1|45|MID_SHUNT _PG7_12|_DFF_P1|A4  2.1704737578552e-12
B_PG7_12|_DFF_P1|6|1 _PG7_12|_DFF_P1|Q1 _PG7_12|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_P1|6|P _PG7_12|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG7_12|_DFF_P1|6|B _PG7_12|_DFF_P1|Q1 _PG7_12|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_P1|6|RB _PG7_12|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_DFF_PG|I_1|B _PG7_12|_DFF_PG|A1 _PG7_12|_DFF_PG|I_1|MID  2e-12
I_PG7_12|_DFF_PG|I_1|B 0 _PG7_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_PG|I_3|B _PG7_12|_DFF_PG|A3 _PG7_12|_DFF_PG|I_3|MID  2e-12
I_PG7_12|_DFF_PG|I_3|B 0 _PG7_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_12|_DFF_PG|I_T|B _PG7_12|_DFF_PG|T1 _PG7_12|_DFF_PG|I_T|MID  2e-12
I_PG7_12|_DFF_PG|I_T|B 0 _PG7_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_PG|I_6|B _PG7_12|_DFF_PG|Q1 _PG7_12|_DFF_PG|I_6|MID  2e-12
I_PG7_12|_DFF_PG|I_6|B 0 _PG7_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_DFF_PG|1|1 _PG7_12|_DFF_PG|A1 _PG7_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_PG|1|P _PG7_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG7_12|_DFF_PG|1|B _PG7_12|_DFF_PG|A1 _PG7_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_PG|1|RB _PG7_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_PG|23|1 _PG7_12|_DFF_PG|A2 _PG7_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_PG|23|B _PG7_12|_DFF_PG|A2 _PG7_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_PG|23|RB _PG7_12|_DFF_PG|23|MID_SHUNT _PG7_12|_DFF_PG|A3  2.1704737578552e-12
B_PG7_12|_DFF_PG|3|1 _PG7_12|_DFF_PG|A3 _PG7_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_PG|3|P _PG7_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG7_12|_DFF_PG|3|B _PG7_12|_DFF_PG|A3 _PG7_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_PG|3|RB _PG7_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_PG|4|1 _PG7_12|_DFF_PG|A4 _PG7_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_PG|4|P _PG7_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG7_12|_DFF_PG|4|B _PG7_12|_DFF_PG|A4 _PG7_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_PG|4|RB _PG7_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_PG|T|1 _PG7_12|_DFF_PG|T1 _PG7_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_PG|T|P _PG7_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG7_12|_DFF_PG|T|B _PG7_12|_DFF_PG|T1 _PG7_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_PG|T|RB _PG7_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_PG|45|1 _PG7_12|_DFF_PG|T2 _PG7_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_PG|45|B _PG7_12|_DFF_PG|T2 _PG7_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_PG|45|RB _PG7_12|_DFF_PG|45|MID_SHUNT _PG7_12|_DFF_PG|A4  2.1704737578552e-12
B_PG7_12|_DFF_PG|6|1 _PG7_12|_DFF_PG|Q1 _PG7_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_PG|6|P _PG7_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG7_12|_DFF_PG|6|B _PG7_12|_DFF_PG|Q1 _PG7_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_PG|6|RB _PG7_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_DFF_GG|I_1|B _PG7_12|_DFF_GG|A1 _PG7_12|_DFF_GG|I_1|MID  2e-12
I_PG7_12|_DFF_GG|I_1|B 0 _PG7_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_GG|I_3|B _PG7_12|_DFF_GG|A3 _PG7_12|_DFF_GG|I_3|MID  2e-12
I_PG7_12|_DFF_GG|I_3|B 0 _PG7_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_12|_DFF_GG|I_T|B _PG7_12|_DFF_GG|T1 _PG7_12|_DFF_GG|I_T|MID  2e-12
I_PG7_12|_DFF_GG|I_T|B 0 _PG7_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_DFF_GG|I_6|B _PG7_12|_DFF_GG|Q1 _PG7_12|_DFF_GG|I_6|MID  2e-12
I_PG7_12|_DFF_GG|I_6|B 0 _PG7_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_DFF_GG|1|1 _PG7_12|_DFF_GG|A1 _PG7_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_GG|1|P _PG7_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG7_12|_DFF_GG|1|B _PG7_12|_DFF_GG|A1 _PG7_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_GG|1|RB _PG7_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_GG|23|1 _PG7_12|_DFF_GG|A2 _PG7_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_GG|23|B _PG7_12|_DFF_GG|A2 _PG7_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_GG|23|RB _PG7_12|_DFF_GG|23|MID_SHUNT _PG7_12|_DFF_GG|A3  2.1704737578552e-12
B_PG7_12|_DFF_GG|3|1 _PG7_12|_DFF_GG|A3 _PG7_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_GG|3|P _PG7_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG7_12|_DFF_GG|3|B _PG7_12|_DFF_GG|A3 _PG7_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_GG|3|RB _PG7_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_GG|4|1 _PG7_12|_DFF_GG|A4 _PG7_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_GG|4|P _PG7_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG7_12|_DFF_GG|4|B _PG7_12|_DFF_GG|A4 _PG7_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_GG|4|RB _PG7_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_GG|T|1 _PG7_12|_DFF_GG|T1 _PG7_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_GG|T|P _PG7_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG7_12|_DFF_GG|T|B _PG7_12|_DFF_GG|T1 _PG7_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_GG|T|RB _PG7_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_DFF_GG|45|1 _PG7_12|_DFF_GG|T2 _PG7_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG7_12|_DFF_GG|45|B _PG7_12|_DFF_GG|T2 _PG7_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG7_12|_DFF_GG|45|RB _PG7_12|_DFF_GG|45|MID_SHUNT _PG7_12|_DFF_GG|A4  2.1704737578552e-12
B_PG7_12|_DFF_GG|6|1 _PG7_12|_DFF_GG|Q1 _PG7_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_DFF_GG|6|P _PG7_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG7_12|_DFF_GG|6|B _PG7_12|_DFF_GG|Q1 _PG7_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG7_12|_DFF_GG|6|RB _PG7_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_AND_G|I_A1|B _PG7_12|_AND_G|A1 _PG7_12|_AND_G|I_A1|MID  2e-12
I_PG7_12|_AND_G|I_A1|B 0 _PG7_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_AND_G|I_B1|B _PG7_12|_AND_G|B1 _PG7_12|_AND_G|I_B1|MID  2e-12
I_PG7_12|_AND_G|I_B1|B 0 _PG7_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_AND_G|I_Q3|B _PG7_12|_AND_G|Q3 _PG7_12|_AND_G|I_Q3|MID  2e-12
I_PG7_12|_AND_G|I_Q3|B 0 _PG7_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG7_12|_AND_G|I_Q2|B _PG7_12|_AND_G|Q2 _PG7_12|_AND_G|I_Q2|MID  2e-12
I_PG7_12|_AND_G|I_Q2|B 0 _PG7_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_AND_G|I_Q1|B _PG7_12|_AND_G|Q1 _PG7_12|_AND_G|I_Q1|MID  2e-12
I_PG7_12|_AND_G|I_Q1|B 0 _PG7_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_AND_G|A1|1 _PG7_12|_AND_G|A1 _PG7_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_G|A1|P _PG7_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG7_12|_AND_G|A1|B _PG7_12|_AND_G|A1 _PG7_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG7_12|_AND_G|A1|RB _PG7_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_G|A2|1 _PG7_12|_AND_G|A2 _PG7_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_G|A2|P _PG7_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG7_12|_AND_G|A2|B _PG7_12|_AND_G|A2 _PG7_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG7_12|_AND_G|A2|RB _PG7_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_G|A12|1 _PG7_12|_AND_G|A2 _PG7_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_AND_G|A12|B _PG7_12|_AND_G|A2 _PG7_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG7_12|_AND_G|A12|RB _PG7_12|_AND_G|A12|MID_SHUNT _PG7_12|_AND_G|A3  2.1704737578552e-12
B_PG7_12|_AND_G|B1|1 _PG7_12|_AND_G|B1 _PG7_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_G|B1|P _PG7_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG7_12|_AND_G|B1|B _PG7_12|_AND_G|B1 _PG7_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG7_12|_AND_G|B1|RB _PG7_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_G|B2|1 _PG7_12|_AND_G|B2 _PG7_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_G|B2|P _PG7_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG7_12|_AND_G|B2|B _PG7_12|_AND_G|B2 _PG7_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG7_12|_AND_G|B2|RB _PG7_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_G|B12|1 _PG7_12|_AND_G|B2 _PG7_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG7_12|_AND_G|B12|B _PG7_12|_AND_G|B2 _PG7_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG7_12|_AND_G|B12|RB _PG7_12|_AND_G|B12|MID_SHUNT _PG7_12|_AND_G|B3  2.1704737578552e-12
B_PG7_12|_AND_G|Q2|1 _PG7_12|_AND_G|Q2 _PG7_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_G|Q2|P _PG7_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG7_12|_AND_G|Q2|B _PG7_12|_AND_G|Q2 _PG7_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG7_12|_AND_G|Q2|RB _PG7_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_G|Q1|1 _PG7_12|_AND_G|Q1 _PG7_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_G|Q1|P _PG7_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG7_12|_AND_G|Q1|B _PG7_12|_AND_G|Q1 _PG7_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG7_12|_AND_G|Q1|RB _PG7_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_12|_AND_P|I_A1|B _PG7_12|_AND_P|A1 _PG7_12|_AND_P|I_A1|MID  2e-12
I_PG7_12|_AND_P|I_A1|B 0 _PG7_12|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_AND_P|I_B1|B _PG7_12|_AND_P|B1 _PG7_12|_AND_P|I_B1|MID  2e-12
I_PG7_12|_AND_P|I_B1|B 0 _PG7_12|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_AND_P|I_Q3|B _PG7_12|_AND_P|Q3 _PG7_12|_AND_P|I_Q3|MID  2e-12
I_PG7_12|_AND_P|I_Q3|B 0 _PG7_12|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG7_12|_AND_P|I_Q2|B _PG7_12|_AND_P|Q2 _PG7_12|_AND_P|I_Q2|MID  2e-12
I_PG7_12|_AND_P|I_Q2|B 0 _PG7_12|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_12|_AND_P|I_Q1|B _PG7_12|_AND_P|Q1 _PG7_12|_AND_P|I_Q1|MID  2e-12
I_PG7_12|_AND_P|I_Q1|B 0 _PG7_12|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_12|_AND_P|A1|1 _PG7_12|_AND_P|A1 _PG7_12|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_P|A1|P _PG7_12|_AND_P|A1|MID_SERIES 0  2e-13
R_PG7_12|_AND_P|A1|B _PG7_12|_AND_P|A1 _PG7_12|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG7_12|_AND_P|A1|RB _PG7_12|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_P|A2|1 _PG7_12|_AND_P|A2 _PG7_12|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_P|A2|P _PG7_12|_AND_P|A2|MID_SERIES 0  2e-13
R_PG7_12|_AND_P|A2|B _PG7_12|_AND_P|A2 _PG7_12|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG7_12|_AND_P|A2|RB _PG7_12|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_P|A12|1 _PG7_12|_AND_P|A2 _PG7_12|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG7_12|_AND_P|A12|B _PG7_12|_AND_P|A2 _PG7_12|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG7_12|_AND_P|A12|RB _PG7_12|_AND_P|A12|MID_SHUNT _PG7_12|_AND_P|A3  2.1704737578552e-12
B_PG7_12|_AND_P|B1|1 _PG7_12|_AND_P|B1 _PG7_12|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_P|B1|P _PG7_12|_AND_P|B1|MID_SERIES 0  2e-13
R_PG7_12|_AND_P|B1|B _PG7_12|_AND_P|B1 _PG7_12|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG7_12|_AND_P|B1|RB _PG7_12|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_P|B2|1 _PG7_12|_AND_P|B2 _PG7_12|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_P|B2|P _PG7_12|_AND_P|B2|MID_SERIES 0  2e-13
R_PG7_12|_AND_P|B2|B _PG7_12|_AND_P|B2 _PG7_12|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG7_12|_AND_P|B2|RB _PG7_12|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_P|B12|1 _PG7_12|_AND_P|B2 _PG7_12|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG7_12|_AND_P|B12|B _PG7_12|_AND_P|B2 _PG7_12|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG7_12|_AND_P|B12|RB _PG7_12|_AND_P|B12|MID_SHUNT _PG7_12|_AND_P|B3  2.1704737578552e-12
B_PG7_12|_AND_P|Q2|1 _PG7_12|_AND_P|Q2 _PG7_12|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_P|Q2|P _PG7_12|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG7_12|_AND_P|Q2|B _PG7_12|_AND_P|Q2 _PG7_12|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG7_12|_AND_P|Q2|RB _PG7_12|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_12|_AND_P|Q1|1 _PG7_12|_AND_P|Q1 _PG7_12|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_12|_AND_P|Q1|P _PG7_12|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG7_12|_AND_P|Q1|B _PG7_12|_AND_P|Q1 _PG7_12|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG7_12|_AND_P|Q1|RB _PG7_12|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PTL_P3_2|_SPL|SPL1|1 _PTL_P3_2|D _PTL_P3_2|_SPL|SPL1|D1  2e-12
L_PTL_P3_2|_SPL|SPL1|2 _PTL_P3_2|_SPL|SPL1|D1 _PTL_P3_2|_SPL|SPL1|D2  4.135667696e-12
L_PTL_P3_2|_SPL|SPL1|3 _PTL_P3_2|_SPL|SPL1|D2 _PTL_P3_2|_SPL|SPL1|JCT  9.84682784761905e-13
L_PTL_P3_2|_SPL|SPL1|4 _PTL_P3_2|_SPL|SPL1|JCT _PTL_P3_2|_SPL|SPL1|QA1  9.84682784761905e-13
L_PTL_P3_2|_SPL|SPL1|5 _PTL_P3_2|_SPL|SPL1|QA1 P3_2_TO4  2e-12
L_PTL_P3_2|_SPL|SPL1|6 _PTL_P3_2|_SPL|SPL1|JCT _PTL_P3_2|_SPL|SPL1|QB1  9.84682784761905e-13
L_PTL_P3_2|_SPL|SPL1|7 _PTL_P3_2|_SPL|SPL1|QB1 _PTL_P3_2|_SPL|QTMP  2e-12
L_PTL_P3_2|_SPL|SPL2|1 _PTL_P3_2|_SPL|QTMP _PTL_P3_2|_SPL|SPL2|D1  2e-12
L_PTL_P3_2|_SPL|SPL2|2 _PTL_P3_2|_SPL|SPL2|D1 _PTL_P3_2|_SPL|SPL2|D2  4.135667696e-12
L_PTL_P3_2|_SPL|SPL2|3 _PTL_P3_2|_SPL|SPL2|D2 _PTL_P3_2|_SPL|SPL2|JCT  9.84682784761905e-13
L_PTL_P3_2|_SPL|SPL2|4 _PTL_P3_2|_SPL|SPL2|JCT _PTL_P3_2|_SPL|SPL2|QA1  9.84682784761905e-13
L_PTL_P3_2|_SPL|SPL2|5 _PTL_P3_2|_SPL|SPL2|QA1 P3_2_TO5  2e-12
L_PTL_P3_2|_SPL|SPL2|6 _PTL_P3_2|_SPL|SPL2|JCT _PTL_P3_2|_SPL|SPL2|QB1  9.84682784761905e-13
L_PTL_P3_2|_SPL|SPL2|7 _PTL_P3_2|_SPL|SPL2|QB1 P3_2_TO7  2e-12
L_PTL_G3_2|_SPL_1|I_D1|B _PTL_G3_2|_SPL_1|D1 _PTL_G3_2|_SPL_1|I_D1|MID  2e-12
I_PTL_G3_2|_SPL_1|I_D1|B 0 _PTL_G3_2|_SPL_1|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_SPL_1|I_D2|B _PTL_G3_2|_SPL_1|D2 _PTL_G3_2|_SPL_1|I_D2|MID  2e-12
I_PTL_G3_2|_SPL_1|I_D2|B 0 _PTL_G3_2|_SPL_1|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G3_2|_SPL_1|I_Q1|B _PTL_G3_2|_SPL_1|QA1 _PTL_G3_2|_SPL_1|I_Q1|MID  2e-12
I_PTL_G3_2|_SPL_1|I_Q1|B 0 _PTL_G3_2|_SPL_1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_SPL_1|I_Q2|B _PTL_G3_2|_SPL_1|QB1 _PTL_G3_2|_SPL_1|I_Q2|MID  2e-12
I_PTL_G3_2|_SPL_1|I_Q2|B 0 _PTL_G3_2|_SPL_1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G3_2|_SPL_1|1|1 _PTL_G3_2|_SPL_1|D1 _PTL_G3_2|_SPL_1|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_1|1|P _PTL_G3_2|_SPL_1|1|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_1|1|B _PTL_G3_2|_SPL_1|D1 _PTL_G3_2|_SPL_1|1|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_1|1|RB _PTL_G3_2|_SPL_1|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_1|2|1 _PTL_G3_2|_SPL_1|D2 _PTL_G3_2|_SPL_1|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_1|2|P _PTL_G3_2|_SPL_1|2|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_1|2|B _PTL_G3_2|_SPL_1|D2 _PTL_G3_2|_SPL_1|2|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_1|2|RB _PTL_G3_2|_SPL_1|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_1|A|1 _PTL_G3_2|_SPL_1|QA1 _PTL_G3_2|_SPL_1|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_1|A|P _PTL_G3_2|_SPL_1|A|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_1|A|B _PTL_G3_2|_SPL_1|QA1 _PTL_G3_2|_SPL_1|A|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_1|A|RB _PTL_G3_2|_SPL_1|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_1|B|1 _PTL_G3_2|_SPL_1|QB1 _PTL_G3_2|_SPL_1|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_1|B|P _PTL_G3_2|_SPL_1|B|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_1|B|B _PTL_G3_2|_SPL_1|QB1 _PTL_G3_2|_SPL_1|B|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_1|B|RB _PTL_G3_2|_SPL_1|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_G3_2|_SPL_2|I_D1|B _PTL_G3_2|_SPL_2|D1 _PTL_G3_2|_SPL_2|I_D1|MID  2e-12
I_PTL_G3_2|_SPL_2|I_D1|B 0 _PTL_G3_2|_SPL_2|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_SPL_2|I_D2|B _PTL_G3_2|_SPL_2|D2 _PTL_G3_2|_SPL_2|I_D2|MID  2e-12
I_PTL_G3_2|_SPL_2|I_D2|B 0 _PTL_G3_2|_SPL_2|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G3_2|_SPL_2|I_Q1|B _PTL_G3_2|_SPL_2|QA1 _PTL_G3_2|_SPL_2|I_Q1|MID  2e-12
I_PTL_G3_2|_SPL_2|I_Q1|B 0 _PTL_G3_2|_SPL_2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_SPL_2|I_Q2|B _PTL_G3_2|_SPL_2|QB1 _PTL_G3_2|_SPL_2|I_Q2|MID  2e-12
I_PTL_G3_2|_SPL_2|I_Q2|B 0 _PTL_G3_2|_SPL_2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G3_2|_SPL_2|1|1 _PTL_G3_2|_SPL_2|D1 _PTL_G3_2|_SPL_2|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_2|1|P _PTL_G3_2|_SPL_2|1|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_2|1|B _PTL_G3_2|_SPL_2|D1 _PTL_G3_2|_SPL_2|1|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_2|1|RB _PTL_G3_2|_SPL_2|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_2|2|1 _PTL_G3_2|_SPL_2|D2 _PTL_G3_2|_SPL_2|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_2|2|P _PTL_G3_2|_SPL_2|2|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_2|2|B _PTL_G3_2|_SPL_2|D2 _PTL_G3_2|_SPL_2|2|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_2|2|RB _PTL_G3_2|_SPL_2|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_2|A|1 _PTL_G3_2|_SPL_2|QA1 _PTL_G3_2|_SPL_2|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_2|A|P _PTL_G3_2|_SPL_2|A|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_2|A|B _PTL_G3_2|_SPL_2|QA1 _PTL_G3_2|_SPL_2|A|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_2|A|RB _PTL_G3_2|_SPL_2|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_2|B|1 _PTL_G3_2|_SPL_2|QB1 _PTL_G3_2|_SPL_2|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_2|B|P _PTL_G3_2|_SPL_2|B|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_2|B|B _PTL_G3_2|_SPL_2|QB1 _PTL_G3_2|_SPL_2|B|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_2|B|RB _PTL_G3_2|_SPL_2|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_G3_2|_SPL_3|I_D1|B _PTL_G3_2|_SPL_3|D1 _PTL_G3_2|_SPL_3|I_D1|MID  2e-12
I_PTL_G3_2|_SPL_3|I_D1|B 0 _PTL_G3_2|_SPL_3|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_SPL_3|I_D2|B _PTL_G3_2|_SPL_3|D2 _PTL_G3_2|_SPL_3|I_D2|MID  2e-12
I_PTL_G3_2|_SPL_3|I_D2|B 0 _PTL_G3_2|_SPL_3|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G3_2|_SPL_3|I_Q1|B _PTL_G3_2|_SPL_3|QA1 _PTL_G3_2|_SPL_3|I_Q1|MID  2e-12
I_PTL_G3_2|_SPL_3|I_Q1|B 0 _PTL_G3_2|_SPL_3|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G3_2|_SPL_3|I_Q2|B _PTL_G3_2|_SPL_3|QB1 _PTL_G3_2|_SPL_3|I_Q2|MID  2e-12
I_PTL_G3_2|_SPL_3|I_Q2|B 0 _PTL_G3_2|_SPL_3|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G3_2|_SPL_3|1|1 _PTL_G3_2|_SPL_3|D1 _PTL_G3_2|_SPL_3|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_3|1|P _PTL_G3_2|_SPL_3|1|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_3|1|B _PTL_G3_2|_SPL_3|D1 _PTL_G3_2|_SPL_3|1|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_3|1|RB _PTL_G3_2|_SPL_3|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_3|2|1 _PTL_G3_2|_SPL_3|D2 _PTL_G3_2|_SPL_3|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_3|2|P _PTL_G3_2|_SPL_3|2|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_3|2|B _PTL_G3_2|_SPL_3|D2 _PTL_G3_2|_SPL_3|2|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_3|2|RB _PTL_G3_2|_SPL_3|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_3|A|1 _PTL_G3_2|_SPL_3|QA1 _PTL_G3_2|_SPL_3|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_3|A|P _PTL_G3_2|_SPL_3|A|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_3|A|B _PTL_G3_2|_SPL_3|QA1 _PTL_G3_2|_SPL_3|A|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_3|A|RB _PTL_G3_2|_SPL_3|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G3_2|_SPL_3|B|1 _PTL_G3_2|_SPL_3|QB1 _PTL_G3_2|_SPL_3|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G3_2|_SPL_3|B|P _PTL_G3_2|_SPL_3|B|MID_SERIES 0  2e-13
R_PTL_G3_2|_SPL_3|B|B _PTL_G3_2|_SPL_3|QB1 _PTL_G3_2|_SPL_3|B|MID_SHUNT  2.7439617672
L_PTL_G3_2|_SPL_3|B|RB _PTL_G3_2|_SPL_3|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_P4_2|_SPL|I_D1|B _PTL_P4_2|_SPL|D1 _PTL_P4_2|_SPL|I_D1|MID  2e-12
I_PTL_P4_2|_SPL|I_D1|B 0 _PTL_P4_2|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P4_2|_SPL|I_D2|B _PTL_P4_2|_SPL|D2 _PTL_P4_2|_SPL|I_D2|MID  2e-12
I_PTL_P4_2|_SPL|I_D2|B 0 _PTL_P4_2|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P4_2|_SPL|I_Q1|B _PTL_P4_2|_SPL|QA1 _PTL_P4_2|_SPL|I_Q1|MID  2e-12
I_PTL_P4_2|_SPL|I_Q1|B 0 _PTL_P4_2|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P4_2|_SPL|I_Q2|B _PTL_P4_2|_SPL|QB1 _PTL_P4_2|_SPL|I_Q2|MID  2e-12
I_PTL_P4_2|_SPL|I_Q2|B 0 _PTL_P4_2|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P4_2|_SPL|1|1 _PTL_P4_2|_SPL|D1 _PTL_P4_2|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P4_2|_SPL|1|P _PTL_P4_2|_SPL|1|MID_SERIES 0  2e-13
R_PTL_P4_2|_SPL|1|B _PTL_P4_2|_SPL|D1 _PTL_P4_2|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_P4_2|_SPL|1|RB _PTL_P4_2|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P4_2|_SPL|2|1 _PTL_P4_2|_SPL|D2 _PTL_P4_2|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P4_2|_SPL|2|P _PTL_P4_2|_SPL|2|MID_SERIES 0  2e-13
R_PTL_P4_2|_SPL|2|B _PTL_P4_2|_SPL|D2 _PTL_P4_2|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_P4_2|_SPL|2|RB _PTL_P4_2|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P4_2|_SPL|A|1 _PTL_P4_2|_SPL|QA1 _PTL_P4_2|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P4_2|_SPL|A|P _PTL_P4_2|_SPL|A|MID_SERIES 0  2e-13
R_PTL_P4_2|_SPL|A|B _PTL_P4_2|_SPL|QA1 _PTL_P4_2|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_P4_2|_SPL|A|RB _PTL_P4_2|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P4_2|_SPL|B|1 _PTL_P4_2|_SPL|QB1 _PTL_P4_2|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P4_2|_SPL|B|P _PTL_P4_2|_SPL|B|MID_SERIES 0  2e-13
R_PTL_P4_2|_SPL|B|B _PTL_P4_2|_SPL|QB1 _PTL_P4_2|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_P4_2|_SPL|B|RB _PTL_P4_2|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_SPL_G1|I_D1|B _PG4_23|_SPL_G1|D1 _PG4_23|_SPL_G1|I_D1|MID  2e-12
I_PG4_23|_SPL_G1|I_D1|B 0 _PG4_23|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG4_23|_SPL_G1|I_D2|B _PG4_23|_SPL_G1|D2 _PG4_23|_SPL_G1|I_D2|MID  2e-12
I_PG4_23|_SPL_G1|I_D2|B 0 _PG4_23|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG4_23|_SPL_G1|I_Q1|B _PG4_23|_SPL_G1|QA1 _PG4_23|_SPL_G1|I_Q1|MID  2e-12
I_PG4_23|_SPL_G1|I_Q1|B 0 _PG4_23|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG4_23|_SPL_G1|I_Q2|B _PG4_23|_SPL_G1|QB1 _PG4_23|_SPL_G1|I_Q2|MID  2e-12
I_PG4_23|_SPL_G1|I_Q2|B 0 _PG4_23|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG4_23|_SPL_G1|1|1 _PG4_23|_SPL_G1|D1 _PG4_23|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_G1|1|P _PG4_23|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG4_23|_SPL_G1|1|B _PG4_23|_SPL_G1|D1 _PG4_23|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_G1|1|RB _PG4_23|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_SPL_G1|2|1 _PG4_23|_SPL_G1|D2 _PG4_23|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_G1|2|P _PG4_23|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG4_23|_SPL_G1|2|B _PG4_23|_SPL_G1|D2 _PG4_23|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_G1|2|RB _PG4_23|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_SPL_G1|A|1 _PG4_23|_SPL_G1|QA1 _PG4_23|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_G1|A|P _PG4_23|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG4_23|_SPL_G1|A|B _PG4_23|_SPL_G1|QA1 _PG4_23|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_G1|A|RB _PG4_23|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_SPL_G1|B|1 _PG4_23|_SPL_G1|QB1 _PG4_23|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_G1|B|P _PG4_23|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG4_23|_SPL_G1|B|B _PG4_23|_SPL_G1|QB1 _PG4_23|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_G1|B|RB _PG4_23|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_SPL_P1|I_D1|B _PG4_23|_SPL_P1|D1 _PG4_23|_SPL_P1|I_D1|MID  2e-12
I_PG4_23|_SPL_P1|I_D1|B 0 _PG4_23|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG4_23|_SPL_P1|I_D2|B _PG4_23|_SPL_P1|D2 _PG4_23|_SPL_P1|I_D2|MID  2e-12
I_PG4_23|_SPL_P1|I_D2|B 0 _PG4_23|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG4_23|_SPL_P1|I_Q1|B _PG4_23|_SPL_P1|QA1 _PG4_23|_SPL_P1|I_Q1|MID  2e-12
I_PG4_23|_SPL_P1|I_Q1|B 0 _PG4_23|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG4_23|_SPL_P1|I_Q2|B _PG4_23|_SPL_P1|QB1 _PG4_23|_SPL_P1|I_Q2|MID  2e-12
I_PG4_23|_SPL_P1|I_Q2|B 0 _PG4_23|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG4_23|_SPL_P1|1|1 _PG4_23|_SPL_P1|D1 _PG4_23|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_P1|1|P _PG4_23|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG4_23|_SPL_P1|1|B _PG4_23|_SPL_P1|D1 _PG4_23|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_P1|1|RB _PG4_23|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_SPL_P1|2|1 _PG4_23|_SPL_P1|D2 _PG4_23|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_P1|2|P _PG4_23|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG4_23|_SPL_P1|2|B _PG4_23|_SPL_P1|D2 _PG4_23|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_P1|2|RB _PG4_23|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_SPL_P1|A|1 _PG4_23|_SPL_P1|QA1 _PG4_23|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_P1|A|P _PG4_23|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG4_23|_SPL_P1|A|B _PG4_23|_SPL_P1|QA1 _PG4_23|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_P1|A|RB _PG4_23|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_SPL_P1|B|1 _PG4_23|_SPL_P1|QB1 _PG4_23|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_SPL_P1|B|P _PG4_23|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG4_23|_SPL_P1|B|B _PG4_23|_SPL_P1|QB1 _PG4_23|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG4_23|_SPL_P1|B|RB _PG4_23|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_PG|I_A1|B _PG4_23|_PG|A1 _PG4_23|_PG|I_A1|MID  2e-12
I_PG4_23|_PG|I_A1|B 0 _PG4_23|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_PG|I_B1|B _PG4_23|_PG|B1 _PG4_23|_PG|I_B1|MID  2e-12
I_PG4_23|_PG|I_B1|B 0 _PG4_23|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_PG|I_Q3|B _PG4_23|_PG|Q3 _PG4_23|_PG|I_Q3|MID  2e-12
I_PG4_23|_PG|I_Q3|B 0 _PG4_23|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_23|_PG|I_Q2|B _PG4_23|_PG|Q2 _PG4_23|_PG|I_Q2|MID  2e-12
I_PG4_23|_PG|I_Q2|B 0 _PG4_23|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_PG|I_Q1|B _PG4_23|_PG|Q1 _PG4_23|_PG|I_Q1|MID  2e-12
I_PG4_23|_PG|I_Q1|B 0 _PG4_23|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_PG|A1|1 _PG4_23|_PG|A1 _PG4_23|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_PG|A1|P _PG4_23|_PG|A1|MID_SERIES 0  2e-13
R_PG4_23|_PG|A1|B _PG4_23|_PG|A1 _PG4_23|_PG|A1|MID_SHUNT  2.7439617672
L_PG4_23|_PG|A1|RB _PG4_23|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_PG|A2|1 _PG4_23|_PG|A2 _PG4_23|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_PG|A2|P _PG4_23|_PG|A2|MID_SERIES 0  2e-13
R_PG4_23|_PG|A2|B _PG4_23|_PG|A2 _PG4_23|_PG|A2|MID_SHUNT  2.7439617672
L_PG4_23|_PG|A2|RB _PG4_23|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_PG|A12|1 _PG4_23|_PG|A2 _PG4_23|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_PG|A12|B _PG4_23|_PG|A2 _PG4_23|_PG|A12|MID_SHUNT  3.84154647408
L_PG4_23|_PG|A12|RB _PG4_23|_PG|A12|MID_SHUNT _PG4_23|_PG|A3  2.1704737578552e-12
B_PG4_23|_PG|B1|1 _PG4_23|_PG|B1 _PG4_23|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_PG|B1|P _PG4_23|_PG|B1|MID_SERIES 0  2e-13
R_PG4_23|_PG|B1|B _PG4_23|_PG|B1 _PG4_23|_PG|B1|MID_SHUNT  2.7439617672
L_PG4_23|_PG|B1|RB _PG4_23|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_PG|B2|1 _PG4_23|_PG|B2 _PG4_23|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_PG|B2|P _PG4_23|_PG|B2|MID_SERIES 0  2e-13
R_PG4_23|_PG|B2|B _PG4_23|_PG|B2 _PG4_23|_PG|B2|MID_SHUNT  2.7439617672
L_PG4_23|_PG|B2|RB _PG4_23|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_PG|B12|1 _PG4_23|_PG|B2 _PG4_23|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG4_23|_PG|B12|B _PG4_23|_PG|B2 _PG4_23|_PG|B12|MID_SHUNT  3.84154647408
L_PG4_23|_PG|B12|RB _PG4_23|_PG|B12|MID_SHUNT _PG4_23|_PG|B3  2.1704737578552e-12
B_PG4_23|_PG|Q2|1 _PG4_23|_PG|Q2 _PG4_23|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_PG|Q2|P _PG4_23|_PG|Q2|MID_SERIES 0  2e-13
R_PG4_23|_PG|Q2|B _PG4_23|_PG|Q2 _PG4_23|_PG|Q2|MID_SHUNT  2.7439617672
L_PG4_23|_PG|Q2|RB _PG4_23|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_PG|Q1|1 _PG4_23|_PG|Q1 _PG4_23|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_PG|Q1|P _PG4_23|_PG|Q1|MID_SERIES 0  2e-13
R_PG4_23|_PG|Q1|B _PG4_23|_PG|Q1 _PG4_23|_PG|Q1|MID_SHUNT  2.7439617672
L_PG4_23|_PG|Q1|RB _PG4_23|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_GG|I_A1|B _PG4_23|_GG|A1 _PG4_23|_GG|I_A1|MID  2e-12
I_PG4_23|_GG|I_A1|B 0 _PG4_23|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_GG|I_B1|B _PG4_23|_GG|B1 _PG4_23|_GG|I_B1|MID  2e-12
I_PG4_23|_GG|I_B1|B 0 _PG4_23|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_GG|I_Q3|B _PG4_23|_GG|Q3 _PG4_23|_GG|I_Q3|MID  2e-12
I_PG4_23|_GG|I_Q3|B 0 _PG4_23|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_23|_GG|I_Q2|B _PG4_23|_GG|Q2 _PG4_23|_GG|I_Q2|MID  2e-12
I_PG4_23|_GG|I_Q2|B 0 _PG4_23|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_GG|I_Q1|B _PG4_23|_GG|Q1 _PG4_23|_GG|I_Q1|MID  2e-12
I_PG4_23|_GG|I_Q1|B 0 _PG4_23|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_GG|A1|1 _PG4_23|_GG|A1 _PG4_23|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_GG|A1|P _PG4_23|_GG|A1|MID_SERIES 0  2e-13
R_PG4_23|_GG|A1|B _PG4_23|_GG|A1 _PG4_23|_GG|A1|MID_SHUNT  2.7439617672
L_PG4_23|_GG|A1|RB _PG4_23|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_GG|A2|1 _PG4_23|_GG|A2 _PG4_23|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_GG|A2|P _PG4_23|_GG|A2|MID_SERIES 0  2e-13
R_PG4_23|_GG|A2|B _PG4_23|_GG|A2 _PG4_23|_GG|A2|MID_SHUNT  2.7439617672
L_PG4_23|_GG|A2|RB _PG4_23|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_GG|A12|1 _PG4_23|_GG|A2 _PG4_23|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_GG|A12|B _PG4_23|_GG|A2 _PG4_23|_GG|A12|MID_SHUNT  3.84154647408
L_PG4_23|_GG|A12|RB _PG4_23|_GG|A12|MID_SHUNT _PG4_23|_GG|A3  2.1704737578552e-12
B_PG4_23|_GG|B1|1 _PG4_23|_GG|B1 _PG4_23|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_GG|B1|P _PG4_23|_GG|B1|MID_SERIES 0  2e-13
R_PG4_23|_GG|B1|B _PG4_23|_GG|B1 _PG4_23|_GG|B1|MID_SHUNT  2.7439617672
L_PG4_23|_GG|B1|RB _PG4_23|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_GG|B2|1 _PG4_23|_GG|B2 _PG4_23|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_GG|B2|P _PG4_23|_GG|B2|MID_SERIES 0  2e-13
R_PG4_23|_GG|B2|B _PG4_23|_GG|B2 _PG4_23|_GG|B2|MID_SHUNT  2.7439617672
L_PG4_23|_GG|B2|RB _PG4_23|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_GG|B12|1 _PG4_23|_GG|B2 _PG4_23|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG4_23|_GG|B12|B _PG4_23|_GG|B2 _PG4_23|_GG|B12|MID_SHUNT  3.84154647408
L_PG4_23|_GG|B12|RB _PG4_23|_GG|B12|MID_SHUNT _PG4_23|_GG|B3  2.1704737578552e-12
B_PG4_23|_GG|Q2|1 _PG4_23|_GG|Q2 _PG4_23|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_GG|Q2|P _PG4_23|_GG|Q2|MID_SERIES 0  2e-13
R_PG4_23|_GG|Q2|B _PG4_23|_GG|Q2 _PG4_23|_GG|Q2|MID_SHUNT  2.7439617672
L_PG4_23|_GG|Q2|RB _PG4_23|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_GG|Q1|1 _PG4_23|_GG|Q1 _PG4_23|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_GG|Q1|P _PG4_23|_GG|Q1|MID_SERIES 0  2e-13
R_PG4_23|_GG|Q1|B _PG4_23|_GG|Q1 _PG4_23|_GG|Q1|MID_SHUNT  2.7439617672
L_PG4_23|_GG|Q1|RB _PG4_23|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_DFF_P0|I_1|B _PG4_23|_DFF_P0|A1 _PG4_23|_DFF_P0|I_1|MID  2e-12
I_PG4_23|_DFF_P0|I_1|B 0 _PG4_23|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_P0|I_3|B _PG4_23|_DFF_P0|A3 _PG4_23|_DFF_P0|I_3|MID  2e-12
I_PG4_23|_DFF_P0|I_3|B 0 _PG4_23|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_23|_DFF_P0|I_T|B _PG4_23|_DFF_P0|T1 _PG4_23|_DFF_P0|I_T|MID  2e-12
I_PG4_23|_DFF_P0|I_T|B 0 _PG4_23|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_P0|I_6|B _PG4_23|_DFF_P0|Q1 _PG4_23|_DFF_P0|I_6|MID  2e-12
I_PG4_23|_DFF_P0|I_6|B 0 _PG4_23|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_DFF_P0|1|1 _PG4_23|_DFF_P0|A1 _PG4_23|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P0|1|P _PG4_23|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P0|1|B _PG4_23|_DFF_P0|A1 _PG4_23|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P0|1|RB _PG4_23|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P0|23|1 _PG4_23|_DFF_P0|A2 _PG4_23|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_P0|23|B _PG4_23|_DFF_P0|A2 _PG4_23|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_P0|23|RB _PG4_23|_DFF_P0|23|MID_SHUNT _PG4_23|_DFF_P0|A3  2.1704737578552e-12
B_PG4_23|_DFF_P0|3|1 _PG4_23|_DFF_P0|A3 _PG4_23|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P0|3|P _PG4_23|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P0|3|B _PG4_23|_DFF_P0|A3 _PG4_23|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P0|3|RB _PG4_23|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P0|4|1 _PG4_23|_DFF_P0|A4 _PG4_23|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P0|4|P _PG4_23|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P0|4|B _PG4_23|_DFF_P0|A4 _PG4_23|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P0|4|RB _PG4_23|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P0|T|1 _PG4_23|_DFF_P0|T1 _PG4_23|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P0|T|P _PG4_23|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P0|T|B _PG4_23|_DFF_P0|T1 _PG4_23|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P0|T|RB _PG4_23|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P0|45|1 _PG4_23|_DFF_P0|T2 _PG4_23|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_P0|45|B _PG4_23|_DFF_P0|T2 _PG4_23|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_P0|45|RB _PG4_23|_DFF_P0|45|MID_SHUNT _PG4_23|_DFF_P0|A4  2.1704737578552e-12
B_PG4_23|_DFF_P0|6|1 _PG4_23|_DFF_P0|Q1 _PG4_23|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P0|6|P _PG4_23|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P0|6|B _PG4_23|_DFF_P0|Q1 _PG4_23|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P0|6|RB _PG4_23|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_DFF_P1|I_1|B _PG4_23|_DFF_P1|A1 _PG4_23|_DFF_P1|I_1|MID  2e-12
I_PG4_23|_DFF_P1|I_1|B 0 _PG4_23|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_P1|I_3|B _PG4_23|_DFF_P1|A3 _PG4_23|_DFF_P1|I_3|MID  2e-12
I_PG4_23|_DFF_P1|I_3|B 0 _PG4_23|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_23|_DFF_P1|I_T|B _PG4_23|_DFF_P1|T1 _PG4_23|_DFF_P1|I_T|MID  2e-12
I_PG4_23|_DFF_P1|I_T|B 0 _PG4_23|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_P1|I_6|B _PG4_23|_DFF_P1|Q1 _PG4_23|_DFF_P1|I_6|MID  2e-12
I_PG4_23|_DFF_P1|I_6|B 0 _PG4_23|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_DFF_P1|1|1 _PG4_23|_DFF_P1|A1 _PG4_23|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P1|1|P _PG4_23|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P1|1|B _PG4_23|_DFF_P1|A1 _PG4_23|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P1|1|RB _PG4_23|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P1|23|1 _PG4_23|_DFF_P1|A2 _PG4_23|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_P1|23|B _PG4_23|_DFF_P1|A2 _PG4_23|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_P1|23|RB _PG4_23|_DFF_P1|23|MID_SHUNT _PG4_23|_DFF_P1|A3  2.1704737578552e-12
B_PG4_23|_DFF_P1|3|1 _PG4_23|_DFF_P1|A3 _PG4_23|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P1|3|P _PG4_23|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P1|3|B _PG4_23|_DFF_P1|A3 _PG4_23|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P1|3|RB _PG4_23|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P1|4|1 _PG4_23|_DFF_P1|A4 _PG4_23|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P1|4|P _PG4_23|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P1|4|B _PG4_23|_DFF_P1|A4 _PG4_23|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P1|4|RB _PG4_23|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P1|T|1 _PG4_23|_DFF_P1|T1 _PG4_23|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P1|T|P _PG4_23|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P1|T|B _PG4_23|_DFF_P1|T1 _PG4_23|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P1|T|RB _PG4_23|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_P1|45|1 _PG4_23|_DFF_P1|T2 _PG4_23|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_P1|45|B _PG4_23|_DFF_P1|T2 _PG4_23|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_P1|45|RB _PG4_23|_DFF_P1|45|MID_SHUNT _PG4_23|_DFF_P1|A4  2.1704737578552e-12
B_PG4_23|_DFF_P1|6|1 _PG4_23|_DFF_P1|Q1 _PG4_23|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_P1|6|P _PG4_23|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG4_23|_DFF_P1|6|B _PG4_23|_DFF_P1|Q1 _PG4_23|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_P1|6|RB _PG4_23|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_DFF_PG|I_1|B _PG4_23|_DFF_PG|A1 _PG4_23|_DFF_PG|I_1|MID  2e-12
I_PG4_23|_DFF_PG|I_1|B 0 _PG4_23|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_PG|I_3|B _PG4_23|_DFF_PG|A3 _PG4_23|_DFF_PG|I_3|MID  2e-12
I_PG4_23|_DFF_PG|I_3|B 0 _PG4_23|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_23|_DFF_PG|I_T|B _PG4_23|_DFF_PG|T1 _PG4_23|_DFF_PG|I_T|MID  2e-12
I_PG4_23|_DFF_PG|I_T|B 0 _PG4_23|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_PG|I_6|B _PG4_23|_DFF_PG|Q1 _PG4_23|_DFF_PG|I_6|MID  2e-12
I_PG4_23|_DFF_PG|I_6|B 0 _PG4_23|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_DFF_PG|1|1 _PG4_23|_DFF_PG|A1 _PG4_23|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_PG|1|P _PG4_23|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG4_23|_DFF_PG|1|B _PG4_23|_DFF_PG|A1 _PG4_23|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_PG|1|RB _PG4_23|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_PG|23|1 _PG4_23|_DFF_PG|A2 _PG4_23|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_PG|23|B _PG4_23|_DFF_PG|A2 _PG4_23|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_PG|23|RB _PG4_23|_DFF_PG|23|MID_SHUNT _PG4_23|_DFF_PG|A3  2.1704737578552e-12
B_PG4_23|_DFF_PG|3|1 _PG4_23|_DFF_PG|A3 _PG4_23|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_PG|3|P _PG4_23|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG4_23|_DFF_PG|3|B _PG4_23|_DFF_PG|A3 _PG4_23|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_PG|3|RB _PG4_23|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_PG|4|1 _PG4_23|_DFF_PG|A4 _PG4_23|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_PG|4|P _PG4_23|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG4_23|_DFF_PG|4|B _PG4_23|_DFF_PG|A4 _PG4_23|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_PG|4|RB _PG4_23|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_PG|T|1 _PG4_23|_DFF_PG|T1 _PG4_23|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_PG|T|P _PG4_23|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG4_23|_DFF_PG|T|B _PG4_23|_DFF_PG|T1 _PG4_23|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_PG|T|RB _PG4_23|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_PG|45|1 _PG4_23|_DFF_PG|T2 _PG4_23|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_PG|45|B _PG4_23|_DFF_PG|T2 _PG4_23|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_PG|45|RB _PG4_23|_DFF_PG|45|MID_SHUNT _PG4_23|_DFF_PG|A4  2.1704737578552e-12
B_PG4_23|_DFF_PG|6|1 _PG4_23|_DFF_PG|Q1 _PG4_23|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_PG|6|P _PG4_23|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG4_23|_DFF_PG|6|B _PG4_23|_DFF_PG|Q1 _PG4_23|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_PG|6|RB _PG4_23|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_DFF_GG|I_1|B _PG4_23|_DFF_GG|A1 _PG4_23|_DFF_GG|I_1|MID  2e-12
I_PG4_23|_DFF_GG|I_1|B 0 _PG4_23|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_GG|I_3|B _PG4_23|_DFF_GG|A3 _PG4_23|_DFF_GG|I_3|MID  2e-12
I_PG4_23|_DFF_GG|I_3|B 0 _PG4_23|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG4_23|_DFF_GG|I_T|B _PG4_23|_DFF_GG|T1 _PG4_23|_DFF_GG|I_T|MID  2e-12
I_PG4_23|_DFF_GG|I_T|B 0 _PG4_23|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_DFF_GG|I_6|B _PG4_23|_DFF_GG|Q1 _PG4_23|_DFF_GG|I_6|MID  2e-12
I_PG4_23|_DFF_GG|I_6|B 0 _PG4_23|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_DFF_GG|1|1 _PG4_23|_DFF_GG|A1 _PG4_23|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_GG|1|P _PG4_23|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG4_23|_DFF_GG|1|B _PG4_23|_DFF_GG|A1 _PG4_23|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_GG|1|RB _PG4_23|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_GG|23|1 _PG4_23|_DFF_GG|A2 _PG4_23|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_GG|23|B _PG4_23|_DFF_GG|A2 _PG4_23|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_GG|23|RB _PG4_23|_DFF_GG|23|MID_SHUNT _PG4_23|_DFF_GG|A3  2.1704737578552e-12
B_PG4_23|_DFF_GG|3|1 _PG4_23|_DFF_GG|A3 _PG4_23|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_GG|3|P _PG4_23|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG4_23|_DFF_GG|3|B _PG4_23|_DFF_GG|A3 _PG4_23|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_GG|3|RB _PG4_23|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_GG|4|1 _PG4_23|_DFF_GG|A4 _PG4_23|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_GG|4|P _PG4_23|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG4_23|_DFF_GG|4|B _PG4_23|_DFF_GG|A4 _PG4_23|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_GG|4|RB _PG4_23|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_GG|T|1 _PG4_23|_DFF_GG|T1 _PG4_23|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_GG|T|P _PG4_23|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG4_23|_DFF_GG|T|B _PG4_23|_DFF_GG|T1 _PG4_23|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_GG|T|RB _PG4_23|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_DFF_GG|45|1 _PG4_23|_DFF_GG|T2 _PG4_23|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG4_23|_DFF_GG|45|B _PG4_23|_DFF_GG|T2 _PG4_23|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG4_23|_DFF_GG|45|RB _PG4_23|_DFF_GG|45|MID_SHUNT _PG4_23|_DFF_GG|A4  2.1704737578552e-12
B_PG4_23|_DFF_GG|6|1 _PG4_23|_DFF_GG|Q1 _PG4_23|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_DFF_GG|6|P _PG4_23|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG4_23|_DFF_GG|6|B _PG4_23|_DFF_GG|Q1 _PG4_23|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG4_23|_DFF_GG|6|RB _PG4_23|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_AND_G|I_A1|B _PG4_23|_AND_G|A1 _PG4_23|_AND_G|I_A1|MID  2e-12
I_PG4_23|_AND_G|I_A1|B 0 _PG4_23|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_AND_G|I_B1|B _PG4_23|_AND_G|B1 _PG4_23|_AND_G|I_B1|MID  2e-12
I_PG4_23|_AND_G|I_B1|B 0 _PG4_23|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_AND_G|I_Q3|B _PG4_23|_AND_G|Q3 _PG4_23|_AND_G|I_Q3|MID  2e-12
I_PG4_23|_AND_G|I_Q3|B 0 _PG4_23|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG4_23|_AND_G|I_Q2|B _PG4_23|_AND_G|Q2 _PG4_23|_AND_G|I_Q2|MID  2e-12
I_PG4_23|_AND_G|I_Q2|B 0 _PG4_23|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_AND_G|I_Q1|B _PG4_23|_AND_G|Q1 _PG4_23|_AND_G|I_Q1|MID  2e-12
I_PG4_23|_AND_G|I_Q1|B 0 _PG4_23|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_AND_G|A1|1 _PG4_23|_AND_G|A1 _PG4_23|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_G|A1|P _PG4_23|_AND_G|A1|MID_SERIES 0  2e-13
R_PG4_23|_AND_G|A1|B _PG4_23|_AND_G|A1 _PG4_23|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG4_23|_AND_G|A1|RB _PG4_23|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_G|A2|1 _PG4_23|_AND_G|A2 _PG4_23|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_G|A2|P _PG4_23|_AND_G|A2|MID_SERIES 0  2e-13
R_PG4_23|_AND_G|A2|B _PG4_23|_AND_G|A2 _PG4_23|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG4_23|_AND_G|A2|RB _PG4_23|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_G|A12|1 _PG4_23|_AND_G|A2 _PG4_23|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_AND_G|A12|B _PG4_23|_AND_G|A2 _PG4_23|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG4_23|_AND_G|A12|RB _PG4_23|_AND_G|A12|MID_SHUNT _PG4_23|_AND_G|A3  2.1704737578552e-12
B_PG4_23|_AND_G|B1|1 _PG4_23|_AND_G|B1 _PG4_23|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_G|B1|P _PG4_23|_AND_G|B1|MID_SERIES 0  2e-13
R_PG4_23|_AND_G|B1|B _PG4_23|_AND_G|B1 _PG4_23|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG4_23|_AND_G|B1|RB _PG4_23|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_G|B2|1 _PG4_23|_AND_G|B2 _PG4_23|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_G|B2|P _PG4_23|_AND_G|B2|MID_SERIES 0  2e-13
R_PG4_23|_AND_G|B2|B _PG4_23|_AND_G|B2 _PG4_23|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG4_23|_AND_G|B2|RB _PG4_23|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_G|B12|1 _PG4_23|_AND_G|B2 _PG4_23|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG4_23|_AND_G|B12|B _PG4_23|_AND_G|B2 _PG4_23|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG4_23|_AND_G|B12|RB _PG4_23|_AND_G|B12|MID_SHUNT _PG4_23|_AND_G|B3  2.1704737578552e-12
B_PG4_23|_AND_G|Q2|1 _PG4_23|_AND_G|Q2 _PG4_23|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_G|Q2|P _PG4_23|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG4_23|_AND_G|Q2|B _PG4_23|_AND_G|Q2 _PG4_23|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG4_23|_AND_G|Q2|RB _PG4_23|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_G|Q1|1 _PG4_23|_AND_G|Q1 _PG4_23|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_G|Q1|P _PG4_23|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG4_23|_AND_G|Q1|B _PG4_23|_AND_G|Q1 _PG4_23|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG4_23|_AND_G|Q1|RB _PG4_23|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG4_23|_AND_P|I_A1|B _PG4_23|_AND_P|A1 _PG4_23|_AND_P|I_A1|MID  2e-12
I_PG4_23|_AND_P|I_A1|B 0 _PG4_23|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_AND_P|I_B1|B _PG4_23|_AND_P|B1 _PG4_23|_AND_P|I_B1|MID  2e-12
I_PG4_23|_AND_P|I_B1|B 0 _PG4_23|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_AND_P|I_Q3|B _PG4_23|_AND_P|Q3 _PG4_23|_AND_P|I_Q3|MID  2e-12
I_PG4_23|_AND_P|I_Q3|B 0 _PG4_23|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG4_23|_AND_P|I_Q2|B _PG4_23|_AND_P|Q2 _PG4_23|_AND_P|I_Q2|MID  2e-12
I_PG4_23|_AND_P|I_Q2|B 0 _PG4_23|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG4_23|_AND_P|I_Q1|B _PG4_23|_AND_P|Q1 _PG4_23|_AND_P|I_Q1|MID  2e-12
I_PG4_23|_AND_P|I_Q1|B 0 _PG4_23|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG4_23|_AND_P|A1|1 _PG4_23|_AND_P|A1 _PG4_23|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_P|A1|P _PG4_23|_AND_P|A1|MID_SERIES 0  2e-13
R_PG4_23|_AND_P|A1|B _PG4_23|_AND_P|A1 _PG4_23|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG4_23|_AND_P|A1|RB _PG4_23|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_P|A2|1 _PG4_23|_AND_P|A2 _PG4_23|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_P|A2|P _PG4_23|_AND_P|A2|MID_SERIES 0  2e-13
R_PG4_23|_AND_P|A2|B _PG4_23|_AND_P|A2 _PG4_23|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG4_23|_AND_P|A2|RB _PG4_23|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_P|A12|1 _PG4_23|_AND_P|A2 _PG4_23|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG4_23|_AND_P|A12|B _PG4_23|_AND_P|A2 _PG4_23|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG4_23|_AND_P|A12|RB _PG4_23|_AND_P|A12|MID_SHUNT _PG4_23|_AND_P|A3  2.1704737578552e-12
B_PG4_23|_AND_P|B1|1 _PG4_23|_AND_P|B1 _PG4_23|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_P|B1|P _PG4_23|_AND_P|B1|MID_SERIES 0  2e-13
R_PG4_23|_AND_P|B1|B _PG4_23|_AND_P|B1 _PG4_23|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG4_23|_AND_P|B1|RB _PG4_23|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_P|B2|1 _PG4_23|_AND_P|B2 _PG4_23|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_P|B2|P _PG4_23|_AND_P|B2|MID_SERIES 0  2e-13
R_PG4_23|_AND_P|B2|B _PG4_23|_AND_P|B2 _PG4_23|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG4_23|_AND_P|B2|RB _PG4_23|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_P|B12|1 _PG4_23|_AND_P|B2 _PG4_23|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG4_23|_AND_P|B12|B _PG4_23|_AND_P|B2 _PG4_23|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG4_23|_AND_P|B12|RB _PG4_23|_AND_P|B12|MID_SHUNT _PG4_23|_AND_P|B3  2.1704737578552e-12
B_PG4_23|_AND_P|Q2|1 _PG4_23|_AND_P|Q2 _PG4_23|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_P|Q2|P _PG4_23|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG4_23|_AND_P|Q2|B _PG4_23|_AND_P|Q2 _PG4_23|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG4_23|_AND_P|Q2|RB _PG4_23|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG4_23|_AND_P|Q1|1 _PG4_23|_AND_P|Q1 _PG4_23|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG4_23|_AND_P|Q1|P _PG4_23|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG4_23|_AND_P|Q1|B _PG4_23|_AND_P|Q1 _PG4_23|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG4_23|_AND_P|Q1|RB _PG4_23|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_SPL_G1|I_D1|B _PG5_23|_SPL_G1|D1 _PG5_23|_SPL_G1|I_D1|MID  2e-12
I_PG5_23|_SPL_G1|I_D1|B 0 _PG5_23|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_23|_SPL_G1|I_D2|B _PG5_23|_SPL_G1|D2 _PG5_23|_SPL_G1|I_D2|MID  2e-12
I_PG5_23|_SPL_G1|I_D2|B 0 _PG5_23|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG5_23|_SPL_G1|I_Q1|B _PG5_23|_SPL_G1|QA1 _PG5_23|_SPL_G1|I_Q1|MID  2e-12
I_PG5_23|_SPL_G1|I_Q1|B 0 _PG5_23|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_23|_SPL_G1|I_Q2|B _PG5_23|_SPL_G1|QB1 _PG5_23|_SPL_G1|I_Q2|MID  2e-12
I_PG5_23|_SPL_G1|I_Q2|B 0 _PG5_23|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG5_23|_SPL_G1|1|1 _PG5_23|_SPL_G1|D1 _PG5_23|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_G1|1|P _PG5_23|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG5_23|_SPL_G1|1|B _PG5_23|_SPL_G1|D1 _PG5_23|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_G1|1|RB _PG5_23|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_SPL_G1|2|1 _PG5_23|_SPL_G1|D2 _PG5_23|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_G1|2|P _PG5_23|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG5_23|_SPL_G1|2|B _PG5_23|_SPL_G1|D2 _PG5_23|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_G1|2|RB _PG5_23|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_SPL_G1|A|1 _PG5_23|_SPL_G1|QA1 _PG5_23|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_G1|A|P _PG5_23|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG5_23|_SPL_G1|A|B _PG5_23|_SPL_G1|QA1 _PG5_23|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_G1|A|RB _PG5_23|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_SPL_G1|B|1 _PG5_23|_SPL_G1|QB1 _PG5_23|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_G1|B|P _PG5_23|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG5_23|_SPL_G1|B|B _PG5_23|_SPL_G1|QB1 _PG5_23|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_G1|B|RB _PG5_23|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_SPL_P1|I_D1|B _PG5_23|_SPL_P1|D1 _PG5_23|_SPL_P1|I_D1|MID  2e-12
I_PG5_23|_SPL_P1|I_D1|B 0 _PG5_23|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_23|_SPL_P1|I_D2|B _PG5_23|_SPL_P1|D2 _PG5_23|_SPL_P1|I_D2|MID  2e-12
I_PG5_23|_SPL_P1|I_D2|B 0 _PG5_23|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG5_23|_SPL_P1|I_Q1|B _PG5_23|_SPL_P1|QA1 _PG5_23|_SPL_P1|I_Q1|MID  2e-12
I_PG5_23|_SPL_P1|I_Q1|B 0 _PG5_23|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG5_23|_SPL_P1|I_Q2|B _PG5_23|_SPL_P1|QB1 _PG5_23|_SPL_P1|I_Q2|MID  2e-12
I_PG5_23|_SPL_P1|I_Q2|B 0 _PG5_23|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG5_23|_SPL_P1|1|1 _PG5_23|_SPL_P1|D1 _PG5_23|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_P1|1|P _PG5_23|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG5_23|_SPL_P1|1|B _PG5_23|_SPL_P1|D1 _PG5_23|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_P1|1|RB _PG5_23|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_SPL_P1|2|1 _PG5_23|_SPL_P1|D2 _PG5_23|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_P1|2|P _PG5_23|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG5_23|_SPL_P1|2|B _PG5_23|_SPL_P1|D2 _PG5_23|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_P1|2|RB _PG5_23|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_SPL_P1|A|1 _PG5_23|_SPL_P1|QA1 _PG5_23|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_P1|A|P _PG5_23|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG5_23|_SPL_P1|A|B _PG5_23|_SPL_P1|QA1 _PG5_23|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_P1|A|RB _PG5_23|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_SPL_P1|B|1 _PG5_23|_SPL_P1|QB1 _PG5_23|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_SPL_P1|B|P _PG5_23|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG5_23|_SPL_P1|B|B _PG5_23|_SPL_P1|QB1 _PG5_23|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG5_23|_SPL_P1|B|RB _PG5_23|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_PG|I_A1|B _PG5_23|_PG|A1 _PG5_23|_PG|I_A1|MID  2e-12
I_PG5_23|_PG|I_A1|B 0 _PG5_23|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_PG|I_B1|B _PG5_23|_PG|B1 _PG5_23|_PG|I_B1|MID  2e-12
I_PG5_23|_PG|I_B1|B 0 _PG5_23|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_PG|I_Q3|B _PG5_23|_PG|Q3 _PG5_23|_PG|I_Q3|MID  2e-12
I_PG5_23|_PG|I_Q3|B 0 _PG5_23|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_23|_PG|I_Q2|B _PG5_23|_PG|Q2 _PG5_23|_PG|I_Q2|MID  2e-12
I_PG5_23|_PG|I_Q2|B 0 _PG5_23|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_PG|I_Q1|B _PG5_23|_PG|Q1 _PG5_23|_PG|I_Q1|MID  2e-12
I_PG5_23|_PG|I_Q1|B 0 _PG5_23|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_PG|A1|1 _PG5_23|_PG|A1 _PG5_23|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_PG|A1|P _PG5_23|_PG|A1|MID_SERIES 0  2e-13
R_PG5_23|_PG|A1|B _PG5_23|_PG|A1 _PG5_23|_PG|A1|MID_SHUNT  2.7439617672
L_PG5_23|_PG|A1|RB _PG5_23|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_PG|A2|1 _PG5_23|_PG|A2 _PG5_23|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_PG|A2|P _PG5_23|_PG|A2|MID_SERIES 0  2e-13
R_PG5_23|_PG|A2|B _PG5_23|_PG|A2 _PG5_23|_PG|A2|MID_SHUNT  2.7439617672
L_PG5_23|_PG|A2|RB _PG5_23|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_PG|A12|1 _PG5_23|_PG|A2 _PG5_23|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_PG|A12|B _PG5_23|_PG|A2 _PG5_23|_PG|A12|MID_SHUNT  3.84154647408
L_PG5_23|_PG|A12|RB _PG5_23|_PG|A12|MID_SHUNT _PG5_23|_PG|A3  2.1704737578552e-12
B_PG5_23|_PG|B1|1 _PG5_23|_PG|B1 _PG5_23|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_PG|B1|P _PG5_23|_PG|B1|MID_SERIES 0  2e-13
R_PG5_23|_PG|B1|B _PG5_23|_PG|B1 _PG5_23|_PG|B1|MID_SHUNT  2.7439617672
L_PG5_23|_PG|B1|RB _PG5_23|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_PG|B2|1 _PG5_23|_PG|B2 _PG5_23|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_PG|B2|P _PG5_23|_PG|B2|MID_SERIES 0  2e-13
R_PG5_23|_PG|B2|B _PG5_23|_PG|B2 _PG5_23|_PG|B2|MID_SHUNT  2.7439617672
L_PG5_23|_PG|B2|RB _PG5_23|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_PG|B12|1 _PG5_23|_PG|B2 _PG5_23|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG5_23|_PG|B12|B _PG5_23|_PG|B2 _PG5_23|_PG|B12|MID_SHUNT  3.84154647408
L_PG5_23|_PG|B12|RB _PG5_23|_PG|B12|MID_SHUNT _PG5_23|_PG|B3  2.1704737578552e-12
B_PG5_23|_PG|Q2|1 _PG5_23|_PG|Q2 _PG5_23|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_PG|Q2|P _PG5_23|_PG|Q2|MID_SERIES 0  2e-13
R_PG5_23|_PG|Q2|B _PG5_23|_PG|Q2 _PG5_23|_PG|Q2|MID_SHUNT  2.7439617672
L_PG5_23|_PG|Q2|RB _PG5_23|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_PG|Q1|1 _PG5_23|_PG|Q1 _PG5_23|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_PG|Q1|P _PG5_23|_PG|Q1|MID_SERIES 0  2e-13
R_PG5_23|_PG|Q1|B _PG5_23|_PG|Q1 _PG5_23|_PG|Q1|MID_SHUNT  2.7439617672
L_PG5_23|_PG|Q1|RB _PG5_23|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_GG|I_A1|B _PG5_23|_GG|A1 _PG5_23|_GG|I_A1|MID  2e-12
I_PG5_23|_GG|I_A1|B 0 _PG5_23|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_GG|I_B1|B _PG5_23|_GG|B1 _PG5_23|_GG|I_B1|MID  2e-12
I_PG5_23|_GG|I_B1|B 0 _PG5_23|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_GG|I_Q3|B _PG5_23|_GG|Q3 _PG5_23|_GG|I_Q3|MID  2e-12
I_PG5_23|_GG|I_Q3|B 0 _PG5_23|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_23|_GG|I_Q2|B _PG5_23|_GG|Q2 _PG5_23|_GG|I_Q2|MID  2e-12
I_PG5_23|_GG|I_Q2|B 0 _PG5_23|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_GG|I_Q1|B _PG5_23|_GG|Q1 _PG5_23|_GG|I_Q1|MID  2e-12
I_PG5_23|_GG|I_Q1|B 0 _PG5_23|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_GG|A1|1 _PG5_23|_GG|A1 _PG5_23|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_GG|A1|P _PG5_23|_GG|A1|MID_SERIES 0  2e-13
R_PG5_23|_GG|A1|B _PG5_23|_GG|A1 _PG5_23|_GG|A1|MID_SHUNT  2.7439617672
L_PG5_23|_GG|A1|RB _PG5_23|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_GG|A2|1 _PG5_23|_GG|A2 _PG5_23|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_GG|A2|P _PG5_23|_GG|A2|MID_SERIES 0  2e-13
R_PG5_23|_GG|A2|B _PG5_23|_GG|A2 _PG5_23|_GG|A2|MID_SHUNT  2.7439617672
L_PG5_23|_GG|A2|RB _PG5_23|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_GG|A12|1 _PG5_23|_GG|A2 _PG5_23|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_GG|A12|B _PG5_23|_GG|A2 _PG5_23|_GG|A12|MID_SHUNT  3.84154647408
L_PG5_23|_GG|A12|RB _PG5_23|_GG|A12|MID_SHUNT _PG5_23|_GG|A3  2.1704737578552e-12
B_PG5_23|_GG|B1|1 _PG5_23|_GG|B1 _PG5_23|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_GG|B1|P _PG5_23|_GG|B1|MID_SERIES 0  2e-13
R_PG5_23|_GG|B1|B _PG5_23|_GG|B1 _PG5_23|_GG|B1|MID_SHUNT  2.7439617672
L_PG5_23|_GG|B1|RB _PG5_23|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_GG|B2|1 _PG5_23|_GG|B2 _PG5_23|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_GG|B2|P _PG5_23|_GG|B2|MID_SERIES 0  2e-13
R_PG5_23|_GG|B2|B _PG5_23|_GG|B2 _PG5_23|_GG|B2|MID_SHUNT  2.7439617672
L_PG5_23|_GG|B2|RB _PG5_23|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_GG|B12|1 _PG5_23|_GG|B2 _PG5_23|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG5_23|_GG|B12|B _PG5_23|_GG|B2 _PG5_23|_GG|B12|MID_SHUNT  3.84154647408
L_PG5_23|_GG|B12|RB _PG5_23|_GG|B12|MID_SHUNT _PG5_23|_GG|B3  2.1704737578552e-12
B_PG5_23|_GG|Q2|1 _PG5_23|_GG|Q2 _PG5_23|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_GG|Q2|P _PG5_23|_GG|Q2|MID_SERIES 0  2e-13
R_PG5_23|_GG|Q2|B _PG5_23|_GG|Q2 _PG5_23|_GG|Q2|MID_SHUNT  2.7439617672
L_PG5_23|_GG|Q2|RB _PG5_23|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_GG|Q1|1 _PG5_23|_GG|Q1 _PG5_23|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_GG|Q1|P _PG5_23|_GG|Q1|MID_SERIES 0  2e-13
R_PG5_23|_GG|Q1|B _PG5_23|_GG|Q1 _PG5_23|_GG|Q1|MID_SHUNT  2.7439617672
L_PG5_23|_GG|Q1|RB _PG5_23|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_DFF_P0|I_1|B _PG5_23|_DFF_P0|A1 _PG5_23|_DFF_P0|I_1|MID  2e-12
I_PG5_23|_DFF_P0|I_1|B 0 _PG5_23|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_P0|I_3|B _PG5_23|_DFF_P0|A3 _PG5_23|_DFF_P0|I_3|MID  2e-12
I_PG5_23|_DFF_P0|I_3|B 0 _PG5_23|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_23|_DFF_P0|I_T|B _PG5_23|_DFF_P0|T1 _PG5_23|_DFF_P0|I_T|MID  2e-12
I_PG5_23|_DFF_P0|I_T|B 0 _PG5_23|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_P0|I_6|B _PG5_23|_DFF_P0|Q1 _PG5_23|_DFF_P0|I_6|MID  2e-12
I_PG5_23|_DFF_P0|I_6|B 0 _PG5_23|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_DFF_P0|1|1 _PG5_23|_DFF_P0|A1 _PG5_23|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P0|1|P _PG5_23|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P0|1|B _PG5_23|_DFF_P0|A1 _PG5_23|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P0|1|RB _PG5_23|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P0|23|1 _PG5_23|_DFF_P0|A2 _PG5_23|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_P0|23|B _PG5_23|_DFF_P0|A2 _PG5_23|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_P0|23|RB _PG5_23|_DFF_P0|23|MID_SHUNT _PG5_23|_DFF_P0|A3  2.1704737578552e-12
B_PG5_23|_DFF_P0|3|1 _PG5_23|_DFF_P0|A3 _PG5_23|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P0|3|P _PG5_23|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P0|3|B _PG5_23|_DFF_P0|A3 _PG5_23|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P0|3|RB _PG5_23|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P0|4|1 _PG5_23|_DFF_P0|A4 _PG5_23|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P0|4|P _PG5_23|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P0|4|B _PG5_23|_DFF_P0|A4 _PG5_23|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P0|4|RB _PG5_23|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P0|T|1 _PG5_23|_DFF_P0|T1 _PG5_23|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P0|T|P _PG5_23|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P0|T|B _PG5_23|_DFF_P0|T1 _PG5_23|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P0|T|RB _PG5_23|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P0|45|1 _PG5_23|_DFF_P0|T2 _PG5_23|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_P0|45|B _PG5_23|_DFF_P0|T2 _PG5_23|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_P0|45|RB _PG5_23|_DFF_P0|45|MID_SHUNT _PG5_23|_DFF_P0|A4  2.1704737578552e-12
B_PG5_23|_DFF_P0|6|1 _PG5_23|_DFF_P0|Q1 _PG5_23|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P0|6|P _PG5_23|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P0|6|B _PG5_23|_DFF_P0|Q1 _PG5_23|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P0|6|RB _PG5_23|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_DFF_P1|I_1|B _PG5_23|_DFF_P1|A1 _PG5_23|_DFF_P1|I_1|MID  2e-12
I_PG5_23|_DFF_P1|I_1|B 0 _PG5_23|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_P1|I_3|B _PG5_23|_DFF_P1|A3 _PG5_23|_DFF_P1|I_3|MID  2e-12
I_PG5_23|_DFF_P1|I_3|B 0 _PG5_23|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_23|_DFF_P1|I_T|B _PG5_23|_DFF_P1|T1 _PG5_23|_DFF_P1|I_T|MID  2e-12
I_PG5_23|_DFF_P1|I_T|B 0 _PG5_23|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_P1|I_6|B _PG5_23|_DFF_P1|Q1 _PG5_23|_DFF_P1|I_6|MID  2e-12
I_PG5_23|_DFF_P1|I_6|B 0 _PG5_23|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_DFF_P1|1|1 _PG5_23|_DFF_P1|A1 _PG5_23|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P1|1|P _PG5_23|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P1|1|B _PG5_23|_DFF_P1|A1 _PG5_23|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P1|1|RB _PG5_23|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P1|23|1 _PG5_23|_DFF_P1|A2 _PG5_23|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_P1|23|B _PG5_23|_DFF_P1|A2 _PG5_23|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_P1|23|RB _PG5_23|_DFF_P1|23|MID_SHUNT _PG5_23|_DFF_P1|A3  2.1704737578552e-12
B_PG5_23|_DFF_P1|3|1 _PG5_23|_DFF_P1|A3 _PG5_23|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P1|3|P _PG5_23|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P1|3|B _PG5_23|_DFF_P1|A3 _PG5_23|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P1|3|RB _PG5_23|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P1|4|1 _PG5_23|_DFF_P1|A4 _PG5_23|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P1|4|P _PG5_23|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P1|4|B _PG5_23|_DFF_P1|A4 _PG5_23|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P1|4|RB _PG5_23|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P1|T|1 _PG5_23|_DFF_P1|T1 _PG5_23|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P1|T|P _PG5_23|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P1|T|B _PG5_23|_DFF_P1|T1 _PG5_23|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P1|T|RB _PG5_23|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_P1|45|1 _PG5_23|_DFF_P1|T2 _PG5_23|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_P1|45|B _PG5_23|_DFF_P1|T2 _PG5_23|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_P1|45|RB _PG5_23|_DFF_P1|45|MID_SHUNT _PG5_23|_DFF_P1|A4  2.1704737578552e-12
B_PG5_23|_DFF_P1|6|1 _PG5_23|_DFF_P1|Q1 _PG5_23|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_P1|6|P _PG5_23|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG5_23|_DFF_P1|6|B _PG5_23|_DFF_P1|Q1 _PG5_23|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_P1|6|RB _PG5_23|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_DFF_PG|I_1|B _PG5_23|_DFF_PG|A1 _PG5_23|_DFF_PG|I_1|MID  2e-12
I_PG5_23|_DFF_PG|I_1|B 0 _PG5_23|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_PG|I_3|B _PG5_23|_DFF_PG|A3 _PG5_23|_DFF_PG|I_3|MID  2e-12
I_PG5_23|_DFF_PG|I_3|B 0 _PG5_23|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_23|_DFF_PG|I_T|B _PG5_23|_DFF_PG|T1 _PG5_23|_DFF_PG|I_T|MID  2e-12
I_PG5_23|_DFF_PG|I_T|B 0 _PG5_23|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_PG|I_6|B _PG5_23|_DFF_PG|Q1 _PG5_23|_DFF_PG|I_6|MID  2e-12
I_PG5_23|_DFF_PG|I_6|B 0 _PG5_23|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_DFF_PG|1|1 _PG5_23|_DFF_PG|A1 _PG5_23|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_PG|1|P _PG5_23|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG5_23|_DFF_PG|1|B _PG5_23|_DFF_PG|A1 _PG5_23|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_PG|1|RB _PG5_23|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_PG|23|1 _PG5_23|_DFF_PG|A2 _PG5_23|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_PG|23|B _PG5_23|_DFF_PG|A2 _PG5_23|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_PG|23|RB _PG5_23|_DFF_PG|23|MID_SHUNT _PG5_23|_DFF_PG|A3  2.1704737578552e-12
B_PG5_23|_DFF_PG|3|1 _PG5_23|_DFF_PG|A3 _PG5_23|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_PG|3|P _PG5_23|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG5_23|_DFF_PG|3|B _PG5_23|_DFF_PG|A3 _PG5_23|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_PG|3|RB _PG5_23|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_PG|4|1 _PG5_23|_DFF_PG|A4 _PG5_23|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_PG|4|P _PG5_23|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG5_23|_DFF_PG|4|B _PG5_23|_DFF_PG|A4 _PG5_23|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_PG|4|RB _PG5_23|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_PG|T|1 _PG5_23|_DFF_PG|T1 _PG5_23|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_PG|T|P _PG5_23|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG5_23|_DFF_PG|T|B _PG5_23|_DFF_PG|T1 _PG5_23|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_PG|T|RB _PG5_23|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_PG|45|1 _PG5_23|_DFF_PG|T2 _PG5_23|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_PG|45|B _PG5_23|_DFF_PG|T2 _PG5_23|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_PG|45|RB _PG5_23|_DFF_PG|45|MID_SHUNT _PG5_23|_DFF_PG|A4  2.1704737578552e-12
B_PG5_23|_DFF_PG|6|1 _PG5_23|_DFF_PG|Q1 _PG5_23|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_PG|6|P _PG5_23|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG5_23|_DFF_PG|6|B _PG5_23|_DFF_PG|Q1 _PG5_23|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_PG|6|RB _PG5_23|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_DFF_GG|I_1|B _PG5_23|_DFF_GG|A1 _PG5_23|_DFF_GG|I_1|MID  2e-12
I_PG5_23|_DFF_GG|I_1|B 0 _PG5_23|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_GG|I_3|B _PG5_23|_DFF_GG|A3 _PG5_23|_DFF_GG|I_3|MID  2e-12
I_PG5_23|_DFF_GG|I_3|B 0 _PG5_23|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG5_23|_DFF_GG|I_T|B _PG5_23|_DFF_GG|T1 _PG5_23|_DFF_GG|I_T|MID  2e-12
I_PG5_23|_DFF_GG|I_T|B 0 _PG5_23|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_DFF_GG|I_6|B _PG5_23|_DFF_GG|Q1 _PG5_23|_DFF_GG|I_6|MID  2e-12
I_PG5_23|_DFF_GG|I_6|B 0 _PG5_23|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_DFF_GG|1|1 _PG5_23|_DFF_GG|A1 _PG5_23|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_GG|1|P _PG5_23|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG5_23|_DFF_GG|1|B _PG5_23|_DFF_GG|A1 _PG5_23|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_GG|1|RB _PG5_23|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_GG|23|1 _PG5_23|_DFF_GG|A2 _PG5_23|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_GG|23|B _PG5_23|_DFF_GG|A2 _PG5_23|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_GG|23|RB _PG5_23|_DFF_GG|23|MID_SHUNT _PG5_23|_DFF_GG|A3  2.1704737578552e-12
B_PG5_23|_DFF_GG|3|1 _PG5_23|_DFF_GG|A3 _PG5_23|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_GG|3|P _PG5_23|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG5_23|_DFF_GG|3|B _PG5_23|_DFF_GG|A3 _PG5_23|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_GG|3|RB _PG5_23|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_GG|4|1 _PG5_23|_DFF_GG|A4 _PG5_23|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_GG|4|P _PG5_23|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG5_23|_DFF_GG|4|B _PG5_23|_DFF_GG|A4 _PG5_23|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_GG|4|RB _PG5_23|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_GG|T|1 _PG5_23|_DFF_GG|T1 _PG5_23|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_GG|T|P _PG5_23|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG5_23|_DFF_GG|T|B _PG5_23|_DFF_GG|T1 _PG5_23|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_GG|T|RB _PG5_23|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_DFF_GG|45|1 _PG5_23|_DFF_GG|T2 _PG5_23|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG5_23|_DFF_GG|45|B _PG5_23|_DFF_GG|T2 _PG5_23|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG5_23|_DFF_GG|45|RB _PG5_23|_DFF_GG|45|MID_SHUNT _PG5_23|_DFF_GG|A4  2.1704737578552e-12
B_PG5_23|_DFF_GG|6|1 _PG5_23|_DFF_GG|Q1 _PG5_23|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_DFF_GG|6|P _PG5_23|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG5_23|_DFF_GG|6|B _PG5_23|_DFF_GG|Q1 _PG5_23|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG5_23|_DFF_GG|6|RB _PG5_23|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_AND_G|I_A1|B _PG5_23|_AND_G|A1 _PG5_23|_AND_G|I_A1|MID  2e-12
I_PG5_23|_AND_G|I_A1|B 0 _PG5_23|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_AND_G|I_B1|B _PG5_23|_AND_G|B1 _PG5_23|_AND_G|I_B1|MID  2e-12
I_PG5_23|_AND_G|I_B1|B 0 _PG5_23|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_AND_G|I_Q3|B _PG5_23|_AND_G|Q3 _PG5_23|_AND_G|I_Q3|MID  2e-12
I_PG5_23|_AND_G|I_Q3|B 0 _PG5_23|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG5_23|_AND_G|I_Q2|B _PG5_23|_AND_G|Q2 _PG5_23|_AND_G|I_Q2|MID  2e-12
I_PG5_23|_AND_G|I_Q2|B 0 _PG5_23|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_AND_G|I_Q1|B _PG5_23|_AND_G|Q1 _PG5_23|_AND_G|I_Q1|MID  2e-12
I_PG5_23|_AND_G|I_Q1|B 0 _PG5_23|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_AND_G|A1|1 _PG5_23|_AND_G|A1 _PG5_23|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_G|A1|P _PG5_23|_AND_G|A1|MID_SERIES 0  2e-13
R_PG5_23|_AND_G|A1|B _PG5_23|_AND_G|A1 _PG5_23|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG5_23|_AND_G|A1|RB _PG5_23|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_G|A2|1 _PG5_23|_AND_G|A2 _PG5_23|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_G|A2|P _PG5_23|_AND_G|A2|MID_SERIES 0  2e-13
R_PG5_23|_AND_G|A2|B _PG5_23|_AND_G|A2 _PG5_23|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG5_23|_AND_G|A2|RB _PG5_23|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_G|A12|1 _PG5_23|_AND_G|A2 _PG5_23|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_AND_G|A12|B _PG5_23|_AND_G|A2 _PG5_23|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG5_23|_AND_G|A12|RB _PG5_23|_AND_G|A12|MID_SHUNT _PG5_23|_AND_G|A3  2.1704737578552e-12
B_PG5_23|_AND_G|B1|1 _PG5_23|_AND_G|B1 _PG5_23|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_G|B1|P _PG5_23|_AND_G|B1|MID_SERIES 0  2e-13
R_PG5_23|_AND_G|B1|B _PG5_23|_AND_G|B1 _PG5_23|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG5_23|_AND_G|B1|RB _PG5_23|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_G|B2|1 _PG5_23|_AND_G|B2 _PG5_23|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_G|B2|P _PG5_23|_AND_G|B2|MID_SERIES 0  2e-13
R_PG5_23|_AND_G|B2|B _PG5_23|_AND_G|B2 _PG5_23|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG5_23|_AND_G|B2|RB _PG5_23|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_G|B12|1 _PG5_23|_AND_G|B2 _PG5_23|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG5_23|_AND_G|B12|B _PG5_23|_AND_G|B2 _PG5_23|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG5_23|_AND_G|B12|RB _PG5_23|_AND_G|B12|MID_SHUNT _PG5_23|_AND_G|B3  2.1704737578552e-12
B_PG5_23|_AND_G|Q2|1 _PG5_23|_AND_G|Q2 _PG5_23|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_G|Q2|P _PG5_23|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG5_23|_AND_G|Q2|B _PG5_23|_AND_G|Q2 _PG5_23|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG5_23|_AND_G|Q2|RB _PG5_23|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_G|Q1|1 _PG5_23|_AND_G|Q1 _PG5_23|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_G|Q1|P _PG5_23|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG5_23|_AND_G|Q1|B _PG5_23|_AND_G|Q1 _PG5_23|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG5_23|_AND_G|Q1|RB _PG5_23|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG5_23|_AND_P|I_A1|B _PG5_23|_AND_P|A1 _PG5_23|_AND_P|I_A1|MID  2e-12
I_PG5_23|_AND_P|I_A1|B 0 _PG5_23|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_AND_P|I_B1|B _PG5_23|_AND_P|B1 _PG5_23|_AND_P|I_B1|MID  2e-12
I_PG5_23|_AND_P|I_B1|B 0 _PG5_23|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_AND_P|I_Q3|B _PG5_23|_AND_P|Q3 _PG5_23|_AND_P|I_Q3|MID  2e-12
I_PG5_23|_AND_P|I_Q3|B 0 _PG5_23|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG5_23|_AND_P|I_Q2|B _PG5_23|_AND_P|Q2 _PG5_23|_AND_P|I_Q2|MID  2e-12
I_PG5_23|_AND_P|I_Q2|B 0 _PG5_23|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG5_23|_AND_P|I_Q1|B _PG5_23|_AND_P|Q1 _PG5_23|_AND_P|I_Q1|MID  2e-12
I_PG5_23|_AND_P|I_Q1|B 0 _PG5_23|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG5_23|_AND_P|A1|1 _PG5_23|_AND_P|A1 _PG5_23|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_P|A1|P _PG5_23|_AND_P|A1|MID_SERIES 0  2e-13
R_PG5_23|_AND_P|A1|B _PG5_23|_AND_P|A1 _PG5_23|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG5_23|_AND_P|A1|RB _PG5_23|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_P|A2|1 _PG5_23|_AND_P|A2 _PG5_23|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_P|A2|P _PG5_23|_AND_P|A2|MID_SERIES 0  2e-13
R_PG5_23|_AND_P|A2|B _PG5_23|_AND_P|A2 _PG5_23|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG5_23|_AND_P|A2|RB _PG5_23|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_P|A12|1 _PG5_23|_AND_P|A2 _PG5_23|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG5_23|_AND_P|A12|B _PG5_23|_AND_P|A2 _PG5_23|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG5_23|_AND_P|A12|RB _PG5_23|_AND_P|A12|MID_SHUNT _PG5_23|_AND_P|A3  2.1704737578552e-12
B_PG5_23|_AND_P|B1|1 _PG5_23|_AND_P|B1 _PG5_23|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_P|B1|P _PG5_23|_AND_P|B1|MID_SERIES 0  2e-13
R_PG5_23|_AND_P|B1|B _PG5_23|_AND_P|B1 _PG5_23|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG5_23|_AND_P|B1|RB _PG5_23|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_P|B2|1 _PG5_23|_AND_P|B2 _PG5_23|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_P|B2|P _PG5_23|_AND_P|B2|MID_SERIES 0  2e-13
R_PG5_23|_AND_P|B2|B _PG5_23|_AND_P|B2 _PG5_23|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG5_23|_AND_P|B2|RB _PG5_23|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_P|B12|1 _PG5_23|_AND_P|B2 _PG5_23|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG5_23|_AND_P|B12|B _PG5_23|_AND_P|B2 _PG5_23|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG5_23|_AND_P|B12|RB _PG5_23|_AND_P|B12|MID_SHUNT _PG5_23|_AND_P|B3  2.1704737578552e-12
B_PG5_23|_AND_P|Q2|1 _PG5_23|_AND_P|Q2 _PG5_23|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_P|Q2|P _PG5_23|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG5_23|_AND_P|Q2|B _PG5_23|_AND_P|Q2 _PG5_23|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG5_23|_AND_P|Q2|RB _PG5_23|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG5_23|_AND_P|Q1|1 _PG5_23|_AND_P|Q1 _PG5_23|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG5_23|_AND_P|Q1|P _PG5_23|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG5_23|_AND_P|Q1|B _PG5_23|_AND_P|Q1 _PG5_23|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG5_23|_AND_P|Q1|RB _PG5_23|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG6_23|P|I_1|B _PG6_23|P|A1 _PG6_23|P|I_1|MID  2e-12
I_PG6_23|P|I_1|B 0 _PG6_23|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_23|P|I_3|B _PG6_23|P|A3 _PG6_23|P|I_3|MID  2e-12
I_PG6_23|P|I_3|B 0 _PG6_23|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_23|P|I_T|B _PG6_23|P|T1 _PG6_23|P|I_T|MID  2e-12
I_PG6_23|P|I_T|B 0 _PG6_23|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_23|P|I_6|B _PG6_23|P|Q1 _PG6_23|P|I_6|MID  2e-12
I_PG6_23|P|I_6|B 0 _PG6_23|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_23|P|1|1 _PG6_23|P|A1 _PG6_23|P|1|MID_SERIES JJMIT AREA=2.5
L_PG6_23|P|1|P _PG6_23|P|1|MID_SERIES 0  2e-13
R_PG6_23|P|1|B _PG6_23|P|A1 _PG6_23|P|1|MID_SHUNT  2.7439617672
L_PG6_23|P|1|RB _PG6_23|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|P|23|1 _PG6_23|P|A2 _PG6_23|P|A3 JJMIT AREA=1.7857142857142858
R_PG6_23|P|23|B _PG6_23|P|A2 _PG6_23|P|23|MID_SHUNT  3.84154647408
L_PG6_23|P|23|RB _PG6_23|P|23|MID_SHUNT _PG6_23|P|A3  2.1704737578552e-12
B_PG6_23|P|3|1 _PG6_23|P|A3 _PG6_23|P|3|MID_SERIES JJMIT AREA=2.5
L_PG6_23|P|3|P _PG6_23|P|3|MID_SERIES 0  2e-13
R_PG6_23|P|3|B _PG6_23|P|A3 _PG6_23|P|3|MID_SHUNT  2.7439617672
L_PG6_23|P|3|RB _PG6_23|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|P|4|1 _PG6_23|P|A4 _PG6_23|P|4|MID_SERIES JJMIT AREA=2.5
L_PG6_23|P|4|P _PG6_23|P|4|MID_SERIES 0  2e-13
R_PG6_23|P|4|B _PG6_23|P|A4 _PG6_23|P|4|MID_SHUNT  2.7439617672
L_PG6_23|P|4|RB _PG6_23|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|P|T|1 _PG6_23|P|T1 _PG6_23|P|T|MID_SERIES JJMIT AREA=2.5
L_PG6_23|P|T|P _PG6_23|P|T|MID_SERIES 0  2e-13
R_PG6_23|P|T|B _PG6_23|P|T1 _PG6_23|P|T|MID_SHUNT  2.7439617672
L_PG6_23|P|T|RB _PG6_23|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|P|45|1 _PG6_23|P|T2 _PG6_23|P|A4 JJMIT AREA=1.7857142857142858
R_PG6_23|P|45|B _PG6_23|P|T2 _PG6_23|P|45|MID_SHUNT  3.84154647408
L_PG6_23|P|45|RB _PG6_23|P|45|MID_SHUNT _PG6_23|P|A4  2.1704737578552e-12
B_PG6_23|P|6|1 _PG6_23|P|Q1 _PG6_23|P|6|MID_SERIES JJMIT AREA=2.5
L_PG6_23|P|6|P _PG6_23|P|6|MID_SERIES 0  2e-13
R_PG6_23|P|6|B _PG6_23|P|Q1 _PG6_23|P|6|MID_SHUNT  2.7439617672
L_PG6_23|P|6|RB _PG6_23|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_23|G|I_1|B _PG6_23|G|A1 _PG6_23|G|I_1|MID  2e-12
I_PG6_23|G|I_1|B 0 _PG6_23|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_23|G|I_3|B _PG6_23|G|A3 _PG6_23|G|I_3|MID  2e-12
I_PG6_23|G|I_3|B 0 _PG6_23|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_23|G|I_T|B _PG6_23|G|T1 _PG6_23|G|I_T|MID  2e-12
I_PG6_23|G|I_T|B 0 _PG6_23|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_23|G|I_6|B _PG6_23|G|Q1 _PG6_23|G|I_6|MID  2e-12
I_PG6_23|G|I_6|B 0 _PG6_23|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_23|G|1|1 _PG6_23|G|A1 _PG6_23|G|1|MID_SERIES JJMIT AREA=2.5
L_PG6_23|G|1|P _PG6_23|G|1|MID_SERIES 0  2e-13
R_PG6_23|G|1|B _PG6_23|G|A1 _PG6_23|G|1|MID_SHUNT  2.7439617672
L_PG6_23|G|1|RB _PG6_23|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|G|23|1 _PG6_23|G|A2 _PG6_23|G|A3 JJMIT AREA=1.7857142857142858
R_PG6_23|G|23|B _PG6_23|G|A2 _PG6_23|G|23|MID_SHUNT  3.84154647408
L_PG6_23|G|23|RB _PG6_23|G|23|MID_SHUNT _PG6_23|G|A3  2.1704737578552e-12
B_PG6_23|G|3|1 _PG6_23|G|A3 _PG6_23|G|3|MID_SERIES JJMIT AREA=2.5
L_PG6_23|G|3|P _PG6_23|G|3|MID_SERIES 0  2e-13
R_PG6_23|G|3|B _PG6_23|G|A3 _PG6_23|G|3|MID_SHUNT  2.7439617672
L_PG6_23|G|3|RB _PG6_23|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|G|4|1 _PG6_23|G|A4 _PG6_23|G|4|MID_SERIES JJMIT AREA=2.5
L_PG6_23|G|4|P _PG6_23|G|4|MID_SERIES 0  2e-13
R_PG6_23|G|4|B _PG6_23|G|A4 _PG6_23|G|4|MID_SHUNT  2.7439617672
L_PG6_23|G|4|RB _PG6_23|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|G|T|1 _PG6_23|G|T1 _PG6_23|G|T|MID_SERIES JJMIT AREA=2.5
L_PG6_23|G|T|P _PG6_23|G|T|MID_SERIES 0  2e-13
R_PG6_23|G|T|B _PG6_23|G|T1 _PG6_23|G|T|MID_SHUNT  2.7439617672
L_PG6_23|G|T|RB _PG6_23|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_23|G|45|1 _PG6_23|G|T2 _PG6_23|G|A4 JJMIT AREA=1.7857142857142858
R_PG6_23|G|45|B _PG6_23|G|T2 _PG6_23|G|45|MID_SHUNT  3.84154647408
L_PG6_23|G|45|RB _PG6_23|G|45|MID_SHUNT _PG6_23|G|A4  2.1704737578552e-12
B_PG6_23|G|6|1 _PG6_23|G|Q1 _PG6_23|G|6|MID_SERIES JJMIT AREA=2.5
L_PG6_23|G|6|P _PG6_23|G|6|MID_SERIES 0  2e-13
R_PG6_23|G|6|B _PG6_23|G|Q1 _PG6_23|G|6|MID_SHUNT  2.7439617672
L_PG6_23|G|6|RB _PG6_23|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_SPL_G1|I_D1|B _PG7_23|_SPL_G1|D1 _PG7_23|_SPL_G1|I_D1|MID  2e-12
I_PG7_23|_SPL_G1|I_D1|B 0 _PG7_23|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_23|_SPL_G1|I_D2|B _PG7_23|_SPL_G1|D2 _PG7_23|_SPL_G1|I_D2|MID  2e-12
I_PG7_23|_SPL_G1|I_D2|B 0 _PG7_23|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG7_23|_SPL_G1|I_Q1|B _PG7_23|_SPL_G1|QA1 _PG7_23|_SPL_G1|I_Q1|MID  2e-12
I_PG7_23|_SPL_G1|I_Q1|B 0 _PG7_23|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_23|_SPL_G1|I_Q2|B _PG7_23|_SPL_G1|QB1 _PG7_23|_SPL_G1|I_Q2|MID  2e-12
I_PG7_23|_SPL_G1|I_Q2|B 0 _PG7_23|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG7_23|_SPL_G1|1|1 _PG7_23|_SPL_G1|D1 _PG7_23|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_G1|1|P _PG7_23|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG7_23|_SPL_G1|1|B _PG7_23|_SPL_G1|D1 _PG7_23|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_G1|1|RB _PG7_23|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_SPL_G1|2|1 _PG7_23|_SPL_G1|D2 _PG7_23|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_G1|2|P _PG7_23|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG7_23|_SPL_G1|2|B _PG7_23|_SPL_G1|D2 _PG7_23|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_G1|2|RB _PG7_23|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_SPL_G1|A|1 _PG7_23|_SPL_G1|QA1 _PG7_23|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_G1|A|P _PG7_23|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG7_23|_SPL_G1|A|B _PG7_23|_SPL_G1|QA1 _PG7_23|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_G1|A|RB _PG7_23|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_SPL_G1|B|1 _PG7_23|_SPL_G1|QB1 _PG7_23|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_G1|B|P _PG7_23|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG7_23|_SPL_G1|B|B _PG7_23|_SPL_G1|QB1 _PG7_23|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_G1|B|RB _PG7_23|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_SPL_P1|I_D1|B _PG7_23|_SPL_P1|D1 _PG7_23|_SPL_P1|I_D1|MID  2e-12
I_PG7_23|_SPL_P1|I_D1|B 0 _PG7_23|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_23|_SPL_P1|I_D2|B _PG7_23|_SPL_P1|D2 _PG7_23|_SPL_P1|I_D2|MID  2e-12
I_PG7_23|_SPL_P1|I_D2|B 0 _PG7_23|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG7_23|_SPL_P1|I_Q1|B _PG7_23|_SPL_P1|QA1 _PG7_23|_SPL_P1|I_Q1|MID  2e-12
I_PG7_23|_SPL_P1|I_Q1|B 0 _PG7_23|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG7_23|_SPL_P1|I_Q2|B _PG7_23|_SPL_P1|QB1 _PG7_23|_SPL_P1|I_Q2|MID  2e-12
I_PG7_23|_SPL_P1|I_Q2|B 0 _PG7_23|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG7_23|_SPL_P1|1|1 _PG7_23|_SPL_P1|D1 _PG7_23|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_P1|1|P _PG7_23|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG7_23|_SPL_P1|1|B _PG7_23|_SPL_P1|D1 _PG7_23|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_P1|1|RB _PG7_23|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_SPL_P1|2|1 _PG7_23|_SPL_P1|D2 _PG7_23|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_P1|2|P _PG7_23|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG7_23|_SPL_P1|2|B _PG7_23|_SPL_P1|D2 _PG7_23|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_P1|2|RB _PG7_23|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_SPL_P1|A|1 _PG7_23|_SPL_P1|QA1 _PG7_23|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_P1|A|P _PG7_23|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG7_23|_SPL_P1|A|B _PG7_23|_SPL_P1|QA1 _PG7_23|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_P1|A|RB _PG7_23|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_SPL_P1|B|1 _PG7_23|_SPL_P1|QB1 _PG7_23|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_SPL_P1|B|P _PG7_23|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG7_23|_SPL_P1|B|B _PG7_23|_SPL_P1|QB1 _PG7_23|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG7_23|_SPL_P1|B|RB _PG7_23|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_PG|I_A1|B _PG7_23|_PG|A1 _PG7_23|_PG|I_A1|MID  2e-12
I_PG7_23|_PG|I_A1|B 0 _PG7_23|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_PG|I_B1|B _PG7_23|_PG|B1 _PG7_23|_PG|I_B1|MID  2e-12
I_PG7_23|_PG|I_B1|B 0 _PG7_23|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_PG|I_Q3|B _PG7_23|_PG|Q3 _PG7_23|_PG|I_Q3|MID  2e-12
I_PG7_23|_PG|I_Q3|B 0 _PG7_23|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_23|_PG|I_Q2|B _PG7_23|_PG|Q2 _PG7_23|_PG|I_Q2|MID  2e-12
I_PG7_23|_PG|I_Q2|B 0 _PG7_23|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_PG|I_Q1|B _PG7_23|_PG|Q1 _PG7_23|_PG|I_Q1|MID  2e-12
I_PG7_23|_PG|I_Q1|B 0 _PG7_23|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_PG|A1|1 _PG7_23|_PG|A1 _PG7_23|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_PG|A1|P _PG7_23|_PG|A1|MID_SERIES 0  2e-13
R_PG7_23|_PG|A1|B _PG7_23|_PG|A1 _PG7_23|_PG|A1|MID_SHUNT  2.7439617672
L_PG7_23|_PG|A1|RB _PG7_23|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_PG|A2|1 _PG7_23|_PG|A2 _PG7_23|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_PG|A2|P _PG7_23|_PG|A2|MID_SERIES 0  2e-13
R_PG7_23|_PG|A2|B _PG7_23|_PG|A2 _PG7_23|_PG|A2|MID_SHUNT  2.7439617672
L_PG7_23|_PG|A2|RB _PG7_23|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_PG|A12|1 _PG7_23|_PG|A2 _PG7_23|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_PG|A12|B _PG7_23|_PG|A2 _PG7_23|_PG|A12|MID_SHUNT  3.84154647408
L_PG7_23|_PG|A12|RB _PG7_23|_PG|A12|MID_SHUNT _PG7_23|_PG|A3  2.1704737578552e-12
B_PG7_23|_PG|B1|1 _PG7_23|_PG|B1 _PG7_23|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_PG|B1|P _PG7_23|_PG|B1|MID_SERIES 0  2e-13
R_PG7_23|_PG|B1|B _PG7_23|_PG|B1 _PG7_23|_PG|B1|MID_SHUNT  2.7439617672
L_PG7_23|_PG|B1|RB _PG7_23|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_PG|B2|1 _PG7_23|_PG|B2 _PG7_23|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_PG|B2|P _PG7_23|_PG|B2|MID_SERIES 0  2e-13
R_PG7_23|_PG|B2|B _PG7_23|_PG|B2 _PG7_23|_PG|B2|MID_SHUNT  2.7439617672
L_PG7_23|_PG|B2|RB _PG7_23|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_PG|B12|1 _PG7_23|_PG|B2 _PG7_23|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG7_23|_PG|B12|B _PG7_23|_PG|B2 _PG7_23|_PG|B12|MID_SHUNT  3.84154647408
L_PG7_23|_PG|B12|RB _PG7_23|_PG|B12|MID_SHUNT _PG7_23|_PG|B3  2.1704737578552e-12
B_PG7_23|_PG|Q2|1 _PG7_23|_PG|Q2 _PG7_23|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_PG|Q2|P _PG7_23|_PG|Q2|MID_SERIES 0  2e-13
R_PG7_23|_PG|Q2|B _PG7_23|_PG|Q2 _PG7_23|_PG|Q2|MID_SHUNT  2.7439617672
L_PG7_23|_PG|Q2|RB _PG7_23|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_PG|Q1|1 _PG7_23|_PG|Q1 _PG7_23|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_PG|Q1|P _PG7_23|_PG|Q1|MID_SERIES 0  2e-13
R_PG7_23|_PG|Q1|B _PG7_23|_PG|Q1 _PG7_23|_PG|Q1|MID_SHUNT  2.7439617672
L_PG7_23|_PG|Q1|RB _PG7_23|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_GG|I_A1|B _PG7_23|_GG|A1 _PG7_23|_GG|I_A1|MID  2e-12
I_PG7_23|_GG|I_A1|B 0 _PG7_23|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_GG|I_B1|B _PG7_23|_GG|B1 _PG7_23|_GG|I_B1|MID  2e-12
I_PG7_23|_GG|I_B1|B 0 _PG7_23|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_GG|I_Q3|B _PG7_23|_GG|Q3 _PG7_23|_GG|I_Q3|MID  2e-12
I_PG7_23|_GG|I_Q3|B 0 _PG7_23|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_23|_GG|I_Q2|B _PG7_23|_GG|Q2 _PG7_23|_GG|I_Q2|MID  2e-12
I_PG7_23|_GG|I_Q2|B 0 _PG7_23|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_GG|I_Q1|B _PG7_23|_GG|Q1 _PG7_23|_GG|I_Q1|MID  2e-12
I_PG7_23|_GG|I_Q1|B 0 _PG7_23|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_GG|A1|1 _PG7_23|_GG|A1 _PG7_23|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_GG|A1|P _PG7_23|_GG|A1|MID_SERIES 0  2e-13
R_PG7_23|_GG|A1|B _PG7_23|_GG|A1 _PG7_23|_GG|A1|MID_SHUNT  2.7439617672
L_PG7_23|_GG|A1|RB _PG7_23|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_GG|A2|1 _PG7_23|_GG|A2 _PG7_23|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_GG|A2|P _PG7_23|_GG|A2|MID_SERIES 0  2e-13
R_PG7_23|_GG|A2|B _PG7_23|_GG|A2 _PG7_23|_GG|A2|MID_SHUNT  2.7439617672
L_PG7_23|_GG|A2|RB _PG7_23|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_GG|A12|1 _PG7_23|_GG|A2 _PG7_23|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_GG|A12|B _PG7_23|_GG|A2 _PG7_23|_GG|A12|MID_SHUNT  3.84154647408
L_PG7_23|_GG|A12|RB _PG7_23|_GG|A12|MID_SHUNT _PG7_23|_GG|A3  2.1704737578552e-12
B_PG7_23|_GG|B1|1 _PG7_23|_GG|B1 _PG7_23|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_GG|B1|P _PG7_23|_GG|B1|MID_SERIES 0  2e-13
R_PG7_23|_GG|B1|B _PG7_23|_GG|B1 _PG7_23|_GG|B1|MID_SHUNT  2.7439617672
L_PG7_23|_GG|B1|RB _PG7_23|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_GG|B2|1 _PG7_23|_GG|B2 _PG7_23|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_GG|B2|P _PG7_23|_GG|B2|MID_SERIES 0  2e-13
R_PG7_23|_GG|B2|B _PG7_23|_GG|B2 _PG7_23|_GG|B2|MID_SHUNT  2.7439617672
L_PG7_23|_GG|B2|RB _PG7_23|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_GG|B12|1 _PG7_23|_GG|B2 _PG7_23|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG7_23|_GG|B12|B _PG7_23|_GG|B2 _PG7_23|_GG|B12|MID_SHUNT  3.84154647408
L_PG7_23|_GG|B12|RB _PG7_23|_GG|B12|MID_SHUNT _PG7_23|_GG|B3  2.1704737578552e-12
B_PG7_23|_GG|Q2|1 _PG7_23|_GG|Q2 _PG7_23|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_GG|Q2|P _PG7_23|_GG|Q2|MID_SERIES 0  2e-13
R_PG7_23|_GG|Q2|B _PG7_23|_GG|Q2 _PG7_23|_GG|Q2|MID_SHUNT  2.7439617672
L_PG7_23|_GG|Q2|RB _PG7_23|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_GG|Q1|1 _PG7_23|_GG|Q1 _PG7_23|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_GG|Q1|P _PG7_23|_GG|Q1|MID_SERIES 0  2e-13
R_PG7_23|_GG|Q1|B _PG7_23|_GG|Q1 _PG7_23|_GG|Q1|MID_SHUNT  2.7439617672
L_PG7_23|_GG|Q1|RB _PG7_23|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_DFF_P0|I_1|B _PG7_23|_DFF_P0|A1 _PG7_23|_DFF_P0|I_1|MID  2e-12
I_PG7_23|_DFF_P0|I_1|B 0 _PG7_23|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_P0|I_3|B _PG7_23|_DFF_P0|A3 _PG7_23|_DFF_P0|I_3|MID  2e-12
I_PG7_23|_DFF_P0|I_3|B 0 _PG7_23|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_23|_DFF_P0|I_T|B _PG7_23|_DFF_P0|T1 _PG7_23|_DFF_P0|I_T|MID  2e-12
I_PG7_23|_DFF_P0|I_T|B 0 _PG7_23|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_P0|I_6|B _PG7_23|_DFF_P0|Q1 _PG7_23|_DFF_P0|I_6|MID  2e-12
I_PG7_23|_DFF_P0|I_6|B 0 _PG7_23|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_DFF_P0|1|1 _PG7_23|_DFF_P0|A1 _PG7_23|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P0|1|P _PG7_23|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P0|1|B _PG7_23|_DFF_P0|A1 _PG7_23|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P0|1|RB _PG7_23|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P0|23|1 _PG7_23|_DFF_P0|A2 _PG7_23|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_P0|23|B _PG7_23|_DFF_P0|A2 _PG7_23|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_P0|23|RB _PG7_23|_DFF_P0|23|MID_SHUNT _PG7_23|_DFF_P0|A3  2.1704737578552e-12
B_PG7_23|_DFF_P0|3|1 _PG7_23|_DFF_P0|A3 _PG7_23|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P0|3|P _PG7_23|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P0|3|B _PG7_23|_DFF_P0|A3 _PG7_23|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P0|3|RB _PG7_23|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P0|4|1 _PG7_23|_DFF_P0|A4 _PG7_23|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P0|4|P _PG7_23|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P0|4|B _PG7_23|_DFF_P0|A4 _PG7_23|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P0|4|RB _PG7_23|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P0|T|1 _PG7_23|_DFF_P0|T1 _PG7_23|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P0|T|P _PG7_23|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P0|T|B _PG7_23|_DFF_P0|T1 _PG7_23|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P0|T|RB _PG7_23|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P0|45|1 _PG7_23|_DFF_P0|T2 _PG7_23|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_P0|45|B _PG7_23|_DFF_P0|T2 _PG7_23|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_P0|45|RB _PG7_23|_DFF_P0|45|MID_SHUNT _PG7_23|_DFF_P0|A4  2.1704737578552e-12
B_PG7_23|_DFF_P0|6|1 _PG7_23|_DFF_P0|Q1 _PG7_23|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P0|6|P _PG7_23|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P0|6|B _PG7_23|_DFF_P0|Q1 _PG7_23|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P0|6|RB _PG7_23|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_DFF_P1|I_1|B _PG7_23|_DFF_P1|A1 _PG7_23|_DFF_P1|I_1|MID  2e-12
I_PG7_23|_DFF_P1|I_1|B 0 _PG7_23|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_P1|I_3|B _PG7_23|_DFF_P1|A3 _PG7_23|_DFF_P1|I_3|MID  2e-12
I_PG7_23|_DFF_P1|I_3|B 0 _PG7_23|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_23|_DFF_P1|I_T|B _PG7_23|_DFF_P1|T1 _PG7_23|_DFF_P1|I_T|MID  2e-12
I_PG7_23|_DFF_P1|I_T|B 0 _PG7_23|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_P1|I_6|B _PG7_23|_DFF_P1|Q1 _PG7_23|_DFF_P1|I_6|MID  2e-12
I_PG7_23|_DFF_P1|I_6|B 0 _PG7_23|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_DFF_P1|1|1 _PG7_23|_DFF_P1|A1 _PG7_23|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P1|1|P _PG7_23|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P1|1|B _PG7_23|_DFF_P1|A1 _PG7_23|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P1|1|RB _PG7_23|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P1|23|1 _PG7_23|_DFF_P1|A2 _PG7_23|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_P1|23|B _PG7_23|_DFF_P1|A2 _PG7_23|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_P1|23|RB _PG7_23|_DFF_P1|23|MID_SHUNT _PG7_23|_DFF_P1|A3  2.1704737578552e-12
B_PG7_23|_DFF_P1|3|1 _PG7_23|_DFF_P1|A3 _PG7_23|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P1|3|P _PG7_23|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P1|3|B _PG7_23|_DFF_P1|A3 _PG7_23|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P1|3|RB _PG7_23|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P1|4|1 _PG7_23|_DFF_P1|A4 _PG7_23|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P1|4|P _PG7_23|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P1|4|B _PG7_23|_DFF_P1|A4 _PG7_23|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P1|4|RB _PG7_23|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P1|T|1 _PG7_23|_DFF_P1|T1 _PG7_23|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P1|T|P _PG7_23|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P1|T|B _PG7_23|_DFF_P1|T1 _PG7_23|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P1|T|RB _PG7_23|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_P1|45|1 _PG7_23|_DFF_P1|T2 _PG7_23|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_P1|45|B _PG7_23|_DFF_P1|T2 _PG7_23|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_P1|45|RB _PG7_23|_DFF_P1|45|MID_SHUNT _PG7_23|_DFF_P1|A4  2.1704737578552e-12
B_PG7_23|_DFF_P1|6|1 _PG7_23|_DFF_P1|Q1 _PG7_23|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_P1|6|P _PG7_23|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG7_23|_DFF_P1|6|B _PG7_23|_DFF_P1|Q1 _PG7_23|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_P1|6|RB _PG7_23|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_DFF_PG|I_1|B _PG7_23|_DFF_PG|A1 _PG7_23|_DFF_PG|I_1|MID  2e-12
I_PG7_23|_DFF_PG|I_1|B 0 _PG7_23|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_PG|I_3|B _PG7_23|_DFF_PG|A3 _PG7_23|_DFF_PG|I_3|MID  2e-12
I_PG7_23|_DFF_PG|I_3|B 0 _PG7_23|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_23|_DFF_PG|I_T|B _PG7_23|_DFF_PG|T1 _PG7_23|_DFF_PG|I_T|MID  2e-12
I_PG7_23|_DFF_PG|I_T|B 0 _PG7_23|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_PG|I_6|B _PG7_23|_DFF_PG|Q1 _PG7_23|_DFF_PG|I_6|MID  2e-12
I_PG7_23|_DFF_PG|I_6|B 0 _PG7_23|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_DFF_PG|1|1 _PG7_23|_DFF_PG|A1 _PG7_23|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_PG|1|P _PG7_23|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG7_23|_DFF_PG|1|B _PG7_23|_DFF_PG|A1 _PG7_23|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_PG|1|RB _PG7_23|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_PG|23|1 _PG7_23|_DFF_PG|A2 _PG7_23|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_PG|23|B _PG7_23|_DFF_PG|A2 _PG7_23|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_PG|23|RB _PG7_23|_DFF_PG|23|MID_SHUNT _PG7_23|_DFF_PG|A3  2.1704737578552e-12
B_PG7_23|_DFF_PG|3|1 _PG7_23|_DFF_PG|A3 _PG7_23|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_PG|3|P _PG7_23|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG7_23|_DFF_PG|3|B _PG7_23|_DFF_PG|A3 _PG7_23|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_PG|3|RB _PG7_23|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_PG|4|1 _PG7_23|_DFF_PG|A4 _PG7_23|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_PG|4|P _PG7_23|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG7_23|_DFF_PG|4|B _PG7_23|_DFF_PG|A4 _PG7_23|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_PG|4|RB _PG7_23|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_PG|T|1 _PG7_23|_DFF_PG|T1 _PG7_23|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_PG|T|P _PG7_23|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG7_23|_DFF_PG|T|B _PG7_23|_DFF_PG|T1 _PG7_23|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_PG|T|RB _PG7_23|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_PG|45|1 _PG7_23|_DFF_PG|T2 _PG7_23|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_PG|45|B _PG7_23|_DFF_PG|T2 _PG7_23|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_PG|45|RB _PG7_23|_DFF_PG|45|MID_SHUNT _PG7_23|_DFF_PG|A4  2.1704737578552e-12
B_PG7_23|_DFF_PG|6|1 _PG7_23|_DFF_PG|Q1 _PG7_23|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_PG|6|P _PG7_23|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG7_23|_DFF_PG|6|B _PG7_23|_DFF_PG|Q1 _PG7_23|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_PG|6|RB _PG7_23|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_DFF_GG|I_1|B _PG7_23|_DFF_GG|A1 _PG7_23|_DFF_GG|I_1|MID  2e-12
I_PG7_23|_DFF_GG|I_1|B 0 _PG7_23|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_GG|I_3|B _PG7_23|_DFF_GG|A3 _PG7_23|_DFF_GG|I_3|MID  2e-12
I_PG7_23|_DFF_GG|I_3|B 0 _PG7_23|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG7_23|_DFF_GG|I_T|B _PG7_23|_DFF_GG|T1 _PG7_23|_DFF_GG|I_T|MID  2e-12
I_PG7_23|_DFF_GG|I_T|B 0 _PG7_23|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_DFF_GG|I_6|B _PG7_23|_DFF_GG|Q1 _PG7_23|_DFF_GG|I_6|MID  2e-12
I_PG7_23|_DFF_GG|I_6|B 0 _PG7_23|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_DFF_GG|1|1 _PG7_23|_DFF_GG|A1 _PG7_23|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_GG|1|P _PG7_23|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG7_23|_DFF_GG|1|B _PG7_23|_DFF_GG|A1 _PG7_23|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_GG|1|RB _PG7_23|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_GG|23|1 _PG7_23|_DFF_GG|A2 _PG7_23|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_GG|23|B _PG7_23|_DFF_GG|A2 _PG7_23|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_GG|23|RB _PG7_23|_DFF_GG|23|MID_SHUNT _PG7_23|_DFF_GG|A3  2.1704737578552e-12
B_PG7_23|_DFF_GG|3|1 _PG7_23|_DFF_GG|A3 _PG7_23|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_GG|3|P _PG7_23|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG7_23|_DFF_GG|3|B _PG7_23|_DFF_GG|A3 _PG7_23|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_GG|3|RB _PG7_23|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_GG|4|1 _PG7_23|_DFF_GG|A4 _PG7_23|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_GG|4|P _PG7_23|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG7_23|_DFF_GG|4|B _PG7_23|_DFF_GG|A4 _PG7_23|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_GG|4|RB _PG7_23|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_GG|T|1 _PG7_23|_DFF_GG|T1 _PG7_23|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_GG|T|P _PG7_23|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG7_23|_DFF_GG|T|B _PG7_23|_DFF_GG|T1 _PG7_23|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_GG|T|RB _PG7_23|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_DFF_GG|45|1 _PG7_23|_DFF_GG|T2 _PG7_23|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG7_23|_DFF_GG|45|B _PG7_23|_DFF_GG|T2 _PG7_23|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG7_23|_DFF_GG|45|RB _PG7_23|_DFF_GG|45|MID_SHUNT _PG7_23|_DFF_GG|A4  2.1704737578552e-12
B_PG7_23|_DFF_GG|6|1 _PG7_23|_DFF_GG|Q1 _PG7_23|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_DFF_GG|6|P _PG7_23|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG7_23|_DFF_GG|6|B _PG7_23|_DFF_GG|Q1 _PG7_23|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG7_23|_DFF_GG|6|RB _PG7_23|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_AND_G|I_A1|B _PG7_23|_AND_G|A1 _PG7_23|_AND_G|I_A1|MID  2e-12
I_PG7_23|_AND_G|I_A1|B 0 _PG7_23|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_AND_G|I_B1|B _PG7_23|_AND_G|B1 _PG7_23|_AND_G|I_B1|MID  2e-12
I_PG7_23|_AND_G|I_B1|B 0 _PG7_23|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_AND_G|I_Q3|B _PG7_23|_AND_G|Q3 _PG7_23|_AND_G|I_Q3|MID  2e-12
I_PG7_23|_AND_G|I_Q3|B 0 _PG7_23|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG7_23|_AND_G|I_Q2|B _PG7_23|_AND_G|Q2 _PG7_23|_AND_G|I_Q2|MID  2e-12
I_PG7_23|_AND_G|I_Q2|B 0 _PG7_23|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_AND_G|I_Q1|B _PG7_23|_AND_G|Q1 _PG7_23|_AND_G|I_Q1|MID  2e-12
I_PG7_23|_AND_G|I_Q1|B 0 _PG7_23|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_AND_G|A1|1 _PG7_23|_AND_G|A1 _PG7_23|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_G|A1|P _PG7_23|_AND_G|A1|MID_SERIES 0  2e-13
R_PG7_23|_AND_G|A1|B _PG7_23|_AND_G|A1 _PG7_23|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG7_23|_AND_G|A1|RB _PG7_23|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_G|A2|1 _PG7_23|_AND_G|A2 _PG7_23|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_G|A2|P _PG7_23|_AND_G|A2|MID_SERIES 0  2e-13
R_PG7_23|_AND_G|A2|B _PG7_23|_AND_G|A2 _PG7_23|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG7_23|_AND_G|A2|RB _PG7_23|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_G|A12|1 _PG7_23|_AND_G|A2 _PG7_23|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_AND_G|A12|B _PG7_23|_AND_G|A2 _PG7_23|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG7_23|_AND_G|A12|RB _PG7_23|_AND_G|A12|MID_SHUNT _PG7_23|_AND_G|A3  2.1704737578552e-12
B_PG7_23|_AND_G|B1|1 _PG7_23|_AND_G|B1 _PG7_23|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_G|B1|P _PG7_23|_AND_G|B1|MID_SERIES 0  2e-13
R_PG7_23|_AND_G|B1|B _PG7_23|_AND_G|B1 _PG7_23|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG7_23|_AND_G|B1|RB _PG7_23|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_G|B2|1 _PG7_23|_AND_G|B2 _PG7_23|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_G|B2|P _PG7_23|_AND_G|B2|MID_SERIES 0  2e-13
R_PG7_23|_AND_G|B2|B _PG7_23|_AND_G|B2 _PG7_23|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG7_23|_AND_G|B2|RB _PG7_23|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_G|B12|1 _PG7_23|_AND_G|B2 _PG7_23|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG7_23|_AND_G|B12|B _PG7_23|_AND_G|B2 _PG7_23|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG7_23|_AND_G|B12|RB _PG7_23|_AND_G|B12|MID_SHUNT _PG7_23|_AND_G|B3  2.1704737578552e-12
B_PG7_23|_AND_G|Q2|1 _PG7_23|_AND_G|Q2 _PG7_23|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_G|Q2|P _PG7_23|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG7_23|_AND_G|Q2|B _PG7_23|_AND_G|Q2 _PG7_23|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG7_23|_AND_G|Q2|RB _PG7_23|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_G|Q1|1 _PG7_23|_AND_G|Q1 _PG7_23|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_G|Q1|P _PG7_23|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG7_23|_AND_G|Q1|B _PG7_23|_AND_G|Q1 _PG7_23|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG7_23|_AND_G|Q1|RB _PG7_23|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG7_23|_AND_P|I_A1|B _PG7_23|_AND_P|A1 _PG7_23|_AND_P|I_A1|MID  2e-12
I_PG7_23|_AND_P|I_A1|B 0 _PG7_23|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_AND_P|I_B1|B _PG7_23|_AND_P|B1 _PG7_23|_AND_P|I_B1|MID  2e-12
I_PG7_23|_AND_P|I_B1|B 0 _PG7_23|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_AND_P|I_Q3|B _PG7_23|_AND_P|Q3 _PG7_23|_AND_P|I_Q3|MID  2e-12
I_PG7_23|_AND_P|I_Q3|B 0 _PG7_23|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG7_23|_AND_P|I_Q2|B _PG7_23|_AND_P|Q2 _PG7_23|_AND_P|I_Q2|MID  2e-12
I_PG7_23|_AND_P|I_Q2|B 0 _PG7_23|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG7_23|_AND_P|I_Q1|B _PG7_23|_AND_P|Q1 _PG7_23|_AND_P|I_Q1|MID  2e-12
I_PG7_23|_AND_P|I_Q1|B 0 _PG7_23|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG7_23|_AND_P|A1|1 _PG7_23|_AND_P|A1 _PG7_23|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_P|A1|P _PG7_23|_AND_P|A1|MID_SERIES 0  2e-13
R_PG7_23|_AND_P|A1|B _PG7_23|_AND_P|A1 _PG7_23|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG7_23|_AND_P|A1|RB _PG7_23|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_P|A2|1 _PG7_23|_AND_P|A2 _PG7_23|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_P|A2|P _PG7_23|_AND_P|A2|MID_SERIES 0  2e-13
R_PG7_23|_AND_P|A2|B _PG7_23|_AND_P|A2 _PG7_23|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG7_23|_AND_P|A2|RB _PG7_23|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_P|A12|1 _PG7_23|_AND_P|A2 _PG7_23|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG7_23|_AND_P|A12|B _PG7_23|_AND_P|A2 _PG7_23|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG7_23|_AND_P|A12|RB _PG7_23|_AND_P|A12|MID_SHUNT _PG7_23|_AND_P|A3  2.1704737578552e-12
B_PG7_23|_AND_P|B1|1 _PG7_23|_AND_P|B1 _PG7_23|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_P|B1|P _PG7_23|_AND_P|B1|MID_SERIES 0  2e-13
R_PG7_23|_AND_P|B1|B _PG7_23|_AND_P|B1 _PG7_23|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG7_23|_AND_P|B1|RB _PG7_23|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_P|B2|1 _PG7_23|_AND_P|B2 _PG7_23|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_P|B2|P _PG7_23|_AND_P|B2|MID_SERIES 0  2e-13
R_PG7_23|_AND_P|B2|B _PG7_23|_AND_P|B2 _PG7_23|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG7_23|_AND_P|B2|RB _PG7_23|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_P|B12|1 _PG7_23|_AND_P|B2 _PG7_23|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG7_23|_AND_P|B12|B _PG7_23|_AND_P|B2 _PG7_23|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG7_23|_AND_P|B12|RB _PG7_23|_AND_P|B12|MID_SHUNT _PG7_23|_AND_P|B3  2.1704737578552e-12
B_PG7_23|_AND_P|Q2|1 _PG7_23|_AND_P|Q2 _PG7_23|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_P|Q2|P _PG7_23|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG7_23|_AND_P|Q2|B _PG7_23|_AND_P|Q2 _PG7_23|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG7_23|_AND_P|Q2|RB _PG7_23|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG7_23|_AND_P|Q1|1 _PG7_23|_AND_P|Q1 _PG7_23|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG7_23|_AND_P|Q1|P _PG7_23|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG7_23|_AND_P|Q1|B _PG7_23|_AND_P|Q1 _PG7_23|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG7_23|_AND_P|Q1|RB _PG7_23|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PTL_G5_3|_SPL|I_D1|B _PTL_G5_3|_SPL|D1 _PTL_G5_3|_SPL|I_D1|MID  2e-12
I_PTL_G5_3|_SPL|I_D1|B 0 _PTL_G5_3|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G5_3|_SPL|I_D2|B _PTL_G5_3|_SPL|D2 _PTL_G5_3|_SPL|I_D2|MID  2e-12
I_PTL_G5_3|_SPL|I_D2|B 0 _PTL_G5_3|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G5_3|_SPL|I_Q1|B _PTL_G5_3|_SPL|QA1 _PTL_G5_3|_SPL|I_Q1|MID  2e-12
I_PTL_G5_3|_SPL|I_Q1|B 0 _PTL_G5_3|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G5_3|_SPL|I_Q2|B _PTL_G5_3|_SPL|QB1 _PTL_G5_3|_SPL|I_Q2|MID  2e-12
I_PTL_G5_3|_SPL|I_Q2|B 0 _PTL_G5_3|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G5_3|_SPL|1|1 _PTL_G5_3|_SPL|D1 _PTL_G5_3|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_3|_SPL|1|P _PTL_G5_3|_SPL|1|MID_SERIES 0  2e-13
R_PTL_G5_3|_SPL|1|B _PTL_G5_3|_SPL|D1 _PTL_G5_3|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_G5_3|_SPL|1|RB _PTL_G5_3|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G5_3|_SPL|2|1 _PTL_G5_3|_SPL|D2 _PTL_G5_3|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_3|_SPL|2|P _PTL_G5_3|_SPL|2|MID_SERIES 0  2e-13
R_PTL_G5_3|_SPL|2|B _PTL_G5_3|_SPL|D2 _PTL_G5_3|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_G5_3|_SPL|2|RB _PTL_G5_3|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G5_3|_SPL|A|1 _PTL_G5_3|_SPL|QA1 _PTL_G5_3|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_3|_SPL|A|P _PTL_G5_3|_SPL|A|MID_SERIES 0  2e-13
R_PTL_G5_3|_SPL|A|B _PTL_G5_3|_SPL|QA1 _PTL_G5_3|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_G5_3|_SPL|A|RB _PTL_G5_3|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G5_3|_SPL|B|1 _PTL_G5_3|_SPL|QB1 _PTL_G5_3|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G5_3|_SPL|B|P _PTL_G5_3|_SPL|B|MID_SERIES 0  2e-13
R_PTL_G5_3|_SPL|B|B _PTL_G5_3|_SPL|QB1 _PTL_G5_3|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_G5_3|_SPL|B|RB _PTL_G5_3|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_P6_3|_SPL|I_D1|B _PTL_P6_3|_SPL|D1 _PTL_P6_3|_SPL|I_D1|MID  2e-12
I_PTL_P6_3|_SPL|I_D1|B 0 _PTL_P6_3|_SPL|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P6_3|_SPL|I_D2|B _PTL_P6_3|_SPL|D2 _PTL_P6_3|_SPL|I_D2|MID  2e-12
I_PTL_P6_3|_SPL|I_D2|B 0 _PTL_P6_3|_SPL|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P6_3|_SPL|I_Q1|B _PTL_P6_3|_SPL|QA1 _PTL_P6_3|_SPL|I_Q1|MID  2e-12
I_PTL_P6_3|_SPL|I_Q1|B 0 _PTL_P6_3|_SPL|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P6_3|_SPL|I_Q2|B _PTL_P6_3|_SPL|QB1 _PTL_P6_3|_SPL|I_Q2|MID  2e-12
I_PTL_P6_3|_SPL|I_Q2|B 0 _PTL_P6_3|_SPL|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P6_3|_SPL|1|1 _PTL_P6_3|_SPL|D1 _PTL_P6_3|_SPL|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P6_3|_SPL|1|P _PTL_P6_3|_SPL|1|MID_SERIES 0  2e-13
R_PTL_P6_3|_SPL|1|B _PTL_P6_3|_SPL|D1 _PTL_P6_3|_SPL|1|MID_SHUNT  2.7439617672
L_PTL_P6_3|_SPL|1|RB _PTL_P6_3|_SPL|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P6_3|_SPL|2|1 _PTL_P6_3|_SPL|D2 _PTL_P6_3|_SPL|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P6_3|_SPL|2|P _PTL_P6_3|_SPL|2|MID_SERIES 0  2e-13
R_PTL_P6_3|_SPL|2|B _PTL_P6_3|_SPL|D2 _PTL_P6_3|_SPL|2|MID_SHUNT  2.7439617672
L_PTL_P6_3|_SPL|2|RB _PTL_P6_3|_SPL|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P6_3|_SPL|A|1 _PTL_P6_3|_SPL|QA1 _PTL_P6_3|_SPL|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P6_3|_SPL|A|P _PTL_P6_3|_SPL|A|MID_SERIES 0  2e-13
R_PTL_P6_3|_SPL|A|B _PTL_P6_3|_SPL|QA1 _PTL_P6_3|_SPL|A|MID_SHUNT  2.7439617672
L_PTL_P6_3|_SPL|A|RB _PTL_P6_3|_SPL|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P6_3|_SPL|B|1 _PTL_P6_3|_SPL|QB1 _PTL_P6_3|_SPL|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P6_3|_SPL|B|P _PTL_P6_3|_SPL|B|MID_SERIES 0  2e-13
R_PTL_P6_3|_SPL|B|B _PTL_P6_3|_SPL|QB1 _PTL_P6_3|_SPL|B|MID_SHUNT  2.7439617672
L_PTL_P6_3|_SPL|B|RB _PTL_P6_3|_SPL|B|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_SPL_G1|I_D1|B _PG6_34|_SPL_G1|D1 _PG6_34|_SPL_G1|I_D1|MID  2e-12
I_PG6_34|_SPL_G1|I_D1|B 0 _PG6_34|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG6_34|_SPL_G1|I_D2|B _PG6_34|_SPL_G1|D2 _PG6_34|_SPL_G1|I_D2|MID  2e-12
I_PG6_34|_SPL_G1|I_D2|B 0 _PG6_34|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG6_34|_SPL_G1|I_Q1|B _PG6_34|_SPL_G1|QA1 _PG6_34|_SPL_G1|I_Q1|MID  2e-12
I_PG6_34|_SPL_G1|I_Q1|B 0 _PG6_34|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG6_34|_SPL_G1|I_Q2|B _PG6_34|_SPL_G1|QB1 _PG6_34|_SPL_G1|I_Q2|MID  2e-12
I_PG6_34|_SPL_G1|I_Q2|B 0 _PG6_34|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG6_34|_SPL_G1|1|1 _PG6_34|_SPL_G1|D1 _PG6_34|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_G1|1|P _PG6_34|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG6_34|_SPL_G1|1|B _PG6_34|_SPL_G1|D1 _PG6_34|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_G1|1|RB _PG6_34|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_SPL_G1|2|1 _PG6_34|_SPL_G1|D2 _PG6_34|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_G1|2|P _PG6_34|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG6_34|_SPL_G1|2|B _PG6_34|_SPL_G1|D2 _PG6_34|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_G1|2|RB _PG6_34|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_SPL_G1|A|1 _PG6_34|_SPL_G1|QA1 _PG6_34|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_G1|A|P _PG6_34|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG6_34|_SPL_G1|A|B _PG6_34|_SPL_G1|QA1 _PG6_34|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_G1|A|RB _PG6_34|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_SPL_G1|B|1 _PG6_34|_SPL_G1|QB1 _PG6_34|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_G1|B|P _PG6_34|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG6_34|_SPL_G1|B|B _PG6_34|_SPL_G1|QB1 _PG6_34|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_G1|B|RB _PG6_34|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_SPL_P1|I_D1|B _PG6_34|_SPL_P1|D1 _PG6_34|_SPL_P1|I_D1|MID  2e-12
I_PG6_34|_SPL_P1|I_D1|B 0 _PG6_34|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG6_34|_SPL_P1|I_D2|B _PG6_34|_SPL_P1|D2 _PG6_34|_SPL_P1|I_D2|MID  2e-12
I_PG6_34|_SPL_P1|I_D2|B 0 _PG6_34|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG6_34|_SPL_P1|I_Q1|B _PG6_34|_SPL_P1|QA1 _PG6_34|_SPL_P1|I_Q1|MID  2e-12
I_PG6_34|_SPL_P1|I_Q1|B 0 _PG6_34|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG6_34|_SPL_P1|I_Q2|B _PG6_34|_SPL_P1|QB1 _PG6_34|_SPL_P1|I_Q2|MID  2e-12
I_PG6_34|_SPL_P1|I_Q2|B 0 _PG6_34|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG6_34|_SPL_P1|1|1 _PG6_34|_SPL_P1|D1 _PG6_34|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_P1|1|P _PG6_34|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG6_34|_SPL_P1|1|B _PG6_34|_SPL_P1|D1 _PG6_34|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_P1|1|RB _PG6_34|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_SPL_P1|2|1 _PG6_34|_SPL_P1|D2 _PG6_34|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_P1|2|P _PG6_34|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG6_34|_SPL_P1|2|B _PG6_34|_SPL_P1|D2 _PG6_34|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_P1|2|RB _PG6_34|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_SPL_P1|A|1 _PG6_34|_SPL_P1|QA1 _PG6_34|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_P1|A|P _PG6_34|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG6_34|_SPL_P1|A|B _PG6_34|_SPL_P1|QA1 _PG6_34|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_P1|A|RB _PG6_34|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_SPL_P1|B|1 _PG6_34|_SPL_P1|QB1 _PG6_34|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_SPL_P1|B|P _PG6_34|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG6_34|_SPL_P1|B|B _PG6_34|_SPL_P1|QB1 _PG6_34|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG6_34|_SPL_P1|B|RB _PG6_34|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_PG|I_A1|B _PG6_34|_PG|A1 _PG6_34|_PG|I_A1|MID  2e-12
I_PG6_34|_PG|I_A1|B 0 _PG6_34|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_PG|I_B1|B _PG6_34|_PG|B1 _PG6_34|_PG|I_B1|MID  2e-12
I_PG6_34|_PG|I_B1|B 0 _PG6_34|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_PG|I_Q3|B _PG6_34|_PG|Q3 _PG6_34|_PG|I_Q3|MID  2e-12
I_PG6_34|_PG|I_Q3|B 0 _PG6_34|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_34|_PG|I_Q2|B _PG6_34|_PG|Q2 _PG6_34|_PG|I_Q2|MID  2e-12
I_PG6_34|_PG|I_Q2|B 0 _PG6_34|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_PG|I_Q1|B _PG6_34|_PG|Q1 _PG6_34|_PG|I_Q1|MID  2e-12
I_PG6_34|_PG|I_Q1|B 0 _PG6_34|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_PG|A1|1 _PG6_34|_PG|A1 _PG6_34|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_PG|A1|P _PG6_34|_PG|A1|MID_SERIES 0  2e-13
R_PG6_34|_PG|A1|B _PG6_34|_PG|A1 _PG6_34|_PG|A1|MID_SHUNT  2.7439617672
L_PG6_34|_PG|A1|RB _PG6_34|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_PG|A2|1 _PG6_34|_PG|A2 _PG6_34|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_PG|A2|P _PG6_34|_PG|A2|MID_SERIES 0  2e-13
R_PG6_34|_PG|A2|B _PG6_34|_PG|A2 _PG6_34|_PG|A2|MID_SHUNT  2.7439617672
L_PG6_34|_PG|A2|RB _PG6_34|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_PG|A12|1 _PG6_34|_PG|A2 _PG6_34|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_PG|A12|B _PG6_34|_PG|A2 _PG6_34|_PG|A12|MID_SHUNT  3.84154647408
L_PG6_34|_PG|A12|RB _PG6_34|_PG|A12|MID_SHUNT _PG6_34|_PG|A3  2.1704737578552e-12
B_PG6_34|_PG|B1|1 _PG6_34|_PG|B1 _PG6_34|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_PG|B1|P _PG6_34|_PG|B1|MID_SERIES 0  2e-13
R_PG6_34|_PG|B1|B _PG6_34|_PG|B1 _PG6_34|_PG|B1|MID_SHUNT  2.7439617672
L_PG6_34|_PG|B1|RB _PG6_34|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_PG|B2|1 _PG6_34|_PG|B2 _PG6_34|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_PG|B2|P _PG6_34|_PG|B2|MID_SERIES 0  2e-13
R_PG6_34|_PG|B2|B _PG6_34|_PG|B2 _PG6_34|_PG|B2|MID_SHUNT  2.7439617672
L_PG6_34|_PG|B2|RB _PG6_34|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_PG|B12|1 _PG6_34|_PG|B2 _PG6_34|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG6_34|_PG|B12|B _PG6_34|_PG|B2 _PG6_34|_PG|B12|MID_SHUNT  3.84154647408
L_PG6_34|_PG|B12|RB _PG6_34|_PG|B12|MID_SHUNT _PG6_34|_PG|B3  2.1704737578552e-12
B_PG6_34|_PG|Q2|1 _PG6_34|_PG|Q2 _PG6_34|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_PG|Q2|P _PG6_34|_PG|Q2|MID_SERIES 0  2e-13
R_PG6_34|_PG|Q2|B _PG6_34|_PG|Q2 _PG6_34|_PG|Q2|MID_SHUNT  2.7439617672
L_PG6_34|_PG|Q2|RB _PG6_34|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_PG|Q1|1 _PG6_34|_PG|Q1 _PG6_34|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_PG|Q1|P _PG6_34|_PG|Q1|MID_SERIES 0  2e-13
R_PG6_34|_PG|Q1|B _PG6_34|_PG|Q1 _PG6_34|_PG|Q1|MID_SHUNT  2.7439617672
L_PG6_34|_PG|Q1|RB _PG6_34|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_GG|I_A1|B _PG6_34|_GG|A1 _PG6_34|_GG|I_A1|MID  2e-12
I_PG6_34|_GG|I_A1|B 0 _PG6_34|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_GG|I_B1|B _PG6_34|_GG|B1 _PG6_34|_GG|I_B1|MID  2e-12
I_PG6_34|_GG|I_B1|B 0 _PG6_34|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_GG|I_Q3|B _PG6_34|_GG|Q3 _PG6_34|_GG|I_Q3|MID  2e-12
I_PG6_34|_GG|I_Q3|B 0 _PG6_34|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_34|_GG|I_Q2|B _PG6_34|_GG|Q2 _PG6_34|_GG|I_Q2|MID  2e-12
I_PG6_34|_GG|I_Q2|B 0 _PG6_34|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_GG|I_Q1|B _PG6_34|_GG|Q1 _PG6_34|_GG|I_Q1|MID  2e-12
I_PG6_34|_GG|I_Q1|B 0 _PG6_34|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_GG|A1|1 _PG6_34|_GG|A1 _PG6_34|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_GG|A1|P _PG6_34|_GG|A1|MID_SERIES 0  2e-13
R_PG6_34|_GG|A1|B _PG6_34|_GG|A1 _PG6_34|_GG|A1|MID_SHUNT  2.7439617672
L_PG6_34|_GG|A1|RB _PG6_34|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_GG|A2|1 _PG6_34|_GG|A2 _PG6_34|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_GG|A2|P _PG6_34|_GG|A2|MID_SERIES 0  2e-13
R_PG6_34|_GG|A2|B _PG6_34|_GG|A2 _PG6_34|_GG|A2|MID_SHUNT  2.7439617672
L_PG6_34|_GG|A2|RB _PG6_34|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_GG|A12|1 _PG6_34|_GG|A2 _PG6_34|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_GG|A12|B _PG6_34|_GG|A2 _PG6_34|_GG|A12|MID_SHUNT  3.84154647408
L_PG6_34|_GG|A12|RB _PG6_34|_GG|A12|MID_SHUNT _PG6_34|_GG|A3  2.1704737578552e-12
B_PG6_34|_GG|B1|1 _PG6_34|_GG|B1 _PG6_34|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_GG|B1|P _PG6_34|_GG|B1|MID_SERIES 0  2e-13
R_PG6_34|_GG|B1|B _PG6_34|_GG|B1 _PG6_34|_GG|B1|MID_SHUNT  2.7439617672
L_PG6_34|_GG|B1|RB _PG6_34|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_GG|B2|1 _PG6_34|_GG|B2 _PG6_34|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_GG|B2|P _PG6_34|_GG|B2|MID_SERIES 0  2e-13
R_PG6_34|_GG|B2|B _PG6_34|_GG|B2 _PG6_34|_GG|B2|MID_SHUNT  2.7439617672
L_PG6_34|_GG|B2|RB _PG6_34|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_GG|B12|1 _PG6_34|_GG|B2 _PG6_34|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG6_34|_GG|B12|B _PG6_34|_GG|B2 _PG6_34|_GG|B12|MID_SHUNT  3.84154647408
L_PG6_34|_GG|B12|RB _PG6_34|_GG|B12|MID_SHUNT _PG6_34|_GG|B3  2.1704737578552e-12
B_PG6_34|_GG|Q2|1 _PG6_34|_GG|Q2 _PG6_34|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_GG|Q2|P _PG6_34|_GG|Q2|MID_SERIES 0  2e-13
R_PG6_34|_GG|Q2|B _PG6_34|_GG|Q2 _PG6_34|_GG|Q2|MID_SHUNT  2.7439617672
L_PG6_34|_GG|Q2|RB _PG6_34|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_GG|Q1|1 _PG6_34|_GG|Q1 _PG6_34|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_GG|Q1|P _PG6_34|_GG|Q1|MID_SERIES 0  2e-13
R_PG6_34|_GG|Q1|B _PG6_34|_GG|Q1 _PG6_34|_GG|Q1|MID_SHUNT  2.7439617672
L_PG6_34|_GG|Q1|RB _PG6_34|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_DFF_P0|I_1|B _PG6_34|_DFF_P0|A1 _PG6_34|_DFF_P0|I_1|MID  2e-12
I_PG6_34|_DFF_P0|I_1|B 0 _PG6_34|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_P0|I_3|B _PG6_34|_DFF_P0|A3 _PG6_34|_DFF_P0|I_3|MID  2e-12
I_PG6_34|_DFF_P0|I_3|B 0 _PG6_34|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_34|_DFF_P0|I_T|B _PG6_34|_DFF_P0|T1 _PG6_34|_DFF_P0|I_T|MID  2e-12
I_PG6_34|_DFF_P0|I_T|B 0 _PG6_34|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_P0|I_6|B _PG6_34|_DFF_P0|Q1 _PG6_34|_DFF_P0|I_6|MID  2e-12
I_PG6_34|_DFF_P0|I_6|B 0 _PG6_34|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_DFF_P0|1|1 _PG6_34|_DFF_P0|A1 _PG6_34|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P0|1|P _PG6_34|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P0|1|B _PG6_34|_DFF_P0|A1 _PG6_34|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P0|1|RB _PG6_34|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P0|23|1 _PG6_34|_DFF_P0|A2 _PG6_34|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_P0|23|B _PG6_34|_DFF_P0|A2 _PG6_34|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_P0|23|RB _PG6_34|_DFF_P0|23|MID_SHUNT _PG6_34|_DFF_P0|A3  2.1704737578552e-12
B_PG6_34|_DFF_P0|3|1 _PG6_34|_DFF_P0|A3 _PG6_34|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P0|3|P _PG6_34|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P0|3|B _PG6_34|_DFF_P0|A3 _PG6_34|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P0|3|RB _PG6_34|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P0|4|1 _PG6_34|_DFF_P0|A4 _PG6_34|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P0|4|P _PG6_34|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P0|4|B _PG6_34|_DFF_P0|A4 _PG6_34|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P0|4|RB _PG6_34|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P0|T|1 _PG6_34|_DFF_P0|T1 _PG6_34|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P0|T|P _PG6_34|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P0|T|B _PG6_34|_DFF_P0|T1 _PG6_34|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P0|T|RB _PG6_34|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P0|45|1 _PG6_34|_DFF_P0|T2 _PG6_34|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_P0|45|B _PG6_34|_DFF_P0|T2 _PG6_34|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_P0|45|RB _PG6_34|_DFF_P0|45|MID_SHUNT _PG6_34|_DFF_P0|A4  2.1704737578552e-12
B_PG6_34|_DFF_P0|6|1 _PG6_34|_DFF_P0|Q1 _PG6_34|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P0|6|P _PG6_34|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P0|6|B _PG6_34|_DFF_P0|Q1 _PG6_34|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P0|6|RB _PG6_34|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_DFF_P1|I_1|B _PG6_34|_DFF_P1|A1 _PG6_34|_DFF_P1|I_1|MID  2e-12
I_PG6_34|_DFF_P1|I_1|B 0 _PG6_34|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_P1|I_3|B _PG6_34|_DFF_P1|A3 _PG6_34|_DFF_P1|I_3|MID  2e-12
I_PG6_34|_DFF_P1|I_3|B 0 _PG6_34|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_34|_DFF_P1|I_T|B _PG6_34|_DFF_P1|T1 _PG6_34|_DFF_P1|I_T|MID  2e-12
I_PG6_34|_DFF_P1|I_T|B 0 _PG6_34|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_P1|I_6|B _PG6_34|_DFF_P1|Q1 _PG6_34|_DFF_P1|I_6|MID  2e-12
I_PG6_34|_DFF_P1|I_6|B 0 _PG6_34|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_DFF_P1|1|1 _PG6_34|_DFF_P1|A1 _PG6_34|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P1|1|P _PG6_34|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P1|1|B _PG6_34|_DFF_P1|A1 _PG6_34|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P1|1|RB _PG6_34|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P1|23|1 _PG6_34|_DFF_P1|A2 _PG6_34|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_P1|23|B _PG6_34|_DFF_P1|A2 _PG6_34|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_P1|23|RB _PG6_34|_DFF_P1|23|MID_SHUNT _PG6_34|_DFF_P1|A3  2.1704737578552e-12
B_PG6_34|_DFF_P1|3|1 _PG6_34|_DFF_P1|A3 _PG6_34|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P1|3|P _PG6_34|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P1|3|B _PG6_34|_DFF_P1|A3 _PG6_34|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P1|3|RB _PG6_34|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P1|4|1 _PG6_34|_DFF_P1|A4 _PG6_34|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P1|4|P _PG6_34|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P1|4|B _PG6_34|_DFF_P1|A4 _PG6_34|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P1|4|RB _PG6_34|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P1|T|1 _PG6_34|_DFF_P1|T1 _PG6_34|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P1|T|P _PG6_34|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P1|T|B _PG6_34|_DFF_P1|T1 _PG6_34|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P1|T|RB _PG6_34|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_P1|45|1 _PG6_34|_DFF_P1|T2 _PG6_34|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_P1|45|B _PG6_34|_DFF_P1|T2 _PG6_34|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_P1|45|RB _PG6_34|_DFF_P1|45|MID_SHUNT _PG6_34|_DFF_P1|A4  2.1704737578552e-12
B_PG6_34|_DFF_P1|6|1 _PG6_34|_DFF_P1|Q1 _PG6_34|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_P1|6|P _PG6_34|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG6_34|_DFF_P1|6|B _PG6_34|_DFF_P1|Q1 _PG6_34|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_P1|6|RB _PG6_34|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_DFF_PG|I_1|B _PG6_34|_DFF_PG|A1 _PG6_34|_DFF_PG|I_1|MID  2e-12
I_PG6_34|_DFF_PG|I_1|B 0 _PG6_34|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_PG|I_3|B _PG6_34|_DFF_PG|A3 _PG6_34|_DFF_PG|I_3|MID  2e-12
I_PG6_34|_DFF_PG|I_3|B 0 _PG6_34|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_34|_DFF_PG|I_T|B _PG6_34|_DFF_PG|T1 _PG6_34|_DFF_PG|I_T|MID  2e-12
I_PG6_34|_DFF_PG|I_T|B 0 _PG6_34|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_PG|I_6|B _PG6_34|_DFF_PG|Q1 _PG6_34|_DFF_PG|I_6|MID  2e-12
I_PG6_34|_DFF_PG|I_6|B 0 _PG6_34|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_DFF_PG|1|1 _PG6_34|_DFF_PG|A1 _PG6_34|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_PG|1|P _PG6_34|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG6_34|_DFF_PG|1|B _PG6_34|_DFF_PG|A1 _PG6_34|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_PG|1|RB _PG6_34|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_PG|23|1 _PG6_34|_DFF_PG|A2 _PG6_34|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_PG|23|B _PG6_34|_DFF_PG|A2 _PG6_34|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_PG|23|RB _PG6_34|_DFF_PG|23|MID_SHUNT _PG6_34|_DFF_PG|A3  2.1704737578552e-12
B_PG6_34|_DFF_PG|3|1 _PG6_34|_DFF_PG|A3 _PG6_34|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_PG|3|P _PG6_34|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG6_34|_DFF_PG|3|B _PG6_34|_DFF_PG|A3 _PG6_34|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_PG|3|RB _PG6_34|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_PG|4|1 _PG6_34|_DFF_PG|A4 _PG6_34|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_PG|4|P _PG6_34|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG6_34|_DFF_PG|4|B _PG6_34|_DFF_PG|A4 _PG6_34|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_PG|4|RB _PG6_34|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_PG|T|1 _PG6_34|_DFF_PG|T1 _PG6_34|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_PG|T|P _PG6_34|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG6_34|_DFF_PG|T|B _PG6_34|_DFF_PG|T1 _PG6_34|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_PG|T|RB _PG6_34|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_PG|45|1 _PG6_34|_DFF_PG|T2 _PG6_34|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_PG|45|B _PG6_34|_DFF_PG|T2 _PG6_34|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_PG|45|RB _PG6_34|_DFF_PG|45|MID_SHUNT _PG6_34|_DFF_PG|A4  2.1704737578552e-12
B_PG6_34|_DFF_PG|6|1 _PG6_34|_DFF_PG|Q1 _PG6_34|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_PG|6|P _PG6_34|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG6_34|_DFF_PG|6|B _PG6_34|_DFF_PG|Q1 _PG6_34|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_PG|6|RB _PG6_34|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_DFF_GG|I_1|B _PG6_34|_DFF_GG|A1 _PG6_34|_DFF_GG|I_1|MID  2e-12
I_PG6_34|_DFF_GG|I_1|B 0 _PG6_34|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_GG|I_3|B _PG6_34|_DFF_GG|A3 _PG6_34|_DFF_GG|I_3|MID  2e-12
I_PG6_34|_DFF_GG|I_3|B 0 _PG6_34|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG6_34|_DFF_GG|I_T|B _PG6_34|_DFF_GG|T1 _PG6_34|_DFF_GG|I_T|MID  2e-12
I_PG6_34|_DFF_GG|I_T|B 0 _PG6_34|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_DFF_GG|I_6|B _PG6_34|_DFF_GG|Q1 _PG6_34|_DFF_GG|I_6|MID  2e-12
I_PG6_34|_DFF_GG|I_6|B 0 _PG6_34|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_DFF_GG|1|1 _PG6_34|_DFF_GG|A1 _PG6_34|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_GG|1|P _PG6_34|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG6_34|_DFF_GG|1|B _PG6_34|_DFF_GG|A1 _PG6_34|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_GG|1|RB _PG6_34|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_GG|23|1 _PG6_34|_DFF_GG|A2 _PG6_34|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_GG|23|B _PG6_34|_DFF_GG|A2 _PG6_34|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_GG|23|RB _PG6_34|_DFF_GG|23|MID_SHUNT _PG6_34|_DFF_GG|A3  2.1704737578552e-12
B_PG6_34|_DFF_GG|3|1 _PG6_34|_DFF_GG|A3 _PG6_34|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_GG|3|P _PG6_34|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG6_34|_DFF_GG|3|B _PG6_34|_DFF_GG|A3 _PG6_34|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_GG|3|RB _PG6_34|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_GG|4|1 _PG6_34|_DFF_GG|A4 _PG6_34|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_GG|4|P _PG6_34|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG6_34|_DFF_GG|4|B _PG6_34|_DFF_GG|A4 _PG6_34|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_GG|4|RB _PG6_34|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_GG|T|1 _PG6_34|_DFF_GG|T1 _PG6_34|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_GG|T|P _PG6_34|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG6_34|_DFF_GG|T|B _PG6_34|_DFF_GG|T1 _PG6_34|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_GG|T|RB _PG6_34|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_DFF_GG|45|1 _PG6_34|_DFF_GG|T2 _PG6_34|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG6_34|_DFF_GG|45|B _PG6_34|_DFF_GG|T2 _PG6_34|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG6_34|_DFF_GG|45|RB _PG6_34|_DFF_GG|45|MID_SHUNT _PG6_34|_DFF_GG|A4  2.1704737578552e-12
B_PG6_34|_DFF_GG|6|1 _PG6_34|_DFF_GG|Q1 _PG6_34|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_DFF_GG|6|P _PG6_34|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG6_34|_DFF_GG|6|B _PG6_34|_DFF_GG|Q1 _PG6_34|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG6_34|_DFF_GG|6|RB _PG6_34|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_AND_G|I_A1|B _PG6_34|_AND_G|A1 _PG6_34|_AND_G|I_A1|MID  2e-12
I_PG6_34|_AND_G|I_A1|B 0 _PG6_34|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_AND_G|I_B1|B _PG6_34|_AND_G|B1 _PG6_34|_AND_G|I_B1|MID  2e-12
I_PG6_34|_AND_G|I_B1|B 0 _PG6_34|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_AND_G|I_Q3|B _PG6_34|_AND_G|Q3 _PG6_34|_AND_G|I_Q3|MID  2e-12
I_PG6_34|_AND_G|I_Q3|B 0 _PG6_34|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG6_34|_AND_G|I_Q2|B _PG6_34|_AND_G|Q2 _PG6_34|_AND_G|I_Q2|MID  2e-12
I_PG6_34|_AND_G|I_Q2|B 0 _PG6_34|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_AND_G|I_Q1|B _PG6_34|_AND_G|Q1 _PG6_34|_AND_G|I_Q1|MID  2e-12
I_PG6_34|_AND_G|I_Q1|B 0 _PG6_34|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_AND_G|A1|1 _PG6_34|_AND_G|A1 _PG6_34|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_G|A1|P _PG6_34|_AND_G|A1|MID_SERIES 0  2e-13
R_PG6_34|_AND_G|A1|B _PG6_34|_AND_G|A1 _PG6_34|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG6_34|_AND_G|A1|RB _PG6_34|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_G|A2|1 _PG6_34|_AND_G|A2 _PG6_34|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_G|A2|P _PG6_34|_AND_G|A2|MID_SERIES 0  2e-13
R_PG6_34|_AND_G|A2|B _PG6_34|_AND_G|A2 _PG6_34|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG6_34|_AND_G|A2|RB _PG6_34|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_G|A12|1 _PG6_34|_AND_G|A2 _PG6_34|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_AND_G|A12|B _PG6_34|_AND_G|A2 _PG6_34|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG6_34|_AND_G|A12|RB _PG6_34|_AND_G|A12|MID_SHUNT _PG6_34|_AND_G|A3  2.1704737578552e-12
B_PG6_34|_AND_G|B1|1 _PG6_34|_AND_G|B1 _PG6_34|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_G|B1|P _PG6_34|_AND_G|B1|MID_SERIES 0  2e-13
R_PG6_34|_AND_G|B1|B _PG6_34|_AND_G|B1 _PG6_34|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG6_34|_AND_G|B1|RB _PG6_34|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_G|B2|1 _PG6_34|_AND_G|B2 _PG6_34|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_G|B2|P _PG6_34|_AND_G|B2|MID_SERIES 0  2e-13
R_PG6_34|_AND_G|B2|B _PG6_34|_AND_G|B2 _PG6_34|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG6_34|_AND_G|B2|RB _PG6_34|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_G|B12|1 _PG6_34|_AND_G|B2 _PG6_34|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG6_34|_AND_G|B12|B _PG6_34|_AND_G|B2 _PG6_34|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG6_34|_AND_G|B12|RB _PG6_34|_AND_G|B12|MID_SHUNT _PG6_34|_AND_G|B3  2.1704737578552e-12
B_PG6_34|_AND_G|Q2|1 _PG6_34|_AND_G|Q2 _PG6_34|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_G|Q2|P _PG6_34|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG6_34|_AND_G|Q2|B _PG6_34|_AND_G|Q2 _PG6_34|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG6_34|_AND_G|Q2|RB _PG6_34|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_G|Q1|1 _PG6_34|_AND_G|Q1 _PG6_34|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_G|Q1|P _PG6_34|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG6_34|_AND_G|Q1|B _PG6_34|_AND_G|Q1 _PG6_34|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG6_34|_AND_G|Q1|RB _PG6_34|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG6_34|_AND_P|I_A1|B _PG6_34|_AND_P|A1 _PG6_34|_AND_P|I_A1|MID  2e-12
I_PG6_34|_AND_P|I_A1|B 0 _PG6_34|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_AND_P|I_B1|B _PG6_34|_AND_P|B1 _PG6_34|_AND_P|I_B1|MID  2e-12
I_PG6_34|_AND_P|I_B1|B 0 _PG6_34|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_AND_P|I_Q3|B _PG6_34|_AND_P|Q3 _PG6_34|_AND_P|I_Q3|MID  2e-12
I_PG6_34|_AND_P|I_Q3|B 0 _PG6_34|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG6_34|_AND_P|I_Q2|B _PG6_34|_AND_P|Q2 _PG6_34|_AND_P|I_Q2|MID  2e-12
I_PG6_34|_AND_P|I_Q2|B 0 _PG6_34|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG6_34|_AND_P|I_Q1|B _PG6_34|_AND_P|Q1 _PG6_34|_AND_P|I_Q1|MID  2e-12
I_PG6_34|_AND_P|I_Q1|B 0 _PG6_34|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG6_34|_AND_P|A1|1 _PG6_34|_AND_P|A1 _PG6_34|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_P|A1|P _PG6_34|_AND_P|A1|MID_SERIES 0  2e-13
R_PG6_34|_AND_P|A1|B _PG6_34|_AND_P|A1 _PG6_34|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG6_34|_AND_P|A1|RB _PG6_34|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_P|A2|1 _PG6_34|_AND_P|A2 _PG6_34|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_P|A2|P _PG6_34|_AND_P|A2|MID_SERIES 0  2e-13
R_PG6_34|_AND_P|A2|B _PG6_34|_AND_P|A2 _PG6_34|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG6_34|_AND_P|A2|RB _PG6_34|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_P|A12|1 _PG6_34|_AND_P|A2 _PG6_34|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG6_34|_AND_P|A12|B _PG6_34|_AND_P|A2 _PG6_34|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG6_34|_AND_P|A12|RB _PG6_34|_AND_P|A12|MID_SHUNT _PG6_34|_AND_P|A3  2.1704737578552e-12
B_PG6_34|_AND_P|B1|1 _PG6_34|_AND_P|B1 _PG6_34|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_P|B1|P _PG6_34|_AND_P|B1|MID_SERIES 0  2e-13
R_PG6_34|_AND_P|B1|B _PG6_34|_AND_P|B1 _PG6_34|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG6_34|_AND_P|B1|RB _PG6_34|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_P|B2|1 _PG6_34|_AND_P|B2 _PG6_34|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_P|B2|P _PG6_34|_AND_P|B2|MID_SERIES 0  2e-13
R_PG6_34|_AND_P|B2|B _PG6_34|_AND_P|B2 _PG6_34|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG6_34|_AND_P|B2|RB _PG6_34|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_P|B12|1 _PG6_34|_AND_P|B2 _PG6_34|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG6_34|_AND_P|B12|B _PG6_34|_AND_P|B2 _PG6_34|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG6_34|_AND_P|B12|RB _PG6_34|_AND_P|B12|MID_SHUNT _PG6_34|_AND_P|B3  2.1704737578552e-12
B_PG6_34|_AND_P|Q2|1 _PG6_34|_AND_P|Q2 _PG6_34|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_P|Q2|P _PG6_34|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG6_34|_AND_P|Q2|B _PG6_34|_AND_P|Q2 _PG6_34|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG6_34|_AND_P|Q2|RB _PG6_34|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG6_34|_AND_P|Q1|1 _PG6_34|_AND_P|Q1 _PG6_34|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG6_34|_AND_P|Q1|P _PG6_34|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG6_34|_AND_P|Q1|B _PG6_34|_AND_P|Q1 _PG6_34|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG6_34|_AND_P|Q1|RB _PG6_34|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
L_PTL_G1_1|_SPL|SPL1|I_D1|B _PTL_G1_1|_SPL|SPL1|D1 _PTL_G1_1|_SPL|SPL1|I_D1|MID  2e-12
I_PTL_G1_1|_SPL|SPL1|I_D1|B 0 _PTL_G1_1|_SPL|SPL1|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_SPL|SPL1|I_D2|B _PTL_G1_1|_SPL|SPL1|D2 _PTL_G1_1|_SPL|SPL1|I_D2|MID  2e-12
I_PTL_G1_1|_SPL|SPL1|I_D2|B 0 _PTL_G1_1|_SPL|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G1_1|_SPL|SPL1|I_Q1|B _PTL_G1_1|_SPL|SPL1|QA1 _PTL_G1_1|_SPL|SPL1|I_Q1|MID  2e-12
I_PTL_G1_1|_SPL|SPL1|I_Q1|B 0 _PTL_G1_1|_SPL|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_SPL|SPL1|I_Q2|B _PTL_G1_1|_SPL|SPL1|QB1 _PTL_G1_1|_SPL|SPL1|I_Q2|MID  2e-12
I_PTL_G1_1|_SPL|SPL1|I_Q2|B 0 _PTL_G1_1|_SPL|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G1_1|_SPL|SPL1|1|1 _PTL_G1_1|_SPL|SPL1|D1 _PTL_G1_1|_SPL|SPL1|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL1|1|P _PTL_G1_1|_SPL|SPL1|1|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL1|1|B _PTL_G1_1|_SPL|SPL1|D1 _PTL_G1_1|_SPL|SPL1|1|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL1|1|RB _PTL_G1_1|_SPL|SPL1|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G1_1|_SPL|SPL1|2|1 _PTL_G1_1|_SPL|SPL1|D2 _PTL_G1_1|_SPL|SPL1|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL1|2|P _PTL_G1_1|_SPL|SPL1|2|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL1|2|B _PTL_G1_1|_SPL|SPL1|D2 _PTL_G1_1|_SPL|SPL1|2|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL1|2|RB _PTL_G1_1|_SPL|SPL1|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G1_1|_SPL|SPL1|A|1 _PTL_G1_1|_SPL|SPL1|QA1 _PTL_G1_1|_SPL|SPL1|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL1|A|P _PTL_G1_1|_SPL|SPL1|A|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL1|A|B _PTL_G1_1|_SPL|SPL1|QA1 _PTL_G1_1|_SPL|SPL1|A|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL1|A|RB _PTL_G1_1|_SPL|SPL1|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G1_1|_SPL|SPL1|B|1 _PTL_G1_1|_SPL|SPL1|QB1 _PTL_G1_1|_SPL|SPL1|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL1|B|P _PTL_G1_1|_SPL|SPL1|B|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL1|B|B _PTL_G1_1|_SPL|SPL1|QB1 _PTL_G1_1|_SPL|SPL1|B|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL1|B|RB _PTL_G1_1|_SPL|SPL1|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_G1_1|_SPL|SPL2|I_D1|B _PTL_G1_1|_SPL|SPL2|D1 _PTL_G1_1|_SPL|SPL2|I_D1|MID  2e-12
I_PTL_G1_1|_SPL|SPL2|I_D1|B 0 _PTL_G1_1|_SPL|SPL2|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_SPL|SPL2|I_D2|B _PTL_G1_1|_SPL|SPL2|D2 _PTL_G1_1|_SPL|SPL2|I_D2|MID  2e-12
I_PTL_G1_1|_SPL|SPL2|I_D2|B 0 _PTL_G1_1|_SPL|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_G1_1|_SPL|SPL2|I_Q1|B _PTL_G1_1|_SPL|SPL2|QA1 _PTL_G1_1|_SPL|SPL2|I_Q1|MID  2e-12
I_PTL_G1_1|_SPL|SPL2|I_Q1|B 0 _PTL_G1_1|_SPL|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_G1_1|_SPL|SPL2|I_Q2|B _PTL_G1_1|_SPL|SPL2|QB1 _PTL_G1_1|_SPL|SPL2|I_Q2|MID  2e-12
I_PTL_G1_1|_SPL|SPL2|I_Q2|B 0 _PTL_G1_1|_SPL|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_G1_1|_SPL|SPL2|1|1 _PTL_G1_1|_SPL|SPL2|D1 _PTL_G1_1|_SPL|SPL2|1|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL2|1|P _PTL_G1_1|_SPL|SPL2|1|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL2|1|B _PTL_G1_1|_SPL|SPL2|D1 _PTL_G1_1|_SPL|SPL2|1|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL2|1|RB _PTL_G1_1|_SPL|SPL2|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_G1_1|_SPL|SPL2|2|1 _PTL_G1_1|_SPL|SPL2|D2 _PTL_G1_1|_SPL|SPL2|2|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL2|2|P _PTL_G1_1|_SPL|SPL2|2|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL2|2|B _PTL_G1_1|_SPL|SPL2|D2 _PTL_G1_1|_SPL|SPL2|2|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL2|2|RB _PTL_G1_1|_SPL|SPL2|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_G1_1|_SPL|SPL2|A|1 _PTL_G1_1|_SPL|SPL2|QA1 _PTL_G1_1|_SPL|SPL2|A|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL2|A|P _PTL_G1_1|_SPL|SPL2|A|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL2|A|B _PTL_G1_1|_SPL|SPL2|QA1 _PTL_G1_1|_SPL|SPL2|A|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL2|A|RB _PTL_G1_1|_SPL|SPL2|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_G1_1|_SPL|SPL2|B|1 _PTL_G1_1|_SPL|SPL2|QB1 _PTL_G1_1|_SPL|SPL2|B|MID_SERIES JJMIT AREA=2.5
L_PTL_G1_1|_SPL|SPL2|B|P _PTL_G1_1|_SPL|SPL2|B|MID_SERIES 0  2e-13
R_PTL_G1_1|_SPL|SPL2|B|B _PTL_G1_1|_SPL|SPL2|QB1 _PTL_G1_1|_SPL|SPL2|B|MID_SHUNT  2.7439617672
L_PTL_G1_1|_SPL|SPL2|B|RB _PTL_G1_1|_SPL|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_P3_2|_SPL|SPL1|I_D1|B _PTL_P3_2|_SPL|SPL1|D1 _PTL_P3_2|_SPL|SPL1|I_D1|MID  2e-12
I_PTL_P3_2|_SPL|SPL1|I_D1|B 0 _PTL_P3_2|_SPL|SPL1|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P3_2|_SPL|SPL1|I_D2|B _PTL_P3_2|_SPL|SPL1|D2 _PTL_P3_2|_SPL|SPL1|I_D2|MID  2e-12
I_PTL_P3_2|_SPL|SPL1|I_D2|B 0 _PTL_P3_2|_SPL|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P3_2|_SPL|SPL1|I_Q1|B _PTL_P3_2|_SPL|SPL1|QA1 _PTL_P3_2|_SPL|SPL1|I_Q1|MID  2e-12
I_PTL_P3_2|_SPL|SPL1|I_Q1|B 0 _PTL_P3_2|_SPL|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P3_2|_SPL|SPL1|I_Q2|B _PTL_P3_2|_SPL|SPL1|QB1 _PTL_P3_2|_SPL|SPL1|I_Q2|MID  2e-12
I_PTL_P3_2|_SPL|SPL1|I_Q2|B 0 _PTL_P3_2|_SPL|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P3_2|_SPL|SPL1|1|1 _PTL_P3_2|_SPL|SPL1|D1 _PTL_P3_2|_SPL|SPL1|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL1|1|P _PTL_P3_2|_SPL|SPL1|1|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL1|1|B _PTL_P3_2|_SPL|SPL1|D1 _PTL_P3_2|_SPL|SPL1|1|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL1|1|RB _PTL_P3_2|_SPL|SPL1|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P3_2|_SPL|SPL1|2|1 _PTL_P3_2|_SPL|SPL1|D2 _PTL_P3_2|_SPL|SPL1|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL1|2|P _PTL_P3_2|_SPL|SPL1|2|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL1|2|B _PTL_P3_2|_SPL|SPL1|D2 _PTL_P3_2|_SPL|SPL1|2|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL1|2|RB _PTL_P3_2|_SPL|SPL1|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P3_2|_SPL|SPL1|A|1 _PTL_P3_2|_SPL|SPL1|QA1 _PTL_P3_2|_SPL|SPL1|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL1|A|P _PTL_P3_2|_SPL|SPL1|A|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL1|A|B _PTL_P3_2|_SPL|SPL1|QA1 _PTL_P3_2|_SPL|SPL1|A|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL1|A|RB _PTL_P3_2|_SPL|SPL1|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P3_2|_SPL|SPL1|B|1 _PTL_P3_2|_SPL|SPL1|QB1 _PTL_P3_2|_SPL|SPL1|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL1|B|P _PTL_P3_2|_SPL|SPL1|B|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL1|B|B _PTL_P3_2|_SPL|SPL1|QB1 _PTL_P3_2|_SPL|SPL1|B|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL1|B|RB _PTL_P3_2|_SPL|SPL1|B|MID_SHUNT 0  1.550338398468e-12
L_PTL_P3_2|_SPL|SPL2|I_D1|B _PTL_P3_2|_SPL|SPL2|D1 _PTL_P3_2|_SPL|SPL2|I_D1|MID  2e-12
I_PTL_P3_2|_SPL|SPL2|I_D1|B 0 _PTL_P3_2|_SPL|SPL2|I_D1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P3_2|_SPL|SPL2|I_D2|B _PTL_P3_2|_SPL|SPL2|D2 _PTL_P3_2|_SPL|SPL2|I_D2|MID  2e-12
I_PTL_P3_2|_SPL|SPL2|I_D2|B 0 _PTL_P3_2|_SPL|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000245)
L_PTL_P3_2|_SPL|SPL2|I_Q1|B _PTL_P3_2|_SPL|SPL2|QA1 _PTL_P3_2|_SPL|SPL2|I_Q1|MID  2e-12
I_PTL_P3_2|_SPL|SPL2|I_Q1|B 0 _PTL_P3_2|_SPL|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
L_PTL_P3_2|_SPL|SPL2|I_Q2|B _PTL_P3_2|_SPL|SPL2|QB1 _PTL_P3_2|_SPL|SPL2|I_Q2|MID  2e-12
I_PTL_P3_2|_SPL|SPL2|I_Q2|B 0 _PTL_P3_2|_SPL|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.000175)
B_PTL_P3_2|_SPL|SPL2|1|1 _PTL_P3_2|_SPL|SPL2|D1 _PTL_P3_2|_SPL|SPL2|1|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL2|1|P _PTL_P3_2|_SPL|SPL2|1|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL2|1|B _PTL_P3_2|_SPL|SPL2|D1 _PTL_P3_2|_SPL|SPL2|1|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL2|1|RB _PTL_P3_2|_SPL|SPL2|1|MID_SHUNT 0  1.550338398468e-12
B_PTL_P3_2|_SPL|SPL2|2|1 _PTL_P3_2|_SPL|SPL2|D2 _PTL_P3_2|_SPL|SPL2|2|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL2|2|P _PTL_P3_2|_SPL|SPL2|2|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL2|2|B _PTL_P3_2|_SPL|SPL2|D2 _PTL_P3_2|_SPL|SPL2|2|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL2|2|RB _PTL_P3_2|_SPL|SPL2|2|MID_SHUNT 0  1.550338398468e-12
B_PTL_P3_2|_SPL|SPL2|A|1 _PTL_P3_2|_SPL|SPL2|QA1 _PTL_P3_2|_SPL|SPL2|A|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL2|A|P _PTL_P3_2|_SPL|SPL2|A|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL2|A|B _PTL_P3_2|_SPL|SPL2|QA1 _PTL_P3_2|_SPL|SPL2|A|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL2|A|RB _PTL_P3_2|_SPL|SPL2|A|MID_SHUNT 0  1.550338398468e-12
B_PTL_P3_2|_SPL|SPL2|B|1 _PTL_P3_2|_SPL|SPL2|QB1 _PTL_P3_2|_SPL|SPL2|B|MID_SERIES JJMIT AREA=2.5
L_PTL_P3_2|_SPL|SPL2|B|P _PTL_P3_2|_SPL|SPL2|B|MID_SERIES 0  2e-13
R_PTL_P3_2|_SPL|SPL2|B|B _PTL_P3_2|_SPL|SPL2|QB1 _PTL_P3_2|_SPL|SPL2|B|MID_SHUNT  2.7439617672
L_PTL_P3_2|_SPL|SPL2|B|RB _PTL_P3_2|_SPL|SPL2|B|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_S0
.print DEVI R_S1
.print DEVI R_S2
.print DEVI R_S3
.print DEVI R_S4
.print DEVI R_S5
.print DEVI R_S6
.print DEVI R_S7
.print DEVI R_S8
.print V B5_RX
.print V G6_3_TO6
.print V B4_TX
.print V T32
.print V IP4_0
.print V G2_2_OUT
.print V G1_1_TO2
.print V T1A
.print V G5_1_TO7
.print V B3_RX
.print V P7_2_TO7
.print V IP0_0
.print V S0_1
.print V IP7_3_OUT
.print V S1_3
.print V G2_2_TX
.print V S8_4
.print V S0_2
.print V T22
.print V P6_1_TX
.print V S0_5
.print V P5_3_TX
.print V IP7_4_OUT_TX
.print V G5_2_TO5
.print V T31
.print V IP6_0_TO6
.print V IP2_0_TO2
.print V P2_1_TO2
.print V P3_2_TX
.print V IP5_3_OUT
.print V S1_5
.print V S0_2_TX
.print V S1_1_TX
.print V S0_3
.print V A3_TX
.print V T54
.print V G4_1_TX
.print V G3_2_TO7
.print V T2A
.print V P6_3_TX
.print V T06
.print V P3_2_TO7
.print V IP0_0_TO1
.print V G5_1_TO5
.print V P4_1_TX
.print V T36
.print V P3_1_TO3
.print V IG2_0_TO2
.print V P7_1_TO7
.print V A5_RX
.print V T11
.print V S4_5_TX
.print V P4_2_TO4
.print V IP6_0
.print V IP5_0_TO5
.print V T28
.print V T24
.print V IG4_0_TO4
.print V T23
.print V IP2_0
.print V T38
.print V IP1_0
.print V B7_TX
.print V S8_4_TX
.print V S8_3
.print V P7_3_TX
.print V T3A
.print V G5_3_TO6
.print V T51
.print V P2_1_TX
.print V IP3_2_OUT
.print V T19
.print V G7_2_TO7
.print V P7_1_TX
.print V T10
.print V P7_2_TX
.print V T47
.print V G4_2_TO4
.print V A6_RX
.print V G2_1_TO2
.print V G4_3_TX
.print V G4_1_TO4
.print V IG1_0_TO1
.print V S0_1_TX
.print V B1_RX
.print V B0_RX
.print V G6_1_TX
.print V T49
.print V S1_2_TX
.print V G7_1_TX
.print V B1_TX
.print V IP5_1_OUT
.print V S3_4
.print V P1_1_TO2
.print V P6_3_OUT
.print V T03
.print V T30
.print V IG4_0_TO5
.print V T21
.print V P5_2_TX
.print V B2_TX
.print V S8_5
.print V T12
.print V A0_TX
.print V IG5_0
.print V T42
.print V A5_TX
.print V IP7_0
.print V S3_4_TX
.print V T04
.print V T26
.print V S8_5_TX
.print V T17
.print V S7_4_TX
.print V IP7_4_OUT
.print V S3_5_TX
.print V P3_2_TO4
.print V G3_2_OUT
.print V S1_5_TX
.print V G7_1_TO7
.print V T57
.print V S8_3_TX
.print V T18
.print V IP2_0_TO3
.print V T56
.print V G3_2_TO5
.print V G5_1_TX
.print V S0_4_TX
.print V A7_RX
.print V IG7_0_TO7
.print V IP5_2_OUT
.print V IP7_2_OUT
.print V S4_5
.print V G1_1_TO3
.print V S3_3_TX
.print V IG7_0
.print V IP3_0
.print V P1_1_TO3
.print V T44
.print V P3_1_TX
.print V P2_1_OUT
.print V T05
.print V B6_RX
.print V IP5_0
.print V G3_1_TX
.print V P4_3_TX
.print V G6_4_TX
.print V S1_1
.print V S2_3
.print V P5_1_TO5
.print V A3_RX
.print V P6_3_TO6
.print V T02
.print V IG0_0_TO1
.print V T52
.print V T1B
.print V IP4_0_TO4
.print V P6_2_TX
.print V S6_5_TX
.print V T14
.print V S2_4_TX
.print V T13
.print V S1_4
.print V IP5_1_OUT_TX
.print V T00
.print V G3_1_TO3
.print V B2_RX
.print V G5_3_OUT
.print V IP5_3_OUT_TX
.print V P4_1_TO4
.print V IP7_2_OUT_TX
.print V IG6_0
.print V S5_5
.print V IP7_1_OUT
.print V A1_RX
.print V P2_2_TX
.print V IP3_0_TO3
.print V P6_4_TX
.print V IP5_0_OUT
.print V T45
.print V P4_2_TX
.print V S3_5
.print V T20
.print V G2_1_TX
.print V G1_1_TX
.print V A4_TX
.print V G6_2_TX
.print V T40
.print V S6_4
.print V IP3_0_OUT
.print V IG3_0
.print V A6_TX
.print V P5_3_TO6
.print V IP6_0_TO7
.print V P5_2_TO5
.print V S6_4_TX
.print V B5_TX
.print V B7_RX
.print V A4_RX
.print V S3_3
.print V P5_1_TO7
.print V B4_RX
.print V S2_2_TX
.print V T01
.print V S2_4
.print V S2_5
.print V IG0_0
.print V G7_2_TX
.print V IP3_2_OUT_TX
.print V P5_1_TX
.print V S1_2
.print V IP7_0_OUT
.print V IP1_0_OUT
.print V IG3_0_TO3
.print V IG1_0
.print V T39
.print V S1_4_TX
.print V B6_TX
.print V IG5_0_TO5
.print V A0_RX
.print V G3_2_TX
.print V S5_5_TX
.print V G6_4_OUT
.print V P6_1_TO6
.print V IG6_0_TO6
.print V IG4_0
.print V S2_5_TX
.print V T2B
.print V T07
.print V A7_TX
.print V G6_2_TO6
.print V S0_5_TX
.print V S5_4_TX
.print V S7_5
.print V T46
.print V T15
.print V T50
.print V T53
.print V S2_3_TX
.print V S6_5
.print V IP7_3_OUT_TX
.print V T16
.print V IP5_2_OUT_TX
.print V G4_2_TX
.print V T29
.print V S5_4
.print V P3_2_TO5
.print V S2_2
.print V G6_3_TX
.print V S0_3_TX
.print V G4_3_OUT
.print V S0_0
.print V IP3_1_OUT
.print V P6_2_TO6
.print V S7_5_TX
.print V T27
.print V P4_2_OUT
.print V T41
.print V G1_1_OUT
.print V T33
.print V T25
.print V S1_3_TX
.print V G5_3_TX
.print V S0_4
.print V S4_4
.print V IP4_0_TO5
.print V T34
.print V IG0_0_TO0
.print V B0_TX
.print V B3_TX
.print V S4_4_TX
.print V T58
.print V A2_TX
.print V IP7_0_TO7
.print V A2_RX
.print V IG6_0_TO7
.print V S4_3_TX
.print V T48
.print V IG2_0
.print V T37
.print V P1_1_TX
.print V G3_2_TO4
.print V T35
.print V IP7_1_OUT_TX
.print V IG2_0_TO3
.print V T43
.print V S4_3
.print V A1_TX
.print V IP1_0_TO1
.print V G6_1_TO6
.print V G5_2_TX
.print V IP3_1_OUT_TX
.print V T55
