*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=1e-10
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.5E-12 12E-09
ROUT1 AB_XOR_CD_1 0  1
ROUT2 NOT_AB_1 0  1
IT1|T 0 T1  PWL(0 0 3.97e-10 0 4e-10 0.001 4.03e-10 0 6.97e-10 0 7e-10 0.001 7.03e-10 0 9.97e-10 0 1e-09 0.001 1.003e-09 0 1.297e-09 0 1.3e-09 0.001 1.303e-09 0 1.597e-09 0 1.6e-09 0.001 1.603e-09 0 1.897e-09 0 1.9e-09 0.001 1.903e-09 0 2.197e-09 0 2.2e-09 0.001 2.203e-09 0 2.497e-09 0 2.5e-09 0.001 2.503e-09 0 2.797e-09 0 2.8e-09 0.001 2.803e-09 0 3.097e-09 0 3.1e-09 0.001 3.103e-09 0 3.397e-09 0 3.4e-09 0.001 3.403e-09 0 3.697e-09 0 3.7e-09 0.001 3.703e-09 0 3.997e-09 0 4e-09 0.001 4.003e-09 0 4.297e-09 0 4.3e-09 0.001 4.303e-09 0 4.597e-09 0 4.6e-09 0.001 4.603e-09 0 4.897e-09 0 4.9e-09 0.001 4.903e-09 0 5.197e-09 0 5.2e-09 0.001 5.203e-09 0 5.497e-09 0 5.5e-09 0.001 5.503e-09 0 5.797e-09 0 5.8e-09 0.001 5.803e-09 0 6.097e-09 0 6.1e-09 0.001 6.103e-09 0 6.397e-09 0 6.4e-09 0.001 6.403e-09 0 6.697e-09 0 6.7e-09 0.001 6.703e-09 0 6.997e-09 0 7e-09 0.001 7.003e-09 0 7.297e-09 0 7.3e-09 0.001 7.303e-09 0 7.597e-09 0 7.6e-09 0.001 7.603e-09 0 7.897e-09 0 7.9e-09 0.001 7.903e-09 0 8.197e-09 0 8.2e-09 0.001 8.203e-09 0 8.497e-09 0 8.5e-09 0.001 8.503e-09 0 8.797e-09 0 8.8e-09 0.001 8.803e-09 0 9.097e-09 0 9.1e-09 0.001 9.103e-09 0 9.397e-09 0 9.4e-09 0.001 9.403e-09 0 9.697e-09 0 9.7e-09 0.001 9.703e-09 0 9.997e-09 0 1e-08 0.001 1.0003e-08 0 1.0297e-08 0 1.03e-08 0.001 1.0303e-08 0 1.0597e-08 0 1.06e-08 0.001 1.0603e-08 0 1.0897e-08 0 1.09e-08 0.001 1.0903e-08 0 1.1197e-08 0 1.12e-08 0.001 1.1203e-08 0 1.1497e-08 0 1.15e-08 0.001 1.1503e-08 0 1.1797e-08 0 1.18e-08 0.001 1.1803e-08 0)
IT2|T 0 T2  PWL(0 0 2.97e-10 0 3e-10 0.001 3.03e-10 0 5.97e-10 0 6e-10 0.001 6.03e-10 0 8.97e-10 0 9e-10 0.001 9.03e-10 0 1.197e-09 0 1.2e-09 0.001 1.203e-09 0 1.497e-09 0 1.5e-09 0.001 1.503e-09 0 1.797e-09 0 1.8e-09 0.001 1.803e-09 0 2.097e-09 0 2.1e-09 0.001 2.103e-09 0 2.397e-09 0 2.4e-09 0.001 2.403e-09 0 2.697e-09 0 2.7e-09 0.001 2.703e-09 0 2.997e-09 0 3e-09 0.001 3.003e-09 0 3.297e-09 0 3.3e-09 0.001 3.303e-09 0 3.597e-09 0 3.6e-09 0.001 3.603e-09 0 3.897e-09 0 3.9e-09 0.001 3.903e-09 0 4.197e-09 0 4.2e-09 0.001 4.203e-09 0 4.497e-09 0 4.5e-09 0.001 4.503e-09 0 4.797e-09 0 4.8e-09 0.001 4.803e-09 0 5.097e-09 0 5.1e-09 0.001 5.103e-09 0 5.397e-09 0 5.4e-09 0.001 5.403e-09 0 5.697e-09 0 5.7e-09 0.001 5.703e-09 0 5.997e-09 0 6e-09 0.001 6.003e-09 0 6.297e-09 0 6.3e-09 0.001 6.303e-09 0 6.597e-09 0 6.6e-09 0.001 6.603e-09 0 6.897e-09 0 6.9e-09 0.001 6.903e-09 0 7.197e-09 0 7.2e-09 0.001 7.203e-09 0 7.497e-09 0 7.5e-09 0.001 7.503e-09 0 7.797e-09 0 7.8e-09 0.001 7.803e-09 0 8.097e-09 0 8.1e-09 0.001 8.103e-09 0 8.397e-09 0 8.4e-09 0.001 8.403e-09 0 8.697e-09 0 8.7e-09 0.001 8.703e-09 0 8.997e-09 0 9e-09 0.001 9.003e-09 0 9.297e-09 0 9.3e-09 0.001 9.303e-09 0 9.597e-09 0 9.6e-09 0.001 9.603e-09 0 9.897e-09 0 9.9e-09 0.001 9.903e-09 0 1.0197e-08 0 1.02e-08 0.001 1.0203e-08 0 1.0497e-08 0 1.05e-08 0.001 1.0503e-08 0 1.0797e-08 0 1.08e-08 0.001 1.0803e-08 0 1.1097e-08 0 1.11e-08 0.001 1.1103e-08 0 1.1397e-08 0 1.14e-08 0.001 1.1403e-08 0 1.1697e-08 0 1.17e-08 0.001 1.1703e-08 0)
IDATA_A1|A 0 A1  PWL(0 0 7.57e-10 0 7.6e-10 0.0005 7.63e-10 0 1.357e-09 0 1.36e-09 0.0005 1.363e-09 0 1.957e-09 0 1.96e-09 0.0005 1.963e-09 0 2.557e-09 0 2.56e-09 0.0005 2.563e-09 0 3.157e-09 0 3.16e-09 0.0005 3.163e-09 0 3.757e-09 0 3.76e-09 0.0005 3.763e-09 0 4.357e-09 0 4.36e-09 0.0005 4.363e-09 0 4.957e-09 0 4.96e-09 0.0005 4.963e-09 0 5.557e-09 0 5.56e-09 0.0005 5.563e-09 0 6.157e-09 0 6.16e-09 0.0005 6.163e-09 0 6.757e-09 0 6.76e-09 0.0005 6.763e-09 0 7.357e-09 0 7.36e-09 0.0005 7.363e-09 0 7.957e-09 0 7.96e-09 0.0005 7.963e-09 0 8.557e-09 0 8.56e-09 0.0005 8.563e-09 0 9.157e-09 0 9.16e-09 0.0005 9.163e-09 0 9.757e-09 0 9.76e-09 0.0005 9.763e-09 0 1.0357e-08 0 1.036e-08 0.0005 1.0363e-08 0 1.0957e-08 0 1.096e-08 0.0005 1.0963e-08 0 1.1557e-08 0 1.156e-08 0.0005 1.1563e-08 0)
IDATA_B1|B 0 B1  PWL(0 0 1.117e-09 0 1.12e-09 0.0005 1.123e-09 0 1.417e-09 0 1.42e-09 0.0005 1.423e-09 0 2.317e-09 0 2.32e-09 0.0005 2.323e-09 0 2.617e-09 0 2.62e-09 0.0005 2.623e-09 0 3.517e-09 0 3.52e-09 0.0005 3.523e-09 0 3.817e-09 0 3.82e-09 0.0005 3.823e-09 0 4.717e-09 0 4.72e-09 0.0005 4.723e-09 0 5.017e-09 0 5.02e-09 0.0005 5.023e-09 0 5.917e-09 0 5.92e-09 0.0005 5.923e-09 0 6.217e-09 0 6.22e-09 0.0005 6.223e-09 0 7.117e-09 0 7.12e-09 0.0005 7.123e-09 0 7.417e-09 0 7.42e-09 0.0005 7.423e-09 0 8.317e-09 0 8.32e-09 0.0005 8.323e-09 0 8.617e-09 0 8.62e-09 0.0005 8.623e-09 0 9.517e-09 0 9.52e-09 0.0005 9.523e-09 0 9.817e-09 0 9.82e-09 0.0005 9.823e-09 0 1.0717e-08 0 1.072e-08 0.0005 1.0723e-08 0 1.1017e-08 0 1.102e-08 0.0005 1.1023e-08 0 1.1917e-08 0 1.192e-08 0.0005 1.1923e-08 0)
IDATA_C1|T 0 C1  PWL(0 0 1.777e-09 0 1.78e-09 0.0005 1.783e-09 0 2.077e-09 0 2.08e-09 0.0005 2.083e-09 0 2.377e-09 0 2.38e-09 0.0005 2.383e-09 0 2.677e-09 0 2.68e-09 0.0005 2.683e-09 0 4.177e-09 0 4.18e-09 0.0005 4.183e-09 0 4.477e-09 0 4.48e-09 0.0005 4.483e-09 0 4.777e-09 0 4.78e-09 0.0005 4.783e-09 0 5.077e-09 0 5.08e-09 0.0005 5.083e-09 0 6.577e-09 0 6.58e-09 0.0005 6.583e-09 0 6.877e-09 0 6.88e-09 0.0005 6.883e-09 0 7.177e-09 0 7.18e-09 0.0005 7.183e-09 0 7.477e-09 0 7.48e-09 0.0005 7.483e-09 0 8.977e-09 0 8.98e-09 0.0005 8.983e-09 0 9.277e-09 0 9.28e-09 0.0005 9.283e-09 0 9.577e-09 0 9.58e-09 0.0005 9.583e-09 0 9.877e-09 0 9.88e-09 0.0005 9.883e-09 0 1.1377e-08 0 1.138e-08 0.0005 1.1383e-08 0 1.1677e-08 0 1.168e-08 0.0005 1.1683e-08 0 1.1977e-08 0 1.198e-08 0.0005 1.1983e-08 0)
IDATA_D1|T 0 D1  PWL(0 0 3.037e-09 0 3.04e-09 0.0005 3.043e-09 0 3.337e-09 0 3.34e-09 0.0005 3.343e-09 0 3.637e-09 0 3.64e-09 0.0005 3.643e-09 0 3.937e-09 0 3.94e-09 0.0005 3.943e-09 0 4.237e-09 0 4.24e-09 0.0005 4.243e-09 0 4.537e-09 0 4.54e-09 0.0005 4.543e-09 0 4.837e-09 0 4.84e-09 0.0005 4.843e-09 0 5.137e-09 0 5.14e-09 0.0005 5.143e-09 0 7.837e-09 0 7.84e-09 0.0005 7.843e-09 0 8.137e-09 0 8.14e-09 0.0005 8.143e-09 0 8.437e-09 0 8.44e-09 0.0005 8.443e-09 0 8.737e-09 0 8.74e-09 0.0005 8.743e-09 0 9.037e-09 0 9.04e-09 0.0005 9.043e-09 0 9.337e-09 0 9.34e-09 0.0005 9.343e-09 0 9.637e-09 0 9.64e-09 0.0005 9.643e-09 0 9.937e-09 0 9.94e-09 0.0005 9.943e-09 0)
L1|_AND_AB|1 A1 1|_AND_AB|A1  2.067833848e-12
L1|_AND_AB|2 1|_AND_AB|A1 1|_AND_AB|A2  4.135667696e-12
L1|_AND_AB|3 1|_AND_AB|A3 1|_AND_AB|A4  8.271335392e-12
L1|_AND_AB|4 1|_AND_AB|TA 1|_AND_AB|T3  1e-12
L1|_AND_AB|5 1|_AND_AB|A4 1|_AND_AB|A5  4.135667696e-12
L1|_AND_AB|6 B1 1|_AND_AB|B1  2.067833848e-12
L1|_AND_AB|7 1|_AND_AB|B1 1|_AND_AB|B2  4.135667696e-12
L1|_AND_AB|8 1|_AND_AB|B3 1|_AND_AB|B4  8.271335392e-12
L1|_AND_AB|9 1|_AND_AB|TB 1|_AND_AB|T3  1e-12
L1|_AND_AB|10 1|_AND_AB|B4 1|_AND_AB|B5  4.135667696e-12
L1|_AND_AB|11 T1 1|_AND_AB|T1  2.067833848e-12
L1|_AND_AB|12 1|_AND_AB|T1 1|_AND_AB|T2  4.135667696e-12
L1|_AND_AB|13 1|_AND_AB|T2 1|_AND_AB|T3  1e-12
L1|_AND_AB|14 1|_AND_AB|Q2 1|_AND_AB|Q1  1e-12
L1|_AND_AB|15 1|_AND_AB|Q1 1|AB_0  2.067833848e-12
L1|_AND_CD|1 C1 1|_AND_CD|A1  2.067833848e-12
L1|_AND_CD|2 1|_AND_CD|A1 1|_AND_CD|A2  4.135667696e-12
L1|_AND_CD|3 1|_AND_CD|A3 1|_AND_CD|A4  8.271335392e-12
L1|_AND_CD|4 1|_AND_CD|TA 1|_AND_CD|T3  1e-12
L1|_AND_CD|5 1|_AND_CD|A4 1|_AND_CD|A5  4.135667696e-12
L1|_AND_CD|6 D1 1|_AND_CD|B1  2.067833848e-12
L1|_AND_CD|7 1|_AND_CD|B1 1|_AND_CD|B2  4.135667696e-12
L1|_AND_CD|8 1|_AND_CD|B3 1|_AND_CD|B4  8.271335392e-12
L1|_AND_CD|9 1|_AND_CD|TB 1|_AND_CD|T3  1e-12
L1|_AND_CD|10 1|_AND_CD|B4 1|_AND_CD|B5  4.135667696e-12
L1|_AND_CD|11 T1 1|_AND_CD|T1  2.067833848e-12
L1|_AND_CD|12 1|_AND_CD|T1 1|_AND_CD|T2  4.135667696e-12
L1|_AND_CD|13 1|_AND_CD|T2 1|_AND_CD|T3  1e-12
L1|_AND_CD|14 1|_AND_CD|Q2 1|_AND_CD|Q1  1e-12
L1|_AND_CD|15 1|_AND_CD|Q1 1|CD_0  2.067833848e-12
B1|D1|1 1|D1|1 1|D1|2 JJMIT AREA=2.5
B1|D1|2 1|D1|4 1|D1|5 JJMIT AREA=2.5
B1|D1|3 1|D1|7 1|D1|8 JJMIT AREA=2.5
B1|D1|4 1|D1|10 1|D1|11 JJMIT AREA=2.5
I1|D1|B1 0 1|D1|3  PWL(0 0 5e-12 0.000175)
I1|D1|B2 0 1|D1|6  PWL(0 0 5e-12 0.0002375)
I1|D1|B3 0 1|D1|9  PWL(0 0 5e-12 0.0002375)
I1|D1|B4 0 1|D1|12  PWL(0 0 5e-12 0.000175)
L1|D1|1 1|AB_0 1|D1|1  2.067833848e-12
L1|D1|2 1|D1|1 1|D1|4  4.135667696e-12
L1|D1|3 1|D1|4 1|D1|7  4.135667696e-12
L1|D1|4 1|D1|7 1|D1|10  4.135667696e-12
L1|D1|5 1|D1|10 1|AB_1  2.067833848e-12
L1|D1|P1 1|D1|2 0  5e-13
L1|D1|P2 1|D1|5 0  5e-13
L1|D1|P3 1|D1|8 0  5e-13
L1|D1|P4 1|D1|11 0  5e-13
L1|D1|B1 1|D1|1 1|D1|3  2e-12
L1|D1|B2 1|D1|4 1|D1|6  2e-12
L1|D1|B3 1|D1|7 1|D1|9  2e-12
L1|D1|B4 1|D1|10 1|D1|12  2e-12
R1|D1|B1 1|D1|1 1|D1|101  2.7439617672
R1|D1|B2 1|D1|4 1|D1|104  2.7439617672
R1|D1|B3 1|D1|7 1|D1|107  2.7439617672
R1|D1|B4 1|D1|10 1|D1|110  2.7439617672
L1|D1|RB1 1|D1|101 0  2.050338398468e-12
L1|D1|RB2 1|D1|104 0  2.050338398468e-12
L1|D1|RB3 1|D1|107 0  2.050338398468e-12
L1|D1|RB4 1|D1|110 0  2.050338398468e-12
B1|D2|1 1|D2|1 1|D2|2 JJMIT AREA=2.5
B1|D2|2 1|D2|4 1|D2|5 JJMIT AREA=2.5
B1|D2|3 1|D2|7 1|D2|8 JJMIT AREA=2.5
B1|D2|4 1|D2|10 1|D2|11 JJMIT AREA=2.5
I1|D2|B1 0 1|D2|3  PWL(0 0 5e-12 0.000175)
I1|D2|B2 0 1|D2|6  PWL(0 0 5e-12 0.0002375)
I1|D2|B3 0 1|D2|9  PWL(0 0 5e-12 0.0002375)
I1|D2|B4 0 1|D2|12  PWL(0 0 5e-12 0.000175)
L1|D2|1 1|CD_0 1|D2|1  2.067833848e-12
L1|D2|2 1|D2|1 1|D2|4  4.135667696e-12
L1|D2|3 1|D2|4 1|D2|7  4.135667696e-12
L1|D2|4 1|D2|7 1|D2|10  4.135667696e-12
L1|D2|5 1|D2|10 1|CD_1  2.067833848e-12
L1|D2|P1 1|D2|2 0  5e-13
L1|D2|P2 1|D2|5 0  5e-13
L1|D2|P3 1|D2|8 0  5e-13
L1|D2|P4 1|D2|11 0  5e-13
L1|D2|B1 1|D2|1 1|D2|3  2e-12
L1|D2|B2 1|D2|4 1|D2|6  2e-12
L1|D2|B3 1|D2|7 1|D2|9  2e-12
L1|D2|B4 1|D2|10 1|D2|12  2e-12
R1|D2|B1 1|D2|1 1|D2|101  2.7439617672
R1|D2|B2 1|D2|4 1|D2|104  2.7439617672
R1|D2|B3 1|D2|7 1|D2|107  2.7439617672
R1|D2|B4 1|D2|10 1|D2|110  2.7439617672
L1|D2|RB1 1|D2|101 0  2.050338398468e-12
L1|D2|RB2 1|D2|104 0  2.050338398468e-12
L1|D2|RB3 1|D2|107 0  2.050338398468e-12
L1|D2|RB4 1|D2|110 0  2.050338398468e-12
B1|D3|1 1|D3|1 1|D3|2 JJMIT AREA=2.5
B1|D3|2 1|D3|6 1|D3|7 JJMIT AREA=2.5
I1|D3|B1 0 1|D3|5  0.00035
L1|D3|1 1|AB_1 1|D3|1  2.067833848e-12
L1|D3|2 1|D3|1 1|D3|4  2.067833848e-12
L1|D3|3 1|D3|4 1|D3|6  2.067833848e-12
L1|D3|4 1|D3|6 1|AB  2.067833848e-12
L1|D3|P1 1|D3|2 0  2e-13
L1|D3|P2 1|D3|7 0  2e-13
L1|D3|B1 1|D3|5 1|D3|4  2e-12
R1|D3|B1 1|D3|1 1|D3|3  2.7439617672
R1|D3|B2 1|D3|6 1|D3|8  2.7439617672
L1|D3|RB1 1|D3|3 0  1.750338398468e-12
L1|D3|RB2 1|D3|8 0  1.750338398468e-12
B1|D4|1 1|D4|1 1|D4|2 JJMIT AREA=2.5
B1|D4|2 1|D4|6 1|D4|7 JJMIT AREA=2.5
I1|D4|B1 0 1|D4|5  0.00035
L1|D4|1 1|CD_1 1|D4|1  2.067833848e-12
L1|D4|2 1|D4|1 1|D4|4  2.067833848e-12
L1|D4|3 1|D4|4 1|D4|6  2.067833848e-12
L1|D4|4 1|D4|6 1|CD  2.067833848e-12
L1|D4|P1 1|D4|2 0  2e-13
L1|D4|P2 1|D4|7 0  2e-13
L1|D4|B1 1|D4|5 1|D4|4  2e-12
R1|D4|B1 1|D4|1 1|D4|3  2.7439617672
R1|D4|B2 1|D4|6 1|D4|8  2.7439617672
L1|D4|RB1 1|D4|3 0  1.750338398468e-12
L1|D4|RB2 1|D4|8 0  1.750338398468e-12
I1|_AB_SPL|B1 0 1|_AB_SPL|3  PWL(0 0 5e-12 0.000175)
I1|_AB_SPL|B2 0 1|_AB_SPL|6  PWL(0 0 5e-12 0.000245)
I1|_AB_SPL|B3 0 1|_AB_SPL|10  PWL(0 0 5e-12 0.000175)
I1|_AB_SPL|B4 0 1|_AB_SPL|13  PWL(0 0 5e-12 0.000175)
L1|_AB_SPL|B1 1|_AB_SPL|3 1|_AB_SPL|1  2e-12
L1|_AB_SPL|B2 1|_AB_SPL|6 1|_AB_SPL|4  2e-12
L1|_AB_SPL|B3 1|_AB_SPL|10 1|_AB_SPL|8  2e-12
L1|_AB_SPL|B4 1|_AB_SPL|13 1|_AB_SPL|11  2e-12
B1|_AB_SPL|1 1|_AB_SPL|1 1|_AB_SPL|2 JJMIT AREA=2.5
B1|_AB_SPL|2 1|_AB_SPL|4 1|_AB_SPL|5 JJMIT AREA=3.5
B1|_AB_SPL|3 1|_AB_SPL|8 1|_AB_SPL|9 JJMIT AREA=2.5
B1|_AB_SPL|4 1|_AB_SPL|11 1|_AB_SPL|12 JJMIT AREA=2.5
L1|_AB_SPL|1 1|AB 1|_AB_SPL|1  2e-12
L1|_AB_SPL|2 1|_AB_SPL|1 1|_AB_SPL|4  4.135667696e-12
L1|_AB_SPL|3 1|_AB_SPL|4 1|_AB_SPL|7  1.4770241771428573e-12
L1|_AB_SPL|4 1|_AB_SPL|7 1|_AB_SPL|8  1.4770241771428573e-12
L1|_AB_SPL|5 1|_AB_SPL|8 1|ABX  2e-12
L1|_AB_SPL|6 1|_AB_SPL|7 1|_AB_SPL|11  1.4770241771428573e-12
L1|_AB_SPL|7 1|_AB_SPL|11 1|ABN  2e-12
L1|_AB_SPL|P1 1|_AB_SPL|2 0  2e-13
L1|_AB_SPL|P2 1|_AB_SPL|5 0  2e-13
L1|_AB_SPL|P3 1|_AB_SPL|9 0  2e-13
L1|_AB_SPL|P4 1|_AB_SPL|12 0  2e-13
R1|_AB_SPL|B1 1|_AB_SPL|1 1|_AB_SPL|101  2.7439617672
L1|_AB_SPL|RB1 1|_AB_SPL|101 0  1.550338398468e-12
R1|_AB_SPL|B2 1|_AB_SPL|4 1|_AB_SPL|104  1.9599726908571429
L1|_AB_SPL|RB2 1|_AB_SPL|104 0  1.1073845703342858e-12
R1|_AB_SPL|B3 1|_AB_SPL|8 1|_AB_SPL|108  2.7439617672
L1|_AB_SPL|RB3 1|_AB_SPL|108 0  1.550338398468e-12
R1|_AB_SPL|B4 1|_AB_SPL|11 1|_AB_SPL|111  2.7439617672
L1|_AB_SPL|RB4 1|_AB_SPL|111 0  1.550338398468e-12
L1|_XOR|A1 1|ABX 1|_XOR|A1  2.067833848e-12
L1|_XOR|A2 1|_XOR|A1 1|_XOR|A2  4.135667696e-12
L1|_XOR|A3 1|_XOR|A3 1|_XOR|AB  8.271335392e-12
L1|_XOR|B1 1|CD 1|_XOR|B1  2.067833848e-12
L1|_XOR|B2 1|_XOR|B1 1|_XOR|B2  4.135667696e-12
L1|_XOR|B3 1|_XOR|B3 1|_XOR|AB  8.271335392e-12
L1|_XOR|T1 T2 1|_XOR|T1  2.067833848e-12
L1|_XOR|T2 1|_XOR|T1 1|_XOR|T2  4.135667696e-12
L1|_XOR|Q2 1|_XOR|ABTQ 1|_XOR|Q1  4.135667696e-12
L1|_XOR|Q1 1|_XOR|Q1 1|ABXCD  2.067833848e-12
B1|_NOT|1 1|_NOT|1 1|_NOT|2 JJMIT AREA=2.5
B1|_NOT|2 1|_NOT|4 1|_NOT|5 JJMIT AREA=2.5
B1|_NOT|3 1|_NOT|7 1|_NOT|8 JJMIT AREA=1.7857142857142858
B1|_NOT|4 1|_NOT|13 1|_NOT|14 JJMIT AREA=2.5
B1|_NOT|5 1|_NOT|17 1|_NOT|18 JJMIT AREA=1.7857142857142858
B1|_NOT|6 1|_NOT|10 1|_NOT|11 JJMIT AREA=2.5
B1|_NOT|7 1|_NOT|20 1|_NOT|18 JJMIT AREA=1.7857142857142858
B1|_NOT|8 1|_NOT|18 1|_NOT|19 JJMIT AREA=2.5
B1|_NOT|9 1|_NOT|21 1|_NOT|22 JJMIT AREA=2.5
I1|_NOT|B1 0 1|_NOT|3  0.00017499999999999997
I1|_NOT|B2 0 1|_NOT|6  0.000125
I1|_NOT|B3 0 1|_NOT|9  0.00017499999999999997
I1|_NOT|B4 0 1|_NOT|15  0.00017499999999999997
I1|_NOT|B5 0 1|_NOT|23  0.00017499999999999997
L1|_NOT|B1 1|_NOT|3 1|_NOT|1  2e-12
L1|_NOT|B2 1|_NOT|6 1|_NOT|4  2e-12
L1|_NOT|B3 1|_NOT|8 1|_NOT|9  2e-12
L1|_NOT|B4 1|_NOT|13 1|_NOT|15  2e-12
L1|_NOT|B5 1|_NOT|21 1|_NOT|23  2e-12
L1|_NOT|1 1|ABN 1|_NOT|1  2.067833848e-12
L1|_NOT|2 1|_NOT|1 1|_NOT|4  4.135667696e-12
L1|_NOT|3 1|_NOT|4 1|_NOT|7  4.135667696e-12
L1|_NOT|4 T2 1|_NOT|13  2.067833848e-12
L1|_NOT|5 1|_NOT|13 1|_NOT|16  1e-12
L1|_NOT|6 1|_NOT|16 1|_NOT|17  4.135667696e-12
L1|_NOT|7 1|_NOT|16 1|_NOT|12  2e-12
L1|_NOT|8 1|_NOT|10 1|_NOT|12  1e-12
L1|_NOT|9 1|_NOT|10 1|_NOT|8  8.271335392e-12
L1|_NOT|10 1|_NOT|8 1|_NOT|20  1e-12
L1|_NOT|11 1|_NOT|18 1|_NOT|21  4.135667696e-12
L1|_NOT|12 1|_NOT|21 1|NOT_AB  2.067833848e-12
L1|_NOT|P1 1|_NOT|2 0  2e-13
L1|_NOT|P2 1|_NOT|5 0  2e-13
L1|_NOT|P4 1|_NOT|14 0  2e-13
L1|_NOT|P6 1|_NOT|11 0  2e-13
L1|_NOT|P8 1|_NOT|19 0  2e-13
L1|_NOT|P9 1|_NOT|22 0  2e-13
R1|_NOT|B1 1|_NOT|1 1|_NOT|101  2.7439617672
L1|_NOT|RB1 1|_NOT|101 0  1.550338398468e-12
R1|_NOT|B2 1|_NOT|4 1|_NOT|104  2.7439617672
L1|_NOT|RB2 1|_NOT|104 1|_NOT|5  1.550338398468e-12
R1|_NOT|B3 1|_NOT|7 1|_NOT|107  3.84154647408
L1|_NOT|RB3 1|_NOT|107 1|_NOT|8  2.1704737578552e-12
R1|_NOT|B4 1|_NOT|13 1|_NOT|113  2.7439617672
L1|_NOT|RB4 1|_NOT|113 0  1.550338398468e-12
R1|_NOT|B5 1|_NOT|17 1|_NOT|117  3.84154647408
L1|_NOT|RB5 1|_NOT|117 1|_NOT|18  2.1704737578552e-12
R1|_NOT|B6 1|_NOT|10 1|_NOT|110  2.7439617672
L1|_NOT|RB6 1|_NOT|110 0  1.550338398468e-12
R1|_NOT|B7 1|_NOT|20 1|_NOT|120  3.84154647408
L1|_NOT|RB7 1|_NOT|120 1|_NOT|18  2.1704737578552e-12
R1|_NOT|B8 1|_NOT|18 1|_NOT|118  2.7439617672
L1|_NOT|RB8 1|_NOT|118 0  1.550338398468e-12
R1|_NOT|B9 1|_NOT|21 1|_NOT|121  2.7439617672
L1|_NOT|RB9 1|_NOT|121 0  1.550338398468e-12
L1|_NOT|RD 1|_NOT|12 1|_NOT|112  2e-12
R1|_NOT|D 1|_NOT|112 0  4
L1|JTLOUT1|1 1|ABXCD 1|JTLOUT1|1  2.067833848e-12
L1|JTLOUT1|2 1|JTLOUT1|1 1|JTLOUT1|4  2.067833848e-12
L1|JTLOUT1|3 1|JTLOUT1|4 1|JTLOUT1|6  2.067833848e-12
L1|JTLOUT1|4 1|JTLOUT1|6 AB_XOR_CD_1  2.067833848e-12
L1|JTLOUT2|1 1|NOT_AB 1|JTLOUT2|1  2.067833848e-12
L1|JTLOUT2|2 1|JTLOUT2|1 1|JTLOUT2|4  2.067833848e-12
L1|JTLOUT2|3 1|JTLOUT2|4 1|JTLOUT2|6  2.067833848e-12
L1|JTLOUT2|4 1|JTLOUT2|6 NOT_AB_1  2.067833848e-12
L1|_AND_AB|I_1|B 1|_AND_AB|A1 1|_AND_AB|I_1|MID  2e-12
I1|_AND_AB|I_1|B 0 1|_AND_AB|I_1|MID  0.000175
L1|_AND_AB|I_5|B 1|_AND_AB|A3 1|_AND_AB|I_5|MID  2e-12
I1|_AND_AB|I_5|B 0 1|_AND_AB|I_5|MID  0.000175
L1|_AND_AB|I_14|B 1|_AND_AB|B1 1|_AND_AB|I_14|MID  2e-12
I1|_AND_AB|I_14|B 0 1|_AND_AB|I_14|MID  0.000175
L1|_AND_AB|I_18|B 1|_AND_AB|B3 1|_AND_AB|I_18|MID  2e-12
I1|_AND_AB|I_18|B 0 1|_AND_AB|I_18|MID  0.000175
L1|_AND_AB|I_25|B 1|_AND_AB|T1 1|_AND_AB|I_25|MID  2e-12
I1|_AND_AB|I_25|B 0 1|_AND_AB|I_25|MID  0.000175
L1|_AND_AB|I_28|B 1|_AND_AB|Q1 1|_AND_AB|I_28|MID  2e-12
I1|_AND_AB|I_28|B 0 1|_AND_AB|I_28|MID  0.000175
L1|_AND_AB|I_31|B 1|_AND_AB|T2 1|_AND_AB|I_31|MID  2e-12
I1|_AND_AB|I_31|B 0 1|_AND_AB|I_31|MID  0.000175
B1|_AND_AB|B1|1 1|_AND_AB|A1 1|_AND_AB|B1|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B1|P 1|_AND_AB|B1|MID_SERIES 0  2e-13
R1|_AND_AB|B1|B 1|_AND_AB|A1 1|_AND_AB|B1|MID_SHUNT  2.7439617672
L1|_AND_AB|B1|RB 1|_AND_AB|B1|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B2|1 1|_AND_AB|A2 1|_AND_AB|A3 JJMIT AREA=1.7857142857142858
R1|_AND_AB|B2|B 1|_AND_AB|A2 1|_AND_AB|B2|MID_SHUNT  3.84154647408
L1|_AND_AB|B2|RB 1|_AND_AB|B2|MID_SHUNT 1|_AND_AB|A3  2.1704737578552e-12
B1|_AND_AB|B3|1 1|_AND_AB|A3 1|_AND_AB|B3|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B3|P 1|_AND_AB|B3|MID_SERIES 0  2e-13
R1|_AND_AB|B3|B 1|_AND_AB|A3 1|_AND_AB|B3|MID_SHUNT  2.7439617672
L1|_AND_AB|B3|RB 1|_AND_AB|B3|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B4|1 1|_AND_AB|A4 1|_AND_AB|TA JJMIT AREA=1.7857142857142858
R1|_AND_AB|B4|B 1|_AND_AB|A4 1|_AND_AB|B4|MID_SHUNT  3.84154647408
L1|_AND_AB|B4|RB 1|_AND_AB|B4|MID_SHUNT 1|_AND_AB|TA  2.1704737578552e-12
B1|_AND_AB|B5|1 1|_AND_AB|A4 1|_AND_AB|B5|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B5|P 1|_AND_AB|B5|MID_SERIES 0  2e-13
R1|_AND_AB|B5|B 1|_AND_AB|A4 1|_AND_AB|B5|MID_SHUNT  2.7439617672
L1|_AND_AB|B5|RB 1|_AND_AB|B5|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B6|1 1|_AND_AB|A5 1|_AND_AB|Q2 JJMIT AREA=1.7857142857142858
R1|_AND_AB|B6|B 1|_AND_AB|A5 1|_AND_AB|B6|MID_SHUNT  3.84154647408
L1|_AND_AB|B6|RB 1|_AND_AB|B6|MID_SHUNT 1|_AND_AB|Q2  2.1704737578552e-12
B1|_AND_AB|B7|1 1|_AND_AB|B1 1|_AND_AB|B7|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B7|P 1|_AND_AB|B7|MID_SERIES 0  2e-13
R1|_AND_AB|B7|B 1|_AND_AB|B1 1|_AND_AB|B7|MID_SHUNT  2.7439617672
L1|_AND_AB|B7|RB 1|_AND_AB|B7|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B8|1 1|_AND_AB|B2 1|_AND_AB|B3 JJMIT AREA=1.7857142857142858
R1|_AND_AB|B8|B 1|_AND_AB|B2 1|_AND_AB|B8|MID_SHUNT  3.84154647408
L1|_AND_AB|B8|RB 1|_AND_AB|B8|MID_SHUNT 1|_AND_AB|B3  2.1704737578552e-12
B1|_AND_AB|B9|1 1|_AND_AB|B3 1|_AND_AB|B9|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B9|P 1|_AND_AB|B9|MID_SERIES 0  2e-13
R1|_AND_AB|B9|B 1|_AND_AB|B3 1|_AND_AB|B9|MID_SHUNT  2.7439617672
L1|_AND_AB|B9|RB 1|_AND_AB|B9|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B10|1 1|_AND_AB|B4 1|_AND_AB|TB JJMIT AREA=1.7857142857142858
R1|_AND_AB|B10|B 1|_AND_AB|B4 1|_AND_AB|B10|MID_SHUNT  3.84154647408
L1|_AND_AB|B10|RB 1|_AND_AB|B10|MID_SHUNT 1|_AND_AB|TB  2.1704737578552e-12
B1|_AND_AB|B11|1 1|_AND_AB|B4 1|_AND_AB|B11|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B11|P 1|_AND_AB|B11|MID_SERIES 0  2e-13
R1|_AND_AB|B11|B 1|_AND_AB|B4 1|_AND_AB|B11|MID_SHUNT  2.7439617672
L1|_AND_AB|B11|RB 1|_AND_AB|B11|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B12|1 1|_AND_AB|B5 1|_AND_AB|Q2 JJMIT AREA=1.7857142857142858
R1|_AND_AB|B12|B 1|_AND_AB|B5 1|_AND_AB|B12|MID_SHUNT  3.84154647408
L1|_AND_AB|B12|RB 1|_AND_AB|B12|MID_SHUNT 1|_AND_AB|Q2  2.1704737578552e-12
B1|_AND_AB|B13|1 1|_AND_AB|T1 1|_AND_AB|B13|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B13|P 1|_AND_AB|B13|MID_SERIES 0  2e-13
R1|_AND_AB|B13|B 1|_AND_AB|T1 1|_AND_AB|B13|MID_SHUNT  2.7439617672
L1|_AND_AB|B13|RB 1|_AND_AB|B13|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B14|1 1|_AND_AB|T2 1|_AND_AB|B14|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B14|P 1|_AND_AB|B14|MID_SERIES 0  2e-13
R1|_AND_AB|B14|B 1|_AND_AB|T2 1|_AND_AB|B14|MID_SHUNT  2.7439617672
L1|_AND_AB|B14|RB 1|_AND_AB|B14|MID_SHUNT 0  1.550338398468e-12
B1|_AND_AB|B15|1 1|_AND_AB|Q1 1|_AND_AB|B15|MID_SERIES JJMIT AREA=2.5
L1|_AND_AB|B15|P 1|_AND_AB|B15|MID_SERIES 0  2e-13
R1|_AND_AB|B15|B 1|_AND_AB|Q1 1|_AND_AB|B15|MID_SHUNT  2.7439617672
L1|_AND_AB|B15|RB 1|_AND_AB|B15|MID_SHUNT 0  1.550338398468e-12
L1|_AND_CD|I_1|B 1|_AND_CD|A1 1|_AND_CD|I_1|MID  2e-12
I1|_AND_CD|I_1|B 0 1|_AND_CD|I_1|MID  0.000175
L1|_AND_CD|I_5|B 1|_AND_CD|A3 1|_AND_CD|I_5|MID  2e-12
I1|_AND_CD|I_5|B 0 1|_AND_CD|I_5|MID  0.000175
L1|_AND_CD|I_14|B 1|_AND_CD|B1 1|_AND_CD|I_14|MID  2e-12
I1|_AND_CD|I_14|B 0 1|_AND_CD|I_14|MID  0.000175
L1|_AND_CD|I_18|B 1|_AND_CD|B3 1|_AND_CD|I_18|MID  2e-12
I1|_AND_CD|I_18|B 0 1|_AND_CD|I_18|MID  0.000175
L1|_AND_CD|I_25|B 1|_AND_CD|T1 1|_AND_CD|I_25|MID  2e-12
I1|_AND_CD|I_25|B 0 1|_AND_CD|I_25|MID  0.000175
L1|_AND_CD|I_28|B 1|_AND_CD|Q1 1|_AND_CD|I_28|MID  2e-12
I1|_AND_CD|I_28|B 0 1|_AND_CD|I_28|MID  0.000175
L1|_AND_CD|I_31|B 1|_AND_CD|T2 1|_AND_CD|I_31|MID  2e-12
I1|_AND_CD|I_31|B 0 1|_AND_CD|I_31|MID  0.000175
B1|_AND_CD|B1|1 1|_AND_CD|A1 1|_AND_CD|B1|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B1|P 1|_AND_CD|B1|MID_SERIES 0  2e-13
R1|_AND_CD|B1|B 1|_AND_CD|A1 1|_AND_CD|B1|MID_SHUNT  2.7439617672
L1|_AND_CD|B1|RB 1|_AND_CD|B1|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B2|1 1|_AND_CD|A2 1|_AND_CD|A3 JJMIT AREA=1.7857142857142858
R1|_AND_CD|B2|B 1|_AND_CD|A2 1|_AND_CD|B2|MID_SHUNT  3.84154647408
L1|_AND_CD|B2|RB 1|_AND_CD|B2|MID_SHUNT 1|_AND_CD|A3  2.1704737578552e-12
B1|_AND_CD|B3|1 1|_AND_CD|A3 1|_AND_CD|B3|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B3|P 1|_AND_CD|B3|MID_SERIES 0  2e-13
R1|_AND_CD|B3|B 1|_AND_CD|A3 1|_AND_CD|B3|MID_SHUNT  2.7439617672
L1|_AND_CD|B3|RB 1|_AND_CD|B3|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B4|1 1|_AND_CD|A4 1|_AND_CD|TA JJMIT AREA=1.7857142857142858
R1|_AND_CD|B4|B 1|_AND_CD|A4 1|_AND_CD|B4|MID_SHUNT  3.84154647408
L1|_AND_CD|B4|RB 1|_AND_CD|B4|MID_SHUNT 1|_AND_CD|TA  2.1704737578552e-12
B1|_AND_CD|B5|1 1|_AND_CD|A4 1|_AND_CD|B5|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B5|P 1|_AND_CD|B5|MID_SERIES 0  2e-13
R1|_AND_CD|B5|B 1|_AND_CD|A4 1|_AND_CD|B5|MID_SHUNT  2.7439617672
L1|_AND_CD|B5|RB 1|_AND_CD|B5|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B6|1 1|_AND_CD|A5 1|_AND_CD|Q2 JJMIT AREA=1.7857142857142858
R1|_AND_CD|B6|B 1|_AND_CD|A5 1|_AND_CD|B6|MID_SHUNT  3.84154647408
L1|_AND_CD|B6|RB 1|_AND_CD|B6|MID_SHUNT 1|_AND_CD|Q2  2.1704737578552e-12
B1|_AND_CD|B7|1 1|_AND_CD|B1 1|_AND_CD|B7|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B7|P 1|_AND_CD|B7|MID_SERIES 0  2e-13
R1|_AND_CD|B7|B 1|_AND_CD|B1 1|_AND_CD|B7|MID_SHUNT  2.7439617672
L1|_AND_CD|B7|RB 1|_AND_CD|B7|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B8|1 1|_AND_CD|B2 1|_AND_CD|B3 JJMIT AREA=1.7857142857142858
R1|_AND_CD|B8|B 1|_AND_CD|B2 1|_AND_CD|B8|MID_SHUNT  3.84154647408
L1|_AND_CD|B8|RB 1|_AND_CD|B8|MID_SHUNT 1|_AND_CD|B3  2.1704737578552e-12
B1|_AND_CD|B9|1 1|_AND_CD|B3 1|_AND_CD|B9|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B9|P 1|_AND_CD|B9|MID_SERIES 0  2e-13
R1|_AND_CD|B9|B 1|_AND_CD|B3 1|_AND_CD|B9|MID_SHUNT  2.7439617672
L1|_AND_CD|B9|RB 1|_AND_CD|B9|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B10|1 1|_AND_CD|B4 1|_AND_CD|TB JJMIT AREA=1.7857142857142858
R1|_AND_CD|B10|B 1|_AND_CD|B4 1|_AND_CD|B10|MID_SHUNT  3.84154647408
L1|_AND_CD|B10|RB 1|_AND_CD|B10|MID_SHUNT 1|_AND_CD|TB  2.1704737578552e-12
B1|_AND_CD|B11|1 1|_AND_CD|B4 1|_AND_CD|B11|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B11|P 1|_AND_CD|B11|MID_SERIES 0  2e-13
R1|_AND_CD|B11|B 1|_AND_CD|B4 1|_AND_CD|B11|MID_SHUNT  2.7439617672
L1|_AND_CD|B11|RB 1|_AND_CD|B11|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B12|1 1|_AND_CD|B5 1|_AND_CD|Q2 JJMIT AREA=1.7857142857142858
R1|_AND_CD|B12|B 1|_AND_CD|B5 1|_AND_CD|B12|MID_SHUNT  3.84154647408
L1|_AND_CD|B12|RB 1|_AND_CD|B12|MID_SHUNT 1|_AND_CD|Q2  2.1704737578552e-12
B1|_AND_CD|B13|1 1|_AND_CD|T1 1|_AND_CD|B13|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B13|P 1|_AND_CD|B13|MID_SERIES 0  2e-13
R1|_AND_CD|B13|B 1|_AND_CD|T1 1|_AND_CD|B13|MID_SHUNT  2.7439617672
L1|_AND_CD|B13|RB 1|_AND_CD|B13|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B14|1 1|_AND_CD|T2 1|_AND_CD|B14|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B14|P 1|_AND_CD|B14|MID_SERIES 0  2e-13
R1|_AND_CD|B14|B 1|_AND_CD|T2 1|_AND_CD|B14|MID_SHUNT  2.7439617672
L1|_AND_CD|B14|RB 1|_AND_CD|B14|MID_SHUNT 0  1.550338398468e-12
B1|_AND_CD|B15|1 1|_AND_CD|Q1 1|_AND_CD|B15|MID_SERIES JJMIT AREA=2.5
L1|_AND_CD|B15|P 1|_AND_CD|B15|MID_SERIES 0  2e-13
R1|_AND_CD|B15|B 1|_AND_CD|Q1 1|_AND_CD|B15|MID_SHUNT  2.7439617672
L1|_AND_CD|B15|RB 1|_AND_CD|B15|MID_SHUNT 0  1.550338398468e-12
L1|_XOR|I_A1|B 1|_XOR|A1 1|_XOR|I_A1|MID  2e-12
I1|_XOR|I_A1|B 0 1|_XOR|I_A1|MID  0.000175
L1|_XOR|I_A3|B 1|_XOR|A3 1|_XOR|I_A3|MID  2e-12
I1|_XOR|I_A3|B 0 1|_XOR|I_A3|MID  0.000175
L1|_XOR|I_B1|B 1|_XOR|B1 1|_XOR|I_B1|MID  2e-12
I1|_XOR|I_B1|B 0 1|_XOR|I_B1|MID  0.000175
L1|_XOR|I_B3|B 1|_XOR|B3 1|_XOR|I_B3|MID  2e-12
I1|_XOR|I_B3|B 0 1|_XOR|I_B3|MID  0.000175
L1|_XOR|I_T1|B 1|_XOR|T1 1|_XOR|I_T1|MID  2e-12
I1|_XOR|I_T1|B 0 1|_XOR|I_T1|MID  0.000175
L1|_XOR|I_Q1|B 1|_XOR|Q1 1|_XOR|I_Q1|MID  2e-12
I1|_XOR|I_Q1|B 0 1|_XOR|I_Q1|MID  0.000175
B1|_XOR|A1|1 1|_XOR|A1 1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
L1|_XOR|A1|P 1|_XOR|A1|MID_SERIES 0  5e-13
R1|_XOR|A1|B 1|_XOR|A1 1|_XOR|A1|MID_SHUNT  2.7439617672
L1|_XOR|A1|RB 1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
B1|_XOR|A2|1 1|_XOR|A2 1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
L1|_XOR|A2|P 1|_XOR|A2|MID_SERIES 0  5e-13
R1|_XOR|A2|B 1|_XOR|A2 1|_XOR|A2|MID_SHUNT  2.7439617672
L1|_XOR|A2|RB 1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
B1|_XOR|A3|1 1|_XOR|A2 1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
L1|_XOR|A3|P 1|_XOR|A3|MID_SERIES 1|_XOR|A3  1.2e-12
R1|_XOR|A3|B 1|_XOR|A2 1|_XOR|A3|MID_SHUNT  2.7439617672
L1|_XOR|A3|RB 1|_XOR|A3|MID_SHUNT 1|_XOR|A3  2.050338398468e-12
B1|_XOR|B1|1 1|_XOR|B1 1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
L1|_XOR|B1|P 1|_XOR|B1|MID_SERIES 0  5e-13
R1|_XOR|B1|B 1|_XOR|B1 1|_XOR|B1|MID_SHUNT  2.7439617672
L1|_XOR|B1|RB 1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
B1|_XOR|B2|1 1|_XOR|B2 1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
L1|_XOR|B2|P 1|_XOR|B2|MID_SERIES 0  5e-13
R1|_XOR|B2|B 1|_XOR|B2 1|_XOR|B2|MID_SHUNT  2.7439617672
L1|_XOR|B2|RB 1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
B1|_XOR|B3|1 1|_XOR|B2 1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
L1|_XOR|B3|P 1|_XOR|B3|MID_SERIES 1|_XOR|B3  1.2e-12
R1|_XOR|B3|B 1|_XOR|B2 1|_XOR|B3|MID_SHUNT  2.7439617672
L1|_XOR|B3|RB 1|_XOR|B3|MID_SHUNT 1|_XOR|B3  2.050338398468e-12
B1|_XOR|T1|1 1|_XOR|T1 1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
L1|_XOR|T1|P 1|_XOR|T1|MID_SERIES 0  5e-13
R1|_XOR|T1|B 1|_XOR|T1 1|_XOR|T1|MID_SHUNT  2.7439617672
L1|_XOR|T1|RB 1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
B1|_XOR|T2|1 1|_XOR|T2 1|_XOR|ABTQ JJMIT AREA=2.5
R1|_XOR|T2|B 1|_XOR|T2 1|_XOR|T2|MID_SHUNT  2.7439617672
L1|_XOR|T2|RB 1|_XOR|T2|MID_SHUNT 1|_XOR|ABTQ  2.050338398468e-12
B1|_XOR|AB|1 1|_XOR|AB 1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
L1|_XOR|AB|P 1|_XOR|AB|MID_SERIES 1|_XOR|ABTQ  1.2e-12
R1|_XOR|AB|B 1|_XOR|AB 1|_XOR|AB|MID_SHUNT  3.429952209
L1|_XOR|AB|RB 1|_XOR|AB|MID_SHUNT 1|_XOR|ABTQ  2.437922998085e-12
B1|_XOR|ABTQ|1 1|_XOR|ABTQ 1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
L1|_XOR|ABTQ|P 1|_XOR|ABTQ|MID_SERIES 0  5e-13
R1|_XOR|ABTQ|B 1|_XOR|ABTQ 1|_XOR|ABTQ|MID_SHUNT  2.7439617672
L1|_XOR|ABTQ|RB 1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
B1|_XOR|Q1|1 1|_XOR|Q1 1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
L1|_XOR|Q1|P 1|_XOR|Q1|MID_SERIES 0  5e-13
R1|_XOR|Q1|B 1|_XOR|Q1 1|_XOR|Q1|MID_SHUNT  2.7439617672
L1|_XOR|Q1|RB 1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
B1|JTLOUT1|1|1 1|JTLOUT1|1 1|JTLOUT1|1|MID_SERIES JJMIT AREA=2.5
L1|JTLOUT1|1|P 1|JTLOUT1|1|MID_SERIES 0  2e-13
R1|JTLOUT1|1|B 1|JTLOUT1|1 1|JTLOUT1|1|MID_SHUNT  2.7439617672
L1|JTLOUT1|1|RB 1|JTLOUT1|1|MID_SHUNT 0  1.750338398468e-12
L1|JTLOUT1|B|B 1|JTLOUT1|4 1|JTLOUT1|B|MID  2e-12
I1|JTLOUT1|B|B 0 1|JTLOUT1|B|MID  0.0005
B1|JTLOUT1|2|1 1|JTLOUT1|6 1|JTLOUT1|2|MID_SERIES JJMIT AREA=2.5
L1|JTLOUT1|2|P 1|JTLOUT1|2|MID_SERIES 0  2e-13
R1|JTLOUT1|2|B 1|JTLOUT1|6 1|JTLOUT1|2|MID_SHUNT  2.7439617672
L1|JTLOUT1|2|RB 1|JTLOUT1|2|MID_SHUNT 0  1.750338398468e-12
B1|JTLOUT2|1|1 1|JTLOUT2|1 1|JTLOUT2|1|MID_SERIES JJMIT AREA=2.5
L1|JTLOUT2|1|P 1|JTLOUT2|1|MID_SERIES 0  2e-13
R1|JTLOUT2|1|B 1|JTLOUT2|1 1|JTLOUT2|1|MID_SHUNT  2.7439617672
L1|JTLOUT2|1|RB 1|JTLOUT2|1|MID_SHUNT 0  1.750338398468e-12
L1|JTLOUT2|B|B 1|JTLOUT2|4 1|JTLOUT2|B|MID  2e-12
I1|JTLOUT2|B|B 0 1|JTLOUT2|B|MID  0.0005
B1|JTLOUT2|2|1 1|JTLOUT2|6 1|JTLOUT2|2|MID_SERIES JJMIT AREA=2.5
L1|JTLOUT2|2|P 1|JTLOUT2|2|MID_SERIES 0  2e-13
R1|JTLOUT2|2|B 1|JTLOUT2|6 1|JTLOUT2|2|MID_SHUNT  2.7439617672
L1|JTLOUT2|2|RB 1|JTLOUT2|2|MID_SHUNT 0  1.750338398468e-12
.print DEVI ROUT1
.print DEVI ROUT2
.print DEVI IT1|T
.print DEVI IT2|T
.print DEVI IDATA_A1|A
.print DEVI IDATA_B1|B
.print DEVI IDATA_C1|T
.print DEVI IDATA_D1|T
.print DEVI L1|_AND_AB|1
.print DEVI L1|_AND_AB|2
.print DEVI L1|_AND_AB|3
.print DEVI L1|_AND_AB|4
.print DEVI L1|_AND_AB|5
.print DEVI L1|_AND_AB|6
.print DEVI L1|_AND_AB|7
.print DEVI L1|_AND_AB|8
.print DEVI L1|_AND_AB|9
.print DEVI L1|_AND_AB|10
.print DEVI L1|_AND_AB|11
.print DEVI L1|_AND_AB|12
.print DEVI L1|_AND_AB|13
.print DEVI L1|_AND_AB|14
.print DEVI L1|_AND_AB|15
.print DEVI L1|_AND_CD|1
.print DEVI L1|_AND_CD|2
.print DEVI L1|_AND_CD|3
.print DEVI L1|_AND_CD|4
.print DEVI L1|_AND_CD|5
.print DEVI L1|_AND_CD|6
.print DEVI L1|_AND_CD|7
.print DEVI L1|_AND_CD|8
.print DEVI L1|_AND_CD|9
.print DEVI L1|_AND_CD|10
.print DEVI L1|_AND_CD|11
.print DEVI L1|_AND_CD|12
.print DEVI L1|_AND_CD|13
.print DEVI L1|_AND_CD|14
.print DEVI L1|_AND_CD|15
.print DEVI B1|D1|1
.print DEVI B1|D1|2
.print DEVI B1|D1|3
.print DEVI B1|D1|4
.print DEVI I1|D1|B1
.print DEVI I1|D1|B2
.print DEVI I1|D1|B3
.print DEVI I1|D1|B4
.print DEVI L1|D1|1
.print DEVI L1|D1|2
.print DEVI L1|D1|3
.print DEVI L1|D1|4
.print DEVI L1|D1|5
.print DEVI L1|D1|P1
.print DEVI L1|D1|P2
.print DEVI L1|D1|P3
.print DEVI L1|D1|P4
.print DEVI L1|D1|B1
.print DEVI L1|D1|B2
.print DEVI L1|D1|B3
.print DEVI L1|D1|B4
.print DEVI R1|D1|B1
.print DEVI R1|D1|B2
.print DEVI R1|D1|B3
.print DEVI R1|D1|B4
.print DEVI L1|D1|RB1
.print DEVI L1|D1|RB2
.print DEVI L1|D1|RB3
.print DEVI L1|D1|RB4
.print DEVI B1|D2|1
.print DEVI B1|D2|2
.print DEVI B1|D2|3
.print DEVI B1|D2|4
.print DEVI I1|D2|B1
.print DEVI I1|D2|B2
.print DEVI I1|D2|B3
.print DEVI I1|D2|B4
.print DEVI L1|D2|1
.print DEVI L1|D2|2
.print DEVI L1|D2|3
.print DEVI L1|D2|4
.print DEVI L1|D2|5
.print DEVI L1|D2|P1
.print DEVI L1|D2|P2
.print DEVI L1|D2|P3
.print DEVI L1|D2|P4
.print DEVI L1|D2|B1
.print DEVI L1|D2|B2
.print DEVI L1|D2|B3
.print DEVI L1|D2|B4
.print DEVI R1|D2|B1
.print DEVI R1|D2|B2
.print DEVI R1|D2|B3
.print DEVI R1|D2|B4
.print DEVI L1|D2|RB1
.print DEVI L1|D2|RB2
.print DEVI L1|D2|RB3
.print DEVI L1|D2|RB4
.print DEVI B1|D3|1
.print DEVI B1|D3|2
.print DEVI I1|D3|B1
.print DEVI L1|D3|1
.print DEVI L1|D3|2
.print DEVI L1|D3|3
.print DEVI L1|D3|4
.print DEVI L1|D3|P1
.print DEVI L1|D3|P2
.print DEVI L1|D3|B1
.print DEVI R1|D3|B1
.print DEVI R1|D3|B2
.print DEVI L1|D3|RB1
.print DEVI L1|D3|RB2
.print DEVI B1|D4|1
.print DEVI B1|D4|2
.print DEVI I1|D4|B1
.print DEVI L1|D4|1
.print DEVI L1|D4|2
.print DEVI L1|D4|3
.print DEVI L1|D4|4
.print DEVI L1|D4|P1
.print DEVI L1|D4|P2
.print DEVI L1|D4|B1
.print DEVI R1|D4|B1
.print DEVI R1|D4|B2
.print DEVI L1|D4|RB1
.print DEVI L1|D4|RB2
.print DEVI I1|_AB_SPL|B1
.print DEVI I1|_AB_SPL|B2
.print DEVI I1|_AB_SPL|B3
.print DEVI I1|_AB_SPL|B4
.print DEVI L1|_AB_SPL|B1
.print DEVI L1|_AB_SPL|B2
.print DEVI L1|_AB_SPL|B3
.print DEVI L1|_AB_SPL|B4
.print DEVI B1|_AB_SPL|1
.print DEVI B1|_AB_SPL|2
.print DEVI B1|_AB_SPL|3
.print DEVI B1|_AB_SPL|4
.print DEVI L1|_AB_SPL|1
.print DEVI L1|_AB_SPL|2
.print DEVI L1|_AB_SPL|3
.print DEVI L1|_AB_SPL|4
.print DEVI L1|_AB_SPL|5
.print DEVI L1|_AB_SPL|6
.print DEVI L1|_AB_SPL|7
.print DEVI L1|_AB_SPL|P1
.print DEVI L1|_AB_SPL|P2
.print DEVI L1|_AB_SPL|P3
.print DEVI L1|_AB_SPL|P4
.print DEVI R1|_AB_SPL|B1
.print DEVI L1|_AB_SPL|RB1
.print DEVI R1|_AB_SPL|B2
.print DEVI L1|_AB_SPL|RB2
.print DEVI R1|_AB_SPL|B3
.print DEVI L1|_AB_SPL|RB3
.print DEVI R1|_AB_SPL|B4
.print DEVI L1|_AB_SPL|RB4
.print DEVI L1|_XOR|A1
.print DEVI L1|_XOR|A2
.print DEVI L1|_XOR|A3
.print DEVI L1|_XOR|B1
.print DEVI L1|_XOR|B2
.print DEVI L1|_XOR|B3
.print DEVI L1|_XOR|T1
.print DEVI L1|_XOR|T2
.print DEVI L1|_XOR|Q2
.print DEVI L1|_XOR|Q1
.print DEVI B1|_NOT|1
.print DEVI B1|_NOT|2
.print DEVI B1|_NOT|3
.print DEVI B1|_NOT|4
.print DEVI B1|_NOT|5
.print DEVI B1|_NOT|6
.print DEVI B1|_NOT|7
.print DEVI B1|_NOT|8
.print DEVI B1|_NOT|9
.print DEVI I1|_NOT|B1
.print DEVI I1|_NOT|B2
.print DEVI I1|_NOT|B3
.print DEVI I1|_NOT|B4
.print DEVI I1|_NOT|B5
.print DEVI L1|_NOT|B1
.print DEVI L1|_NOT|B2
.print DEVI L1|_NOT|B3
.print DEVI L1|_NOT|B4
.print DEVI L1|_NOT|B5
.print DEVI L1|_NOT|1
.print DEVI L1|_NOT|2
.print DEVI L1|_NOT|3
.print DEVI L1|_NOT|4
.print DEVI L1|_NOT|5
.print DEVI L1|_NOT|6
.print DEVI L1|_NOT|7
.print DEVI L1|_NOT|8
.print DEVI L1|_NOT|9
.print DEVI L1|_NOT|10
.print DEVI L1|_NOT|11
.print DEVI L1|_NOT|12
.print DEVI L1|_NOT|P1
.print DEVI L1|_NOT|P2
.print DEVI L1|_NOT|P4
.print DEVI L1|_NOT|P6
.print DEVI L1|_NOT|P8
.print DEVI L1|_NOT|P9
.print DEVI R1|_NOT|B1
.print DEVI L1|_NOT|RB1
.print DEVI R1|_NOT|B2
.print DEVI L1|_NOT|RB2
.print DEVI R1|_NOT|B3
.print DEVI L1|_NOT|RB3
.print DEVI R1|_NOT|B4
.print DEVI L1|_NOT|RB4
.print DEVI R1|_NOT|B5
.print DEVI L1|_NOT|RB5
.print DEVI R1|_NOT|B6
.print DEVI L1|_NOT|RB6
.print DEVI R1|_NOT|B7
.print DEVI L1|_NOT|RB7
.print DEVI R1|_NOT|B8
.print DEVI L1|_NOT|RB8
.print DEVI R1|_NOT|B9
.print DEVI L1|_NOT|RB9
.print DEVI L1|_NOT|RD
.print DEVI R1|_NOT|D
.print DEVI L1|JTLOUT1|1
.print DEVI L1|JTLOUT1|2
.print DEVI L1|JTLOUT1|3
.print DEVI L1|JTLOUT1|4
.print DEVI L1|JTLOUT2|1
.print DEVI L1|JTLOUT2|2
.print DEVI L1|JTLOUT2|3
.print DEVI L1|JTLOUT2|4
.print DEVI L1|_AND_AB|I_1|B
.print DEVI I1|_AND_AB|I_1|B
.print DEVI L1|_AND_AB|I_5|B
.print DEVI I1|_AND_AB|I_5|B
.print DEVI L1|_AND_AB|I_14|B
.print DEVI I1|_AND_AB|I_14|B
.print DEVI L1|_AND_AB|I_18|B
.print DEVI I1|_AND_AB|I_18|B
.print DEVI L1|_AND_AB|I_25|B
.print DEVI I1|_AND_AB|I_25|B
.print DEVI L1|_AND_AB|I_28|B
.print DEVI I1|_AND_AB|I_28|B
.print DEVI L1|_AND_AB|I_31|B
.print DEVI I1|_AND_AB|I_31|B
.print DEVI B1|_AND_AB|B1|1
.print DEVI L1|_AND_AB|B1|P
.print DEVI R1|_AND_AB|B1|B
.print DEVI L1|_AND_AB|B1|RB
.print DEVI B1|_AND_AB|B2|1
.print DEVI R1|_AND_AB|B2|B
.print DEVI L1|_AND_AB|B2|RB
.print DEVI B1|_AND_AB|B3|1
.print DEVI L1|_AND_AB|B3|P
.print DEVI R1|_AND_AB|B3|B
.print DEVI L1|_AND_AB|B3|RB
.print DEVI B1|_AND_AB|B4|1
.print DEVI R1|_AND_AB|B4|B
.print DEVI L1|_AND_AB|B4|RB
.print DEVI B1|_AND_AB|B5|1
.print DEVI L1|_AND_AB|B5|P
.print DEVI R1|_AND_AB|B5|B
.print DEVI L1|_AND_AB|B5|RB
.print DEVI B1|_AND_AB|B6|1
.print DEVI R1|_AND_AB|B6|B
.print DEVI L1|_AND_AB|B6|RB
.print DEVI B1|_AND_AB|B7|1
.print DEVI L1|_AND_AB|B7|P
.print DEVI R1|_AND_AB|B7|B
.print DEVI L1|_AND_AB|B7|RB
.print DEVI B1|_AND_AB|B8|1
.print DEVI R1|_AND_AB|B8|B
.print DEVI L1|_AND_AB|B8|RB
.print DEVI B1|_AND_AB|B9|1
.print DEVI L1|_AND_AB|B9|P
.print DEVI R1|_AND_AB|B9|B
.print DEVI L1|_AND_AB|B9|RB
.print DEVI B1|_AND_AB|B10|1
.print DEVI R1|_AND_AB|B10|B
.print DEVI L1|_AND_AB|B10|RB
.print DEVI B1|_AND_AB|B11|1
.print DEVI L1|_AND_AB|B11|P
.print DEVI R1|_AND_AB|B11|B
.print DEVI L1|_AND_AB|B11|RB
.print DEVI B1|_AND_AB|B12|1
.print DEVI R1|_AND_AB|B12|B
.print DEVI L1|_AND_AB|B12|RB
.print DEVI B1|_AND_AB|B13|1
.print DEVI L1|_AND_AB|B13|P
.print DEVI R1|_AND_AB|B13|B
.print DEVI L1|_AND_AB|B13|RB
.print DEVI B1|_AND_AB|B14|1
.print DEVI L1|_AND_AB|B14|P
.print DEVI R1|_AND_AB|B14|B
.print DEVI L1|_AND_AB|B14|RB
.print DEVI B1|_AND_AB|B15|1
.print DEVI L1|_AND_AB|B15|P
.print DEVI R1|_AND_AB|B15|B
.print DEVI L1|_AND_AB|B15|RB
.print DEVI L1|_AND_CD|I_1|B
.print DEVI I1|_AND_CD|I_1|B
.print DEVI L1|_AND_CD|I_5|B
.print DEVI I1|_AND_CD|I_5|B
.print DEVI L1|_AND_CD|I_14|B
.print DEVI I1|_AND_CD|I_14|B
.print DEVI L1|_AND_CD|I_18|B
.print DEVI I1|_AND_CD|I_18|B
.print DEVI L1|_AND_CD|I_25|B
.print DEVI I1|_AND_CD|I_25|B
.print DEVI L1|_AND_CD|I_28|B
.print DEVI I1|_AND_CD|I_28|B
.print DEVI L1|_AND_CD|I_31|B
.print DEVI I1|_AND_CD|I_31|B
.print DEVI B1|_AND_CD|B1|1
.print DEVI L1|_AND_CD|B1|P
.print DEVI R1|_AND_CD|B1|B
.print DEVI L1|_AND_CD|B1|RB
.print DEVI B1|_AND_CD|B2|1
.print DEVI R1|_AND_CD|B2|B
.print DEVI L1|_AND_CD|B2|RB
.print DEVI B1|_AND_CD|B3|1
.print DEVI L1|_AND_CD|B3|P
.print DEVI R1|_AND_CD|B3|B
.print DEVI L1|_AND_CD|B3|RB
.print DEVI B1|_AND_CD|B4|1
.print DEVI R1|_AND_CD|B4|B
.print DEVI L1|_AND_CD|B4|RB
.print DEVI B1|_AND_CD|B5|1
.print DEVI L1|_AND_CD|B5|P
.print DEVI R1|_AND_CD|B5|B
.print DEVI L1|_AND_CD|B5|RB
.print DEVI B1|_AND_CD|B6|1
.print DEVI R1|_AND_CD|B6|B
.print DEVI L1|_AND_CD|B6|RB
.print DEVI B1|_AND_CD|B7|1
.print DEVI L1|_AND_CD|B7|P
.print DEVI R1|_AND_CD|B7|B
.print DEVI L1|_AND_CD|B7|RB
.print DEVI B1|_AND_CD|B8|1
.print DEVI R1|_AND_CD|B8|B
.print DEVI L1|_AND_CD|B8|RB
.print DEVI B1|_AND_CD|B9|1
.print DEVI L1|_AND_CD|B9|P
.print DEVI R1|_AND_CD|B9|B
.print DEVI L1|_AND_CD|B9|RB
.print DEVI B1|_AND_CD|B10|1
.print DEVI R1|_AND_CD|B10|B
.print DEVI L1|_AND_CD|B10|RB
.print DEVI B1|_AND_CD|B11|1
.print DEVI L1|_AND_CD|B11|P
.print DEVI R1|_AND_CD|B11|B
.print DEVI L1|_AND_CD|B11|RB
.print DEVI B1|_AND_CD|B12|1
.print DEVI R1|_AND_CD|B12|B
.print DEVI L1|_AND_CD|B12|RB
.print DEVI B1|_AND_CD|B13|1
.print DEVI L1|_AND_CD|B13|P
.print DEVI R1|_AND_CD|B13|B
.print DEVI L1|_AND_CD|B13|RB
.print DEVI B1|_AND_CD|B14|1
.print DEVI L1|_AND_CD|B14|P
.print DEVI R1|_AND_CD|B14|B
.print DEVI L1|_AND_CD|B14|RB
.print DEVI B1|_AND_CD|B15|1
.print DEVI L1|_AND_CD|B15|P
.print DEVI R1|_AND_CD|B15|B
.print DEVI L1|_AND_CD|B15|RB
.print DEVI L1|_XOR|I_A1|B
.print DEVI I1|_XOR|I_A1|B
.print DEVI L1|_XOR|I_A3|B
.print DEVI I1|_XOR|I_A3|B
.print DEVI L1|_XOR|I_B1|B
.print DEVI I1|_XOR|I_B1|B
.print DEVI L1|_XOR|I_B3|B
.print DEVI I1|_XOR|I_B3|B
.print DEVI L1|_XOR|I_T1|B
.print DEVI I1|_XOR|I_T1|B
.print DEVI L1|_XOR|I_Q1|B
.print DEVI I1|_XOR|I_Q1|B
.print DEVI B1|_XOR|A1|1
.print DEVI L1|_XOR|A1|P
.print DEVI R1|_XOR|A1|B
.print DEVI L1|_XOR|A1|RB
.print DEVI B1|_XOR|A2|1
.print DEVI L1|_XOR|A2|P
.print DEVI R1|_XOR|A2|B
.print DEVI L1|_XOR|A2|RB
.print DEVI B1|_XOR|A3|1
.print DEVI L1|_XOR|A3|P
.print DEVI R1|_XOR|A3|B
.print DEVI L1|_XOR|A3|RB
.print DEVI B1|_XOR|B1|1
.print DEVI L1|_XOR|B1|P
.print DEVI R1|_XOR|B1|B
.print DEVI L1|_XOR|B1|RB
.print DEVI B1|_XOR|B2|1
.print DEVI L1|_XOR|B2|P
.print DEVI R1|_XOR|B2|B
.print DEVI L1|_XOR|B2|RB
.print DEVI B1|_XOR|B3|1
.print DEVI L1|_XOR|B3|P
.print DEVI R1|_XOR|B3|B
.print DEVI L1|_XOR|B3|RB
.print DEVI B1|_XOR|T1|1
.print DEVI L1|_XOR|T1|P
.print DEVI R1|_XOR|T1|B
.print DEVI L1|_XOR|T1|RB
.print DEVI B1|_XOR|T2|1
.print DEVI R1|_XOR|T2|B
.print DEVI L1|_XOR|T2|RB
.print DEVI B1|_XOR|AB|1
.print DEVI L1|_XOR|AB|P
.print DEVI R1|_XOR|AB|B
.print DEVI L1|_XOR|AB|RB
.print DEVI B1|_XOR|ABTQ|1
.print DEVI L1|_XOR|ABTQ|P
.print DEVI R1|_XOR|ABTQ|B
.print DEVI L1|_XOR|ABTQ|RB
.print DEVI B1|_XOR|Q1|1
.print DEVI L1|_XOR|Q1|P
.print DEVI R1|_XOR|Q1|B
.print DEVI L1|_XOR|Q1|RB
.print DEVI B1|JTLOUT1|1|1
.print DEVI L1|JTLOUT1|1|P
.print DEVI R1|JTLOUT1|1|B
.print DEVI L1|JTLOUT1|1|RB
.print DEVI L1|JTLOUT1|B|B
.print DEVI I1|JTLOUT1|B|B
.print DEVI B1|JTLOUT1|2|1
.print DEVI L1|JTLOUT1|2|P
.print DEVI R1|JTLOUT1|2|B
.print DEVI L1|JTLOUT1|2|RB
.print DEVI B1|JTLOUT2|1|1
.print DEVI L1|JTLOUT2|1|P
.print DEVI R1|JTLOUT2|1|B
.print DEVI L1|JTLOUT2|1|RB
.print DEVI L1|JTLOUT2|B|B
.print DEVI I1|JTLOUT2|B|B
.print DEVI B1|JTLOUT2|2|1
.print DEVI L1|JTLOUT2|2|P
.print DEVI R1|JTLOUT2|2|B
.print DEVI L1|JTLOUT2|2|RB
.print V 1|_AND_CD|I_5|MID
.print V 1|_AND_CD|B13|MID_SHUNT
.print V 1|D3|1
.print V 1|_NOT|112
.print V 1|_NOT|101
.print V 1|_AND_AB|I_18|MID
.print V 1|_AND_CD|I_1|MID
.print V 1|_XOR|B1|MID_SHUNT
.print V 1|_AND_AB|B4
.print V 1|D2|6
.print V 1|_NOT|8
.print V 1|_AND_CD|B6|MID_SHUNT
.print V 1|_AND_CD|I_31|MID
.print V 1|JTLOUT2|1|MID_SHUNT
.print V 1|_AND_AB|B4|MID_SHUNT
.print V 1|_AND_AB|A5
.print V 1|_NOT|10
.print V 1|_AND_AB|B1
.print V 1|_AND_CD|A5
.print V 1|_AND_CD|T2
.print V 1|D2|2
.print V 1|D2|10
.print V 1|_XOR|B3|MID_SHUNT
.print V 1|JTLOUT2|2|MID_SERIES
.print V 1|ABX
.print V T2
.print V 1|_AND_CD|B4
.print V 1|_NOT|113
.print V 1|D1|11
.print V 1|D3|4
.print V 1|_XOR|B2|MID_SHUNT
.print V 1|_XOR|T2
.print V 1|_NOT|1
.print V 1|_AND_CD|A4
.print V 1|D1|4
.print V 1|_AND_AB|B8|MID_SHUNT
.print V 1|_XOR|A3|MID_SHUNT
.print V 1|D4|7
.print V 1|_NOT|2
.print V 1|_AB_SPL|1
.print V 1|_NOT|14
.print V 1|CD_1
.print V 1|_AND_AB|TB
.print V 1|D1|5
.print V 1|_AND_CD|B3|MID_SERIES
.print V 1|_XOR|I_Q1|MID
.print V 1|_NOT|12
.print V 1|_AND_CD|B3|MID_SHUNT
.print V 1|_AND_AB|B2|MID_SHUNT
.print V 1|_XOR|A3
.print V 1|D4|5
.print V 1|D3|6
.print V 1|_AB_SPL|111
.print V 1|AB_0
.print V 1|_AB_SPL|10
.print V 1|_AB_SPL|8
.print V 1|_AND_AB|A1
.print V 1|_NOT|9
.print V 1|_XOR|T2|MID_SHUNT
.print V 1|_AB_SPL|12
.print V 1|_XOR|I_T1|MID
.print V 1|_XOR|AB|MID_SHUNT
.print V 1|_NOT|121
.print V 1|_AB_SPL|6
.print V 1|_NOT|5
.print V 1|_XOR|B2|MID_SERIES
.print V 1|_XOR|B1
.print V 1|_NOT|11
.print V 1|D1|101
.print V 1|JTLOUT1|6
.print V 1|_AB_SPL|7
.print V 1|_XOR|Q1|MID_SERIES
.print V 1|JTLOUT1|1|MID_SHUNT
.print V 1|JTLOUT2|1|MID_SERIES
.print V 1|_NOT|18
.print V 1|_AND_AB|A4
.print V 1|_XOR|T1
.print V 1|_NOT|104
.print V 1|JTLOUT1|B|MID
.print V 1|_AB_SPL|101
.print V 1|_AND_AB|B3|MID_SERIES
.print V 1|_AND_AB|B15|MID_SERIES
.print V 1|_AND_CD|I_28|MID
.print V 1|D2|11
.print V 1|_NOT|19
.print V 1|D1|9
.print V 1|JTLOUT1|2|MID_SERIES
.print V 1|CD
.print V 1|_NOT|23
.print V 1|_AND_AB|B6|MID_SHUNT
.print V 1|_XOR|A1|MID_SERIES
.print V 1|_NOT|107
.print V 1|_AND_AB|Q1
.print V 1|D4|8
.print V 1|_XOR|AB
.print V 1|D4|2
.print V 1|JTLOUT1|4
.print V 1|_XOR|I_B3|MID
.print V 1|JTLOUT1|2|MID_SHUNT
.print V 1|_XOR|B2
.print V 1|_AND_AB|I_25|MID
.print V 1|_AND_AB|B10|MID_SHUNT
.print V 1|_XOR|ABTQ
.print V 1|D2|4
.print V 1|_AND_CD|B1|MID_SHUNT
.print V 1|D2|104
.print V 1|_AB_SPL|3
.print V 1|_XOR|B3
.print V 1|_XOR|A2|MID_SERIES
.print V 1|_AB_SPL|11
.print V 1|D3|5
.print V 1|_XOR|B1|MID_SERIES
.print V 1|_XOR|A2|MID_SHUNT
.print V 1|_XOR|AB|MID_SERIES
.print V 1|D1|12
.print V 1|_AND_AB|B5|MID_SHUNT
.print V 1|D1|107
.print V D1
.print V 1|_AND_AB|B11|MID_SHUNT
.print V 1|_AND_CD|A2
.print V 1|_AND_AB|B3|MID_SHUNT
.print V B1
.print V 1|D2|107
.print V 1|_AND_AB|B5|MID_SERIES
.print V 1|_AND_CD|I_14|MID
.print V 1|_AND_CD|I_18|MID
.print V 1|_XOR|I_B1|MID
.print V 1|_XOR|B3|MID_SERIES
.print V 1|_AND_CD|TB
.print V 1|D1|3
.print V 1|AB
.print V 1|_AND_CD|I_25|MID
.print V 1|_AND_CD|B11|MID_SHUNT
.print V A1
.print V 1|_XOR|Q1
.print V 1|_AND_CD|B5|MID_SHUNT
.print V 1|_XOR|T1|MID_SERIES
.print V 1|_XOR|A3|MID_SERIES
.print V 1|_AND_CD|B7|MID_SERIES
.print V 1|NOT_AB
.print V 1|D4|3
.print V 1|_AND_AB|TA
.print V 1|AB_1
.print V 1|D3|7
.print V 1|_AND_AB|B12|MID_SHUNT
.print V 1|D4|4
.print V 1|_AND_CD|B11|MID_SERIES
.print V 1|JTLOUT2|B|MID
.print V 1|_AND_AB|B2
.print V 1|_AND_AB|B9|MID_SHUNT
.print V 1|D3|8
.print V 1|_AND_CD|B1
.print V 1|D1|6
.print V 1|_AND_CD|B15|MID_SHUNT
.print V 1|_XOR|T1|MID_SHUNT
.print V AB_XOR_CD_1
.print V 1|_AND_AB|B1|MID_SHUNT
.print V 1|_NOT|15
.print V 1|_NOT|7
.print V 1|_AND_AB|B13|MID_SERIES
.print V 1|_AND_AB|B11|MID_SERIES
.print V 1|_AND_AB|I_31|MID
.print V 1|_AND_CD|B8|MID_SHUNT
.print V 1|_AND_CD|B12|MID_SHUNT
.print V 1|_AND_CD|B10|MID_SHUNT
.print V 1|D1|8
.print V 1|_AB_SPL|4
.print V 1|_AB_SPL|2
.print V 1|_AND_AB|I_5|MID
.print V 1|JTLOUT1|1
.print V 1|JTLOUT2|6
.print V 1|_AND_AB|I_28|MID
.print V 1|_AND_AB|T3
.print V 1|_AND_AB|B1|MID_SERIES
.print V 1|_AND_AB|A3
.print V 1|_AND_CD|B9|MID_SHUNT
.print V 1|_AND_CD|B4|MID_SHUNT
.print V 1|D2|12
.print V 1|_NOT|4
.print V 1|_AND_CD|B1|MID_SERIES
.print V 1|D1|1
.print V 1|CD_0
.print V 1|_AND_CD|T3
.print V 1|D4|6
.print V 1|_AND_CD|B9|MID_SERIES
.print V 1|_AND_CD|Q1
.print V 1|_AND_CD|B2
.print V 1|D2|9
.print V 1|_AND_AB|B13|MID_SHUNT
.print V 1|_NOT|117
.print V 1|_NOT|13
.print V 1|D2|7
.print V 1|_XOR|ABTQ|MID_SERIES
.print V 1|_XOR|I_A1|MID
.print V 1|D2|8
.print V 1|_NOT|120
.print V 1|_AND_CD|B5
.print V 1|D1|104
.print V 1|_AND_AB|T1
.print V 1|_AB_SPL|5
.print V 1|_XOR|I_A3|MID
.print V 1|D1|7
.print V 1|_AND_AB|A2
.print V 1|_AND_AB|B15|MID_SHUNT
.print V 1|D1|110
.print V 1|_AND_CD|B7|MID_SHUNT
.print V 1|D2|101
.print V 1|_XOR|A1
.print V 1|_AND_AB|B14|MID_SHUNT
.print V 1|_NOT|118
.print V 1|_AND_AB|Q2
.print V 1|_AND_AB|B3
.print V C1
.print V 1|_AND_CD|Q2
.print V 1|_AB_SPL|104
.print V 1|_AND_AB|I_14|MID
.print V 1|_XOR|A1|MID_SHUNT
.print V 1|D1|2
.print V 1|_AB_SPL|9
.print V 1|_AND_CD|B2|MID_SHUNT
.print V 1|_NOT|20
.print V 1|_XOR|ABTQ|MID_SHUNT
.print V 1|_AND_AB|B9|MID_SERIES
.print V 1|_AND_CD|A1
.print V 1|_AB_SPL|13
.print V 1|_NOT|3
.print V 1|D4|1
.print V 1|_AND_AB|B5
.print V 1|JTLOUT2|2|MID_SHUNT
.print V 1|_AND_AB|T2
.print V 1|_NOT|6
.print V 1|_AND_CD|B5|MID_SERIES
.print V 1|D2|1
.print V 1|D3|3
.print V 1|ABN
.print V 1|ABXCD
.print V 1|_AND_AB|B7|MID_SERIES
.print V 1|_AND_AB|B14|MID_SERIES
.print V 1|_AND_AB|B7|MID_SHUNT
.print V 1|_NOT|21
.print V 1|_AND_CD|TA
.print V 1|_NOT|16
.print V 1|_AND_CD|T1
.print V 1|D3|2
.print V 1|JTLOUT2|1
.print V T1
.print V 1|D2|5
.print V 1|_AND_AB|I_1|MID
.print V 1|_AND_CD|B13|MID_SERIES
.print V NOT_AB_1
.print V 1|D2|110
.print V 1|_NOT|17
.print V 1|JTLOUT1|1|MID_SERIES
.print V 1|_AND_CD|B14|MID_SERIES
.print V 1|_AND_CD|B3
.print V 1|D2|3
.print V 1|JTLOUT2|4
.print V 1|_NOT|110
.print V 1|_AND_CD|B14|MID_SHUNT
.print V 1|_AND_CD|B15|MID_SERIES
.print V 1|_XOR|Q1|MID_SHUNT
.print V 1|_AND_CD|A3
.print V 1|_NOT|22
.print V 1|_AB_SPL|108
.print V 1|_XOR|A2
.print V 1|D1|10
.print DEVP B1|D1|1
.print DEVP B1|D1|2
.print DEVP B1|D1|3
.print DEVP B1|D1|4
.print DEVP B1|D2|1
.print DEVP B1|D2|2
.print DEVP B1|D2|3
.print DEVP B1|D2|4
.print DEVP B1|D3|1
.print DEVP B1|D3|2
.print DEVP B1|D4|1
.print DEVP B1|D4|2
.print DEVP B1|_AB_SPL|1
.print DEVP B1|_AB_SPL|2
.print DEVP B1|_AB_SPL|3
.print DEVP B1|_AB_SPL|4
.print DEVP B1|_NOT|1
.print DEVP B1|_NOT|2
.print DEVP B1|_NOT|3
.print DEVP B1|_NOT|4
.print DEVP B1|_NOT|5
.print DEVP B1|_NOT|6
.print DEVP B1|_NOT|7
.print DEVP B1|_NOT|8
.print DEVP B1|_NOT|9
.print DEVP B1|_AND_AB|B1|1
.print DEVP B1|_AND_AB|B2|1
.print DEVP B1|_AND_AB|B3|1
.print DEVP B1|_AND_AB|B4|1
.print DEVP B1|_AND_AB|B5|1
.print DEVP B1|_AND_AB|B6|1
.print DEVP B1|_AND_AB|B7|1
.print DEVP B1|_AND_AB|B8|1
.print DEVP B1|_AND_AB|B9|1
.print DEVP B1|_AND_AB|B10|1
.print DEVP B1|_AND_AB|B11|1
.print DEVP B1|_AND_AB|B12|1
.print DEVP B1|_AND_AB|B13|1
.print DEVP B1|_AND_AB|B14|1
.print DEVP B1|_AND_AB|B15|1
.print DEVP B1|_AND_CD|B1|1
.print DEVP B1|_AND_CD|B2|1
.print DEVP B1|_AND_CD|B3|1
.print DEVP B1|_AND_CD|B4|1
.print DEVP B1|_AND_CD|B5|1
.print DEVP B1|_AND_CD|B6|1
.print DEVP B1|_AND_CD|B7|1
.print DEVP B1|_AND_CD|B8|1
.print DEVP B1|_AND_CD|B9|1
.print DEVP B1|_AND_CD|B10|1
.print DEVP B1|_AND_CD|B11|1
.print DEVP B1|_AND_CD|B12|1
.print DEVP B1|_AND_CD|B13|1
.print DEVP B1|_AND_CD|B14|1
.print DEVP B1|_AND_CD|B15|1
.print DEVP B1|_XOR|A1|1
.print DEVP B1|_XOR|A2|1
.print DEVP B1|_XOR|A3|1
.print DEVP B1|_XOR|B1|1
.print DEVP B1|_XOR|B2|1
.print DEVP B1|_XOR|B3|1
.print DEVP B1|_XOR|T1|1
.print DEVP B1|_XOR|T2|1
.print DEVP B1|_XOR|AB|1
.print DEVP B1|_XOR|ABTQ|1
.print DEVP B1|_XOR|Q1|1
.print DEVP B1|JTLOUT1|1|1
.print DEVP B1|JTLOUT1|2|1
.print DEVP B1|JTLOUT2|1|1
.print DEVP B1|JTLOUT2|2|1
