*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM TCLOCK=2e-10
.PARAM OS=5.0000000000000005e-12
.PARAM STEP=0.08
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 1E-12 52000E-12
R_S0 S0 0  1
R_S1 S1 0  1
R_S2 S2 0  1
R_S3 S3 0  1
R_S4 S4 0  1
IA0|A 0 A0  PWL(0 0 3.4e-11 0 3.7e-11 0.0007 4e-11 0 4.34e-10 0 4.37e-10 0.0007 4.4e-10 0 8.34e-10 0 8.37e-10 0.0007 8.4e-10 0 1.234e-09 0 1.237e-09 0.0007 1.24e-09 0 1.634e-09 0 1.637e-09 0.0007 1.64e-09 0 2.034e-09 0 2.037e-09 0.0007 2.04e-09 0 2.434e-09 0 2.437e-09 0.0007 2.44e-09 0 2.834e-09 0 2.837e-09 0.0007 2.84e-09 0 3.234e-09 0 3.237e-09 0.0007 3.24e-09 0 3.634e-09 0 3.637e-09 0.0007 3.64e-09 0 4.034e-09 0 4.037e-09 0.0007 4.04e-09 0 4.434e-09 0 4.437e-09 0.0007 4.44e-09 0 4.834e-09 0 4.837e-09 0.0007 4.84e-09 0 5.234e-09 0 5.237e-09 0.0007 5.24e-09 0 5.634e-09 0 5.637e-09 0.0007 5.64e-09 0 6.034e-09 0 6.037e-09 0.0007 6.04e-09 0 6.434e-09 0 6.437e-09 0.0007 6.44e-09 0 6.834e-09 0 6.837e-09 0.0007 6.84e-09 0 7.234e-09 0 7.237e-09 0.0007 7.24e-09 0 7.634e-09 0 7.637e-09 0.0007 7.64e-09 0 8.034e-09 0 8.037e-09 0.0007 8.04e-09 0 8.434e-09 0 8.437e-09 0.0007 8.44e-09 0 8.834e-09 0 8.837e-09 0.0007 8.84e-09 0 9.234e-09 0 9.237e-09 0.0007 9.24e-09 0 9.634e-09 0 9.637e-09 0.0007 9.64e-09 0 1.0034e-08 0 1.0037e-08 0.0007 1.004e-08 0 1.0434e-08 0 1.0437e-08 0.0007 1.044e-08 0 1.0834e-08 0 1.0837e-08 0.0007 1.084e-08 0 1.1234e-08 0 1.1237e-08 0.0007 1.124e-08 0 1.1634e-08 0 1.1637e-08 0.0007 1.164e-08 0 1.2034e-08 0 1.2037e-08 0.0007 1.204e-08 0 1.2434e-08 0 1.2437e-08 0.0007 1.244e-08 0 1.2834e-08 0 1.2837e-08 0.0007 1.284e-08 0 1.3234e-08 0 1.3237e-08 0.0007 1.324e-08 0 1.3634e-08 0 1.3637e-08 0.0007 1.364e-08 0 1.4034e-08 0 1.4037e-08 0.0007 1.404e-08 0 1.4434e-08 0 1.4437e-08 0.0007 1.444e-08 0 1.4834e-08 0 1.4837e-08 0.0007 1.484e-08 0 1.5234e-08 0 1.5237e-08 0.0007 1.524e-08 0 1.5634e-08 0 1.5637e-08 0.0007 1.564e-08 0 1.6034e-08 0 1.6037e-08 0.0007 1.604e-08 0 1.6434e-08 0 1.6437e-08 0.0007 1.644e-08 0 1.6834e-08 0 1.6837e-08 0.0007 1.684e-08 0 1.7234e-08 0 1.7237e-08 0.0007 1.724e-08 0 1.7634e-08 0 1.7637e-08 0.0007 1.764e-08 0 1.8034e-08 0 1.8037e-08 0.0007 1.804e-08 0 1.8434e-08 0 1.8437e-08 0.0007 1.844e-08 0 1.8834e-08 0 1.8837e-08 0.0007 1.884e-08 0 1.9234e-08 0 1.9237e-08 0.0007 1.924e-08 0 1.9634e-08 0 1.9637e-08 0.0007 1.964e-08 0 2.0034e-08 0 2.0037e-08 0.0007 2.004e-08 0 2.0434e-08 0 2.0437e-08 0.0007 2.044e-08 0 2.0834e-08 0 2.0837e-08 0.0007 2.084e-08 0 2.1234e-08 0 2.1237e-08 0.0007 2.124e-08 0 2.1634e-08 0 2.1637e-08 0.0007 2.164e-08 0 2.2034e-08 0 2.2037e-08 0.0007 2.204e-08 0 2.2434e-08 0 2.2437e-08 0.0007 2.244e-08 0 2.2834e-08 0 2.2837e-08 0.0007 2.284e-08 0 2.3234e-08 0 2.3237e-08 0.0007 2.324e-08 0 2.3634e-08 0 2.3637e-08 0.0007 2.364e-08 0 2.4034e-08 0 2.4037e-08 0.0007 2.404e-08 0 2.4434e-08 0 2.4437e-08 0.0007 2.444e-08 0 2.4834e-08 0 2.4837e-08 0.0007 2.484e-08 0 2.5234e-08 0 2.5237e-08 0.0007 2.524e-08 0 2.5634e-08 0 2.5637e-08 0.0007 2.564e-08 0 2.6034e-08 0 2.6037e-08 0.0007 2.604e-08 0 2.6434e-08 0 2.6437e-08 0.0007 2.644e-08 0 2.6834e-08 0 2.6837e-08 0.0007 2.684e-08 0 2.7234e-08 0 2.7237e-08 0.0007 2.724e-08 0 2.7634e-08 0 2.7637e-08 0.0007 2.764e-08 0 2.8034e-08 0 2.8037e-08 0.0007 2.804e-08 0 2.8434e-08 0 2.8437e-08 0.0007 2.844e-08 0 2.8834e-08 0 2.8837e-08 0.0007 2.884e-08 0 2.9234e-08 0 2.9237e-08 0.0007 2.924e-08 0 2.9634e-08 0 2.9637e-08 0.0007 2.964e-08 0 3.0034e-08 0 3.0037e-08 0.0007 3.004e-08 0 3.0434e-08 0 3.0437e-08 0.0007 3.044e-08 0 3.0834e-08 0 3.0837e-08 0.0007 3.084e-08 0 3.1234e-08 0 3.1237e-08 0.0007 3.124e-08 0 3.1634e-08 0 3.1637e-08 0.0007 3.164e-08 0 3.2034e-08 0 3.2037e-08 0.0007 3.204e-08 0 3.2434e-08 0 3.2437e-08 0.0007 3.244e-08 0 3.2834e-08 0 3.2837e-08 0.0007 3.284e-08 0 3.3234e-08 0 3.3237e-08 0.0007 3.324e-08 0 3.3634e-08 0 3.3637e-08 0.0007 3.364e-08 0 3.4034e-08 0 3.4037e-08 0.0007 3.404e-08 0 3.4434e-08 0 3.4437e-08 0.0007 3.444e-08 0 3.4834e-08 0 3.4837e-08 0.0007 3.484e-08 0 3.5234e-08 0 3.5237e-08 0.0007 3.524e-08 0 3.5634e-08 0 3.5637e-08 0.0007 3.564e-08 0 3.6034e-08 0 3.6037e-08 0.0007 3.604e-08 0 3.6434e-08 0 3.6437e-08 0.0007 3.644e-08 0 3.6834e-08 0 3.6837e-08 0.0007 3.684e-08 0 3.7234e-08 0 3.7237e-08 0.0007 3.724e-08 0 3.7634e-08 0 3.7637e-08 0.0007 3.764e-08 0 3.8034e-08 0 3.8037e-08 0.0007 3.804e-08 0 3.8434e-08 0 3.8437e-08 0.0007 3.844e-08 0 3.8834e-08 0 3.8837e-08 0.0007 3.884e-08 0 3.9234e-08 0 3.9237e-08 0.0007 3.924e-08 0 3.9634e-08 0 3.9637e-08 0.0007 3.964e-08 0 4.0034e-08 0 4.0037e-08 0.0007 4.004e-08 0 4.0434e-08 0 4.0437e-08 0.0007 4.044e-08 0 4.0834e-08 0 4.0837e-08 0.0007 4.084e-08 0 4.1234e-08 0 4.1237e-08 0.0007 4.124e-08 0 4.1634e-08 0 4.1637e-08 0.0007 4.164e-08 0 4.2034e-08 0 4.2037e-08 0.0007 4.204e-08 0 4.2434e-08 0 4.2437e-08 0.0007 4.244e-08 0 4.2834e-08 0 4.2837e-08 0.0007 4.284e-08 0 4.3234e-08 0 4.3237e-08 0.0007 4.324e-08 0 4.3634e-08 0 4.3637e-08 0.0007 4.364e-08 0 4.4034e-08 0 4.4037e-08 0.0007 4.404e-08 0 4.4434e-08 0 4.4437e-08 0.0007 4.444e-08 0 4.4834e-08 0 4.4837e-08 0.0007 4.484e-08 0 4.5234e-08 0 4.5237e-08 0.0007 4.524e-08 0 4.5634e-08 0 4.5637e-08 0.0007 4.564e-08 0 4.6034e-08 0 4.6037e-08 0.0007 4.604e-08 0 4.6434e-08 0 4.6437e-08 0.0007 4.644e-08 0 4.6834e-08 0 4.6837e-08 0.0007 4.684e-08 0 4.7234e-08 0 4.7237e-08 0.0007 4.724e-08 0 4.7634e-08 0 4.7637e-08 0.0007 4.764e-08 0 4.8034e-08 0 4.8037e-08 0.0007 4.804e-08 0 4.8434e-08 0 4.8437e-08 0.0007 4.844e-08 0 4.8834e-08 0 4.8837e-08 0.0007 4.884e-08 0 4.9234e-08 0 4.9237e-08 0.0007 4.924e-08 0 4.9634e-08 0 4.9637e-08 0.0007 4.964e-08 0 5.0034e-08 0 5.0037e-08 0.0007 5.004e-08 0 5.0434e-08 0 5.0437e-08 0.0007 5.044e-08 0 5.0834e-08 0 5.0837e-08 0.0007 5.084e-08 0)
IB0|B 0 B0  PWL(0 0 5e-11 0 5.3e-11 0.0007 5.6e-11 0 2.5e-10 0 2.53e-10 0.0007 2.56e-10 0 8.5e-10 0 8.53e-10 0.0007 8.56e-10 0 1.05e-09 0 1.053e-09 0.0007 1.056e-09 0 1.65e-09 0 1.653e-09 0.0007 1.656e-09 0 1.85e-09 0 1.853e-09 0.0007 1.856e-09 0 2.45e-09 0 2.453e-09 0.0007 2.456e-09 0 2.65e-09 0 2.653e-09 0.0007 2.656e-09 0 3.25e-09 0 3.253e-09 0.0007 3.256e-09 0 3.45e-09 0 3.453e-09 0.0007 3.456e-09 0 4.05e-09 0 4.053e-09 0.0007 4.056e-09 0 4.25e-09 0 4.253e-09 0.0007 4.256e-09 0 4.85e-09 0 4.853e-09 0.0007 4.856e-09 0 5.05e-09 0 5.053e-09 0.0007 5.056e-09 0 5.65e-09 0 5.653e-09 0.0007 5.656e-09 0 5.85e-09 0 5.853e-09 0.0007 5.856e-09 0 6.45e-09 0 6.453e-09 0.0007 6.456e-09 0 6.65e-09 0 6.653e-09 0.0007 6.656e-09 0 7.25e-09 0 7.253e-09 0.0007 7.256e-09 0 7.45e-09 0 7.453e-09 0.0007 7.456e-09 0 8.05e-09 0 8.053e-09 0.0007 8.056e-09 0 8.25e-09 0 8.253e-09 0.0007 8.256e-09 0 8.85e-09 0 8.853e-09 0.0007 8.856e-09 0 9.05e-09 0 9.053e-09 0.0007 9.056e-09 0 9.65e-09 0 9.653e-09 0.0007 9.656e-09 0 9.85e-09 0 9.853e-09 0.0007 9.856e-09 0 1.045e-08 0 1.0453e-08 0.0007 1.0456e-08 0 1.065e-08 0 1.0653e-08 0.0007 1.0656e-08 0 1.125e-08 0 1.1253e-08 0.0007 1.1256e-08 0 1.145e-08 0 1.1453e-08 0.0007 1.1456e-08 0 1.205e-08 0 1.2053e-08 0.0007 1.2056e-08 0 1.225e-08 0 1.2253e-08 0.0007 1.2256e-08 0 1.285e-08 0 1.2853e-08 0.0007 1.2856e-08 0 1.305e-08 0 1.3053e-08 0.0007 1.3056e-08 0 1.365e-08 0 1.3653e-08 0.0007 1.3656e-08 0 1.385e-08 0 1.3853e-08 0.0007 1.3856e-08 0 1.445e-08 0 1.4453e-08 0.0007 1.4456e-08 0 1.465e-08 0 1.4653e-08 0.0007 1.4656e-08 0 1.525e-08 0 1.5253e-08 0.0007 1.5256e-08 0 1.545e-08 0 1.5453e-08 0.0007 1.5456e-08 0 1.605e-08 0 1.6053e-08 0.0007 1.6056e-08 0 1.625e-08 0 1.6253e-08 0.0007 1.6256e-08 0 1.685e-08 0 1.6853e-08 0.0007 1.6856e-08 0 1.705e-08 0 1.7053e-08 0.0007 1.7056e-08 0 1.765e-08 0 1.7653e-08 0.0007 1.7656e-08 0 1.785e-08 0 1.7853e-08 0.0007 1.7856e-08 0 1.845e-08 0 1.8453e-08 0.0007 1.8456e-08 0 1.865e-08 0 1.8653e-08 0.0007 1.8656e-08 0 1.925e-08 0 1.9253e-08 0.0007 1.9256e-08 0 1.945e-08 0 1.9453e-08 0.0007 1.9456e-08 0 2.005e-08 0 2.0053e-08 0.0007 2.0056e-08 0 2.025e-08 0 2.0253e-08 0.0007 2.0256e-08 0 2.085e-08 0 2.0853e-08 0.0007 2.0856e-08 0 2.105e-08 0 2.1053e-08 0.0007 2.1056e-08 0 2.165e-08 0 2.1653e-08 0.0007 2.1656e-08 0 2.185e-08 0 2.1853e-08 0.0007 2.1856e-08 0 2.245e-08 0 2.2453e-08 0.0007 2.2456e-08 0 2.265e-08 0 2.2653e-08 0.0007 2.2656e-08 0 2.325e-08 0 2.3253e-08 0.0007 2.3256e-08 0 2.345e-08 0 2.3453e-08 0.0007 2.3456e-08 0 2.405e-08 0 2.4053e-08 0.0007 2.4056e-08 0 2.425e-08 0 2.4253e-08 0.0007 2.4256e-08 0 2.485e-08 0 2.4853e-08 0.0007 2.4856e-08 0 2.505e-08 0 2.5053e-08 0.0007 2.5056e-08 0 2.565e-08 0 2.5653e-08 0.0007 2.5656e-08 0 2.585e-08 0 2.5853e-08 0.0007 2.5856e-08 0 2.645e-08 0 2.6453e-08 0.0007 2.6456e-08 0 2.665e-08 0 2.6653e-08 0.0007 2.6656e-08 0 2.725e-08 0 2.7253e-08 0.0007 2.7256e-08 0 2.745e-08 0 2.7453e-08 0.0007 2.7456e-08 0 2.805e-08 0 2.8053e-08 0.0007 2.8056e-08 0 2.825e-08 0 2.8253e-08 0.0007 2.8256e-08 0 2.885e-08 0 2.8853e-08 0.0007 2.8856e-08 0 2.905e-08 0 2.9053e-08 0.0007 2.9056e-08 0 2.965e-08 0 2.9653e-08 0.0007 2.9656e-08 0 2.985e-08 0 2.9853e-08 0.0007 2.9856e-08 0 3.045e-08 0 3.0453e-08 0.0007 3.0456e-08 0 3.065e-08 0 3.0653e-08 0.0007 3.0656e-08 0 3.125e-08 0 3.1253e-08 0.0007 3.1256e-08 0 3.145e-08 0 3.1453e-08 0.0007 3.1456e-08 0 3.205e-08 0 3.2053e-08 0.0007 3.2056e-08 0 3.225e-08 0 3.2253e-08 0.0007 3.2256e-08 0 3.285e-08 0 3.2853e-08 0.0007 3.2856e-08 0 3.305e-08 0 3.3053e-08 0.0007 3.3056e-08 0 3.365e-08 0 3.3653e-08 0.0007 3.3656e-08 0 3.385e-08 0 3.3853e-08 0.0007 3.3856e-08 0 3.445e-08 0 3.4453e-08 0.0007 3.4456e-08 0 3.465e-08 0 3.4653e-08 0.0007 3.4656e-08 0 3.525e-08 0 3.5253e-08 0.0007 3.5256e-08 0 3.545e-08 0 3.5453e-08 0.0007 3.5456e-08 0 3.605e-08 0 3.6053e-08 0.0007 3.6056e-08 0 3.625e-08 0 3.6253e-08 0.0007 3.6256e-08 0 3.685e-08 0 3.6853e-08 0.0007 3.6856e-08 0 3.705e-08 0 3.7053e-08 0.0007 3.7056e-08 0 3.765e-08 0 3.7653e-08 0.0007 3.7656e-08 0 3.785e-08 0 3.7853e-08 0.0007 3.7856e-08 0 3.845e-08 0 3.8453e-08 0.0007 3.8456e-08 0 3.865e-08 0 3.8653e-08 0.0007 3.8656e-08 0 3.925e-08 0 3.9253e-08 0.0007 3.9256e-08 0 3.945e-08 0 3.9453e-08 0.0007 3.9456e-08 0 4.005e-08 0 4.0053e-08 0.0007 4.0056e-08 0 4.025e-08 0 4.0253e-08 0.0007 4.0256e-08 0 4.085e-08 0 4.0853e-08 0.0007 4.0856e-08 0 4.105e-08 0 4.1053e-08 0.0007 4.1056e-08 0 4.165e-08 0 4.1653e-08 0.0007 4.1656e-08 0 4.185e-08 0 4.1853e-08 0.0007 4.1856e-08 0 4.245e-08 0 4.2453e-08 0.0007 4.2456e-08 0 4.265e-08 0 4.2653e-08 0.0007 4.2656e-08 0 4.325e-08 0 4.3253e-08 0.0007 4.3256e-08 0 4.345e-08 0 4.3453e-08 0.0007 4.3456e-08 0 4.405e-08 0 4.4053e-08 0.0007 4.4056e-08 0 4.425e-08 0 4.4253e-08 0.0007 4.4256e-08 0 4.485e-08 0 4.4853e-08 0.0007 4.4856e-08 0 4.505e-08 0 4.5053e-08 0.0007 4.5056e-08 0 4.565e-08 0 4.5653e-08 0.0007 4.5656e-08 0 4.585e-08 0 4.5853e-08 0.0007 4.5856e-08 0 4.645e-08 0 4.6453e-08 0.0007 4.6456e-08 0 4.665e-08 0 4.6653e-08 0.0007 4.6656e-08 0 4.725e-08 0 4.7253e-08 0.0007 4.7256e-08 0 4.745e-08 0 4.7453e-08 0.0007 4.7456e-08 0 4.805e-08 0 4.8053e-08 0.0007 4.8056e-08 0 4.825e-08 0 4.8253e-08 0.0007 4.8256e-08 0 4.885e-08 0 4.8853e-08 0.0007 4.8856e-08 0 4.905e-08 0 4.9053e-08 0.0007 4.9056e-08 0 4.965e-08 0 4.9653e-08 0.0007 4.9656e-08 0 4.985e-08 0 4.9853e-08 0.0007 4.9856e-08 0 5.045e-08 0 5.0453e-08 0.0007 5.0456e-08 0 5.065e-08 0 5.0653e-08 0.0007 5.0656e-08 0)
IA1|C 0 A1  PWL(0 0 6.6e-11 0 6.9e-11 0.0007 7.2e-11 0 2.66e-10 0 2.69e-10 0.0007 2.72e-10 0 4.66e-10 0 4.69e-10 0.0007 4.72e-10 0 6.66e-10 0 6.69e-10 0.0007 6.72e-10 0 1.666e-09 0 1.669e-09 0.0007 1.672e-09 0 1.866e-09 0 1.869e-09 0.0007 1.872e-09 0 2.066e-09 0 2.069e-09 0.0007 2.072e-09 0 2.266e-09 0 2.269e-09 0.0007 2.272e-09 0 3.266e-09 0 3.269e-09 0.0007 3.272e-09 0 3.466e-09 0 3.469e-09 0.0007 3.472e-09 0 3.666e-09 0 3.669e-09 0.0007 3.672e-09 0 3.866e-09 0 3.869e-09 0.0007 3.872e-09 0 4.866e-09 0 4.869e-09 0.0007 4.872e-09 0 5.066e-09 0 5.069e-09 0.0007 5.072e-09 0 5.266e-09 0 5.269e-09 0.0007 5.272e-09 0 5.466e-09 0 5.469e-09 0.0007 5.472e-09 0 6.466e-09 0 6.469e-09 0.0007 6.472e-09 0 6.666e-09 0 6.669e-09 0.0007 6.672e-09 0 6.866e-09 0 6.869e-09 0.0007 6.872e-09 0 7.066e-09 0 7.069e-09 0.0007 7.072e-09 0 8.066e-09 0 8.069e-09 0.0007 8.072e-09 0 8.266e-09 0 8.269e-09 0.0007 8.272e-09 0 8.466e-09 0 8.469e-09 0.0007 8.472e-09 0 8.666e-09 0 8.669e-09 0.0007 8.672e-09 0 9.666e-09 0 9.669e-09 0.0007 9.672e-09 0 9.866e-09 0 9.869e-09 0.0007 9.872e-09 0 1.0066e-08 0 1.0069e-08 0.0007 1.0072e-08 0 1.0266e-08 0 1.0269e-08 0.0007 1.0272e-08 0 1.1266e-08 0 1.1269e-08 0.0007 1.1272e-08 0 1.1466e-08 0 1.1469e-08 0.0007 1.1472e-08 0 1.1666e-08 0 1.1669e-08 0.0007 1.1672e-08 0 1.1866e-08 0 1.1869e-08 0.0007 1.1872e-08 0 1.2866e-08 0 1.2869e-08 0.0007 1.2872e-08 0 1.3066e-08 0 1.3069e-08 0.0007 1.3072e-08 0 1.3266e-08 0 1.3269e-08 0.0007 1.3272e-08 0 1.3466e-08 0 1.3469e-08 0.0007 1.3472e-08 0 1.4466e-08 0 1.4469e-08 0.0007 1.4472e-08 0 1.4666e-08 0 1.4669e-08 0.0007 1.4672e-08 0 1.4866e-08 0 1.4869e-08 0.0007 1.4872e-08 0 1.5066e-08 0 1.5069e-08 0.0007 1.5072e-08 0 1.6066e-08 0 1.6069e-08 0.0007 1.6072e-08 0 1.6266e-08 0 1.6269e-08 0.0007 1.6272e-08 0 1.6466e-08 0 1.6469e-08 0.0007 1.6472e-08 0 1.6666e-08 0 1.6669e-08 0.0007 1.6672e-08 0 1.7666e-08 0 1.7669e-08 0.0007 1.7672e-08 0 1.7866e-08 0 1.7869e-08 0.0007 1.7872e-08 0 1.8066e-08 0 1.8069e-08 0.0007 1.8072e-08 0 1.8266e-08 0 1.8269e-08 0.0007 1.8272e-08 0 1.9266e-08 0 1.9269e-08 0.0007 1.9272e-08 0 1.9466e-08 0 1.9469e-08 0.0007 1.9472e-08 0 1.9666e-08 0 1.9669e-08 0.0007 1.9672e-08 0 1.9866e-08 0 1.9869e-08 0.0007 1.9872e-08 0 2.0866e-08 0 2.0869e-08 0.0007 2.0872e-08 0 2.1066e-08 0 2.1069e-08 0.0007 2.1072e-08 0 2.1266e-08 0 2.1269e-08 0.0007 2.1272e-08 0 2.1466e-08 0 2.1469e-08 0.0007 2.1472e-08 0 2.2466e-08 0 2.2469e-08 0.0007 2.2472e-08 0 2.2666e-08 0 2.2669e-08 0.0007 2.2672e-08 0 2.2866e-08 0 2.2869e-08 0.0007 2.2872e-08 0 2.3066e-08 0 2.3069e-08 0.0007 2.3072e-08 0 2.4066e-08 0 2.4069e-08 0.0007 2.4072e-08 0 2.4266e-08 0 2.4269e-08 0.0007 2.4272e-08 0 2.4466e-08 0 2.4469e-08 0.0007 2.4472e-08 0 2.4666e-08 0 2.4669e-08 0.0007 2.4672e-08 0 2.5666e-08 0 2.5669e-08 0.0007 2.5672e-08 0 2.5866e-08 0 2.5869e-08 0.0007 2.5872e-08 0 2.6066e-08 0 2.6069e-08 0.0007 2.6072e-08 0 2.6266e-08 0 2.6269e-08 0.0007 2.6272e-08 0 2.7266e-08 0 2.7269e-08 0.0007 2.7272e-08 0 2.7466e-08 0 2.7469e-08 0.0007 2.7472e-08 0 2.7666e-08 0 2.7669e-08 0.0007 2.7672e-08 0 2.7866e-08 0 2.7869e-08 0.0007 2.7872e-08 0 2.8866e-08 0 2.8869e-08 0.0007 2.8872e-08 0 2.9066e-08 0 2.9069e-08 0.0007 2.9072e-08 0 2.9266e-08 0 2.9269e-08 0.0007 2.9272e-08 0 2.9466e-08 0 2.9469e-08 0.0007 2.9472e-08 0 3.0466e-08 0 3.0469e-08 0.0007 3.0472e-08 0 3.0666e-08 0 3.0669e-08 0.0007 3.0672e-08 0 3.0866e-08 0 3.0869e-08 0.0007 3.0872e-08 0 3.1066e-08 0 3.1069e-08 0.0007 3.1072e-08 0 3.2066e-08 0 3.2069e-08 0.0007 3.2072e-08 0 3.2266e-08 0 3.2269e-08 0.0007 3.2272e-08 0 3.2466e-08 0 3.2469e-08 0.0007 3.2472e-08 0 3.2666e-08 0 3.2669e-08 0.0007 3.2672e-08 0 3.3666e-08 0 3.3669e-08 0.0007 3.3672e-08 0 3.3866e-08 0 3.3869e-08 0.0007 3.3872e-08 0 3.4066e-08 0 3.4069e-08 0.0007 3.4072e-08 0 3.4266e-08 0 3.4269e-08 0.0007 3.4272e-08 0 3.5266e-08 0 3.5269e-08 0.0007 3.5272e-08 0 3.5466e-08 0 3.5469e-08 0.0007 3.5472e-08 0 3.5666e-08 0 3.5669e-08 0.0007 3.5672e-08 0 3.5866e-08 0 3.5869e-08 0.0007 3.5872e-08 0 3.6866e-08 0 3.6869e-08 0.0007 3.6872e-08 0 3.7066e-08 0 3.7069e-08 0.0007 3.7072e-08 0 3.7266e-08 0 3.7269e-08 0.0007 3.7272e-08 0 3.7466e-08 0 3.7469e-08 0.0007 3.7472e-08 0 3.8466e-08 0 3.8469e-08 0.0007 3.8472e-08 0 3.8666e-08 0 3.8669e-08 0.0007 3.8672e-08 0 3.8866e-08 0 3.8869e-08 0.0007 3.8872e-08 0 3.9066e-08 0 3.9069e-08 0.0007 3.9072e-08 0 4.0066e-08 0 4.0069e-08 0.0007 4.0072e-08 0 4.0266e-08 0 4.0269e-08 0.0007 4.0272e-08 0 4.0466e-08 0 4.0469e-08 0.0007 4.0472e-08 0 4.0666e-08 0 4.0669e-08 0.0007 4.0672e-08 0 4.1666e-08 0 4.1669e-08 0.0007 4.1672e-08 0 4.1866e-08 0 4.1869e-08 0.0007 4.1872e-08 0 4.2066e-08 0 4.2069e-08 0.0007 4.2072e-08 0 4.2266e-08 0 4.2269e-08 0.0007 4.2272e-08 0 4.3266e-08 0 4.3269e-08 0.0007 4.3272e-08 0 4.3466e-08 0 4.3469e-08 0.0007 4.3472e-08 0 4.3666e-08 0 4.3669e-08 0.0007 4.3672e-08 0 4.3866e-08 0 4.3869e-08 0.0007 4.3872e-08 0 4.4866e-08 0 4.4869e-08 0.0007 4.4872e-08 0 4.5066e-08 0 4.5069e-08 0.0007 4.5072e-08 0 4.5266e-08 0 4.5269e-08 0.0007 4.5272e-08 0 4.5466e-08 0 4.5469e-08 0.0007 4.5472e-08 0 4.6466e-08 0 4.6469e-08 0.0007 4.6472e-08 0 4.6666e-08 0 4.6669e-08 0.0007 4.6672e-08 0 4.6866e-08 0 4.6869e-08 0.0007 4.6872e-08 0 4.7066e-08 0 4.7069e-08 0.0007 4.7072e-08 0 4.8066e-08 0 4.8069e-08 0.0007 4.8072e-08 0 4.8266e-08 0 4.8269e-08 0.0007 4.8272e-08 0 4.8466e-08 0 4.8469e-08 0.0007 4.8472e-08 0 4.8666e-08 0 4.8669e-08 0.0007 4.8672e-08 0 4.9666e-08 0 4.9669e-08 0.0007 4.9672e-08 0 4.9866e-08 0 4.9869e-08 0.0007 4.9872e-08 0 5.0066e-08 0 5.0069e-08 0.0007 5.0072e-08 0 5.0266e-08 0 5.0269e-08 0.0007 5.0272e-08 0)
IB1|D 0 B1  PWL(0 0 8.2e-11 0 8.5e-11 0.0007 8.8e-11 0 2.82e-10 0 2.85e-10 0.0007 2.88e-10 0 4.82e-10 0 4.85e-10 0.0007 4.88e-10 0 6.82e-10 0 6.85e-10 0.0007 6.88e-10 0 8.82e-10 0 8.85e-10 0.0007 8.88e-10 0 1.082e-09 0 1.085e-09 0.0007 1.088e-09 0 1.282e-09 0 1.285e-09 0.0007 1.288e-09 0 1.482e-09 0 1.485e-09 0.0007 1.488e-09 0 3.282e-09 0 3.285e-09 0.0007 3.288e-09 0 3.482e-09 0 3.485e-09 0.0007 3.488e-09 0 3.682e-09 0 3.685e-09 0.0007 3.688e-09 0 3.882e-09 0 3.885e-09 0.0007 3.888e-09 0 4.082e-09 0 4.085e-09 0.0007 4.088e-09 0 4.282e-09 0 4.285e-09 0.0007 4.288e-09 0 4.482e-09 0 4.485e-09 0.0007 4.488e-09 0 4.682e-09 0 4.685e-09 0.0007 4.688e-09 0 6.482e-09 0 6.485e-09 0.0007 6.488e-09 0 6.682e-09 0 6.685e-09 0.0007 6.688e-09 0 6.882e-09 0 6.885e-09 0.0007 6.888e-09 0 7.082e-09 0 7.085e-09 0.0007 7.088e-09 0 7.282e-09 0 7.285e-09 0.0007 7.288e-09 0 7.482e-09 0 7.485e-09 0.0007 7.488e-09 0 7.682e-09 0 7.685e-09 0.0007 7.688e-09 0 7.882e-09 0 7.885e-09 0.0007 7.888e-09 0 9.682e-09 0 9.685e-09 0.0007 9.688e-09 0 9.882e-09 0 9.885e-09 0.0007 9.888e-09 0 1.0082e-08 0 1.0085e-08 0.0007 1.0088e-08 0 1.0282e-08 0 1.0285e-08 0.0007 1.0288e-08 0 1.0482e-08 0 1.0485e-08 0.0007 1.0488e-08 0 1.0682e-08 0 1.0685e-08 0.0007 1.0688e-08 0 1.0882e-08 0 1.0885e-08 0.0007 1.0888e-08 0 1.1082e-08 0 1.1085e-08 0.0007 1.1088e-08 0 1.2882e-08 0 1.2885e-08 0.0007 1.2888e-08 0 1.3082e-08 0 1.3085e-08 0.0007 1.3088e-08 0 1.3282e-08 0 1.3285e-08 0.0007 1.3288e-08 0 1.3482e-08 0 1.3485e-08 0.0007 1.3488e-08 0 1.3682e-08 0 1.3685e-08 0.0007 1.3688e-08 0 1.3882e-08 0 1.3885e-08 0.0007 1.3888e-08 0 1.4082e-08 0 1.4085e-08 0.0007 1.4088e-08 0 1.4282e-08 0 1.4285e-08 0.0007 1.4288e-08 0 1.6082e-08 0 1.6085e-08 0.0007 1.6088e-08 0 1.6282e-08 0 1.6285e-08 0.0007 1.6288e-08 0 1.6482e-08 0 1.6485e-08 0.0007 1.6488e-08 0 1.6682e-08 0 1.6685e-08 0.0007 1.6688e-08 0 1.6882e-08 0 1.6885e-08 0.0007 1.6888e-08 0 1.7082e-08 0 1.7085e-08 0.0007 1.7088e-08 0 1.7282e-08 0 1.7285e-08 0.0007 1.7288e-08 0 1.7482e-08 0 1.7485e-08 0.0007 1.7488e-08 0 1.9282e-08 0 1.9285e-08 0.0007 1.9288e-08 0 1.9482e-08 0 1.9485e-08 0.0007 1.9488e-08 0 1.9682e-08 0 1.9685e-08 0.0007 1.9688e-08 0 1.9882e-08 0 1.9885e-08 0.0007 1.9888e-08 0 2.0082e-08 0 2.0085e-08 0.0007 2.0088e-08 0 2.0282e-08 0 2.0285e-08 0.0007 2.0288e-08 0 2.0482e-08 0 2.0485e-08 0.0007 2.0488e-08 0 2.0682e-08 0 2.0685e-08 0.0007 2.0688e-08 0 2.2482e-08 0 2.2485e-08 0.0007 2.2488e-08 0 2.2682e-08 0 2.2685e-08 0.0007 2.2688e-08 0 2.2882e-08 0 2.2885e-08 0.0007 2.2888e-08 0 2.3082e-08 0 2.3085e-08 0.0007 2.3088e-08 0 2.3282e-08 0 2.3285e-08 0.0007 2.3288e-08 0 2.3482e-08 0 2.3485e-08 0.0007 2.3488e-08 0 2.3682e-08 0 2.3685e-08 0.0007 2.3688e-08 0 2.3882e-08 0 2.3885e-08 0.0007 2.3888e-08 0 2.5682e-08 0 2.5685e-08 0.0007 2.5688e-08 0 2.5882e-08 0 2.5885e-08 0.0007 2.5888e-08 0 2.6082e-08 0 2.6085e-08 0.0007 2.6088e-08 0 2.6282e-08 0 2.6285e-08 0.0007 2.6288e-08 0 2.6482e-08 0 2.6485e-08 0.0007 2.6488e-08 0 2.6682e-08 0 2.6685e-08 0.0007 2.6688e-08 0 2.6882e-08 0 2.6885e-08 0.0007 2.6888e-08 0 2.7082e-08 0 2.7085e-08 0.0007 2.7088e-08 0 2.8882e-08 0 2.8885e-08 0.0007 2.8888e-08 0 2.9082e-08 0 2.9085e-08 0.0007 2.9088e-08 0 2.9282e-08 0 2.9285e-08 0.0007 2.9288e-08 0 2.9482e-08 0 2.9485e-08 0.0007 2.9488e-08 0 2.9682e-08 0 2.9685e-08 0.0007 2.9688e-08 0 2.9882e-08 0 2.9885e-08 0.0007 2.9888e-08 0 3.0082e-08 0 3.0085e-08 0.0007 3.0088e-08 0 3.0282e-08 0 3.0285e-08 0.0007 3.0288e-08 0 3.2082e-08 0 3.2085e-08 0.0007 3.2088e-08 0 3.2282e-08 0 3.2285e-08 0.0007 3.2288e-08 0 3.2482e-08 0 3.2485e-08 0.0007 3.2488e-08 0 3.2682e-08 0 3.2685e-08 0.0007 3.2688e-08 0 3.2882e-08 0 3.2885e-08 0.0007 3.2888e-08 0 3.3082e-08 0 3.3085e-08 0.0007 3.3088e-08 0 3.3282e-08 0 3.3285e-08 0.0007 3.3288e-08 0 3.3482e-08 0 3.3485e-08 0.0007 3.3488e-08 0 3.5282e-08 0 3.5285e-08 0.0007 3.5288e-08 0 3.5482e-08 0 3.5485e-08 0.0007 3.5488e-08 0 3.5682e-08 0 3.5685e-08 0.0007 3.5688e-08 0 3.5882e-08 0 3.5885e-08 0.0007 3.5888e-08 0 3.6082e-08 0 3.6085e-08 0.0007 3.6088e-08 0 3.6282e-08 0 3.6285e-08 0.0007 3.6288e-08 0 3.6482e-08 0 3.6485e-08 0.0007 3.6488e-08 0 3.6682e-08 0 3.6685e-08 0.0007 3.6688e-08 0 3.8482e-08 0 3.8485e-08 0.0007 3.8488e-08 0 3.8682e-08 0 3.8685e-08 0.0007 3.8688e-08 0 3.8882e-08 0 3.8885e-08 0.0007 3.8888e-08 0 3.9082e-08 0 3.9085e-08 0.0007 3.9088e-08 0 3.9282e-08 0 3.9285e-08 0.0007 3.9288e-08 0 3.9482e-08 0 3.9485e-08 0.0007 3.9488e-08 0 3.9682e-08 0 3.9685e-08 0.0007 3.9688e-08 0 3.9882e-08 0 3.9885e-08 0.0007 3.9888e-08 0 4.1682e-08 0 4.1685e-08 0.0007 4.1688e-08 0 4.1882e-08 0 4.1885e-08 0.0007 4.1888e-08 0 4.2082e-08 0 4.2085e-08 0.0007 4.2088e-08 0 4.2282e-08 0 4.2285e-08 0.0007 4.2288e-08 0 4.2482e-08 0 4.2485e-08 0.0007 4.2488e-08 0 4.2682e-08 0 4.2685e-08 0.0007 4.2688e-08 0 4.2882e-08 0 4.2885e-08 0.0007 4.2888e-08 0 4.3082e-08 0 4.3085e-08 0.0007 4.3088e-08 0 4.4882e-08 0 4.4885e-08 0.0007 4.4888e-08 0 4.5082e-08 0 4.5085e-08 0.0007 4.5088e-08 0 4.5282e-08 0 4.5285e-08 0.0007 4.5288e-08 0 4.5482e-08 0 4.5485e-08 0.0007 4.5488e-08 0 4.5682e-08 0 4.5685e-08 0.0007 4.5688e-08 0 4.5882e-08 0 4.5885e-08 0.0007 4.5888e-08 0 4.6082e-08 0 4.6085e-08 0.0007 4.6088e-08 0 4.6282e-08 0 4.6285e-08 0.0007 4.6288e-08 0 4.8082e-08 0 4.8085e-08 0.0007 4.8088e-08 0 4.8282e-08 0 4.8285e-08 0.0007 4.8288e-08 0 4.8482e-08 0 4.8485e-08 0.0007 4.8488e-08 0 4.8682e-08 0 4.8685e-08 0.0007 4.8688e-08 0 4.8882e-08 0 4.8885e-08 0.0007 4.8888e-08 0 4.9082e-08 0 4.9085e-08 0.0007 4.9088e-08 0 4.9282e-08 0 4.9285e-08 0.0007 4.9288e-08 0 4.9482e-08 0 4.9485e-08 0.0007 4.9488e-08 0)
IA2|E 0 A2  PWL(0 0 9.8e-11 0 1.01e-10 0.0007 1.04e-10 0 2.98e-10 0 3.01e-10 0.0007 3.04e-10 0 4.98e-10 0 5.01e-10 0.0007 5.04e-10 0 6.98e-10 0 7.01e-10 0.0007 7.04e-10 0 8.98e-10 0 9.01e-10 0.0007 9.04e-10 0 1.098e-09 0 1.101e-09 0.0007 1.104e-09 0 1.298e-09 0 1.301e-09 0.0007 1.304e-09 0 1.498e-09 0 1.501e-09 0.0007 1.504e-09 0 1.698e-09 0 1.701e-09 0.0007 1.704e-09 0 1.898e-09 0 1.901e-09 0.0007 1.904e-09 0 2.098e-09 0 2.101e-09 0.0007 2.104e-09 0 2.298e-09 0 2.301e-09 0.0007 2.304e-09 0 2.498e-09 0 2.501e-09 0.0007 2.504e-09 0 2.698e-09 0 2.701e-09 0.0007 2.704e-09 0 2.898e-09 0 2.901e-09 0.0007 2.904e-09 0 3.098e-09 0 3.101e-09 0.0007 3.104e-09 0 6.498e-09 0 6.501e-09 0.0007 6.504e-09 0 6.698e-09 0 6.701e-09 0.0007 6.704e-09 0 6.898e-09 0 6.901e-09 0.0007 6.904e-09 0 7.098e-09 0 7.101e-09 0.0007 7.104e-09 0 7.298e-09 0 7.301e-09 0.0007 7.304e-09 0 7.498e-09 0 7.501e-09 0.0007 7.504e-09 0 7.698e-09 0 7.701e-09 0.0007 7.704e-09 0 7.898e-09 0 7.901e-09 0.0007 7.904e-09 0 8.098e-09 0 8.101e-09 0.0007 8.104e-09 0 8.298e-09 0 8.301e-09 0.0007 8.304e-09 0 8.498e-09 0 8.501e-09 0.0007 8.504e-09 0 8.698e-09 0 8.701e-09 0.0007 8.704e-09 0 8.898e-09 0 8.901e-09 0.0007 8.904e-09 0 9.098e-09 0 9.101e-09 0.0007 9.104e-09 0 9.298e-09 0 9.301e-09 0.0007 9.304e-09 0 9.498e-09 0 9.501e-09 0.0007 9.504e-09 0 1.2898e-08 0 1.2901e-08 0.0007 1.2904e-08 0 1.3098e-08 0 1.3101e-08 0.0007 1.3104e-08 0 1.3298e-08 0 1.3301e-08 0.0007 1.3304e-08 0 1.3498e-08 0 1.3501e-08 0.0007 1.3504e-08 0 1.3698e-08 0 1.3701e-08 0.0007 1.3704e-08 0 1.3898e-08 0 1.3901e-08 0.0007 1.3904e-08 0 1.4098e-08 0 1.4101e-08 0.0007 1.4104e-08 0 1.4298e-08 0 1.4301e-08 0.0007 1.4304e-08 0 1.4498e-08 0 1.4501e-08 0.0007 1.4504e-08 0 1.4698e-08 0 1.4701e-08 0.0007 1.4704e-08 0 1.4898e-08 0 1.4901e-08 0.0007 1.4904e-08 0 1.5098e-08 0 1.5101e-08 0.0007 1.5104e-08 0 1.5298e-08 0 1.5301e-08 0.0007 1.5304e-08 0 1.5498e-08 0 1.5501e-08 0.0007 1.5504e-08 0 1.5698e-08 0 1.5701e-08 0.0007 1.5704e-08 0 1.5898e-08 0 1.5901e-08 0.0007 1.5904e-08 0 1.9298e-08 0 1.9301e-08 0.0007 1.9304e-08 0 1.9498e-08 0 1.9501e-08 0.0007 1.9504e-08 0 1.9698e-08 0 1.9701e-08 0.0007 1.9704e-08 0 1.9898e-08 0 1.9901e-08 0.0007 1.9904e-08 0 2.0098e-08 0 2.0101e-08 0.0007 2.0104e-08 0 2.0298e-08 0 2.0301e-08 0.0007 2.0304e-08 0 2.0498e-08 0 2.0501e-08 0.0007 2.0504e-08 0 2.0698e-08 0 2.0701e-08 0.0007 2.0704e-08 0 2.0898e-08 0 2.0901e-08 0.0007 2.0904e-08 0 2.1098e-08 0 2.1101e-08 0.0007 2.1104e-08 0 2.1298e-08 0 2.1301e-08 0.0007 2.1304e-08 0 2.1498e-08 0 2.1501e-08 0.0007 2.1504e-08 0 2.1698e-08 0 2.1701e-08 0.0007 2.1704e-08 0 2.1898e-08 0 2.1901e-08 0.0007 2.1904e-08 0 2.2098e-08 0 2.2101e-08 0.0007 2.2104e-08 0 2.2298e-08 0 2.2301e-08 0.0007 2.2304e-08 0 2.5698e-08 0 2.5701e-08 0.0007 2.5704e-08 0 2.5898e-08 0 2.5901e-08 0.0007 2.5904e-08 0 2.6098e-08 0 2.6101e-08 0.0007 2.6104e-08 0 2.6298e-08 0 2.6301e-08 0.0007 2.6304e-08 0 2.6498e-08 0 2.6501e-08 0.0007 2.6504e-08 0 2.6698e-08 0 2.6701e-08 0.0007 2.6704e-08 0 2.6898e-08 0 2.6901e-08 0.0007 2.6904e-08 0 2.7098e-08 0 2.7101e-08 0.0007 2.7104e-08 0 2.7298e-08 0 2.7301e-08 0.0007 2.7304e-08 0 2.7498e-08 0 2.7501e-08 0.0007 2.7504e-08 0 2.7698e-08 0 2.7701e-08 0.0007 2.7704e-08 0 2.7898e-08 0 2.7901e-08 0.0007 2.7904e-08 0 2.8098e-08 0 2.8101e-08 0.0007 2.8104e-08 0 2.8298e-08 0 2.8301e-08 0.0007 2.8304e-08 0 2.8498e-08 0 2.8501e-08 0.0007 2.8504e-08 0 2.8698e-08 0 2.8701e-08 0.0007 2.8704e-08 0 3.2098e-08 0 3.2101e-08 0.0007 3.2104e-08 0 3.2298e-08 0 3.2301e-08 0.0007 3.2304e-08 0 3.2498e-08 0 3.2501e-08 0.0007 3.2504e-08 0 3.2698e-08 0 3.2701e-08 0.0007 3.2704e-08 0 3.2898e-08 0 3.2901e-08 0.0007 3.2904e-08 0 3.3098e-08 0 3.3101e-08 0.0007 3.3104e-08 0 3.3298e-08 0 3.3301e-08 0.0007 3.3304e-08 0 3.3498e-08 0 3.3501e-08 0.0007 3.3504e-08 0 3.3698e-08 0 3.3701e-08 0.0007 3.3704e-08 0 3.3898e-08 0 3.3901e-08 0.0007 3.3904e-08 0 3.4098e-08 0 3.4101e-08 0.0007 3.4104e-08 0 3.4298e-08 0 3.4301e-08 0.0007 3.4304e-08 0 3.4498e-08 0 3.4501e-08 0.0007 3.4504e-08 0 3.4698e-08 0 3.4701e-08 0.0007 3.4704e-08 0 3.4898e-08 0 3.4901e-08 0.0007 3.4904e-08 0 3.5098e-08 0 3.5101e-08 0.0007 3.5104e-08 0 3.8498e-08 0 3.8501e-08 0.0007 3.8504e-08 0 3.8698e-08 0 3.8701e-08 0.0007 3.8704e-08 0 3.8898e-08 0 3.8901e-08 0.0007 3.8904e-08 0 3.9098e-08 0 3.9101e-08 0.0007 3.9104e-08 0 3.9298e-08 0 3.9301e-08 0.0007 3.9304e-08 0 3.9498e-08 0 3.9501e-08 0.0007 3.9504e-08 0 3.9698e-08 0 3.9701e-08 0.0007 3.9704e-08 0 3.9898e-08 0 3.9901e-08 0.0007 3.9904e-08 0 4.0098e-08 0 4.0101e-08 0.0007 4.0104e-08 0 4.0298e-08 0 4.0301e-08 0.0007 4.0304e-08 0 4.0498e-08 0 4.0501e-08 0.0007 4.0504e-08 0 4.0698e-08 0 4.0701e-08 0.0007 4.0704e-08 0 4.0898e-08 0 4.0901e-08 0.0007 4.0904e-08 0 4.1098e-08 0 4.1101e-08 0.0007 4.1104e-08 0 4.1298e-08 0 4.1301e-08 0.0007 4.1304e-08 0 4.1498e-08 0 4.1501e-08 0.0007 4.1504e-08 0 4.4898e-08 0 4.4901e-08 0.0007 4.4904e-08 0 4.5098e-08 0 4.5101e-08 0.0007 4.5104e-08 0 4.5298e-08 0 4.5301e-08 0.0007 4.5304e-08 0 4.5498e-08 0 4.5501e-08 0.0007 4.5504e-08 0 4.5698e-08 0 4.5701e-08 0.0007 4.5704e-08 0 4.5898e-08 0 4.5901e-08 0.0007 4.5904e-08 0 4.6098e-08 0 4.6101e-08 0.0007 4.6104e-08 0 4.6298e-08 0 4.6301e-08 0.0007 4.6304e-08 0 4.6498e-08 0 4.6501e-08 0.0007 4.6504e-08 0 4.6698e-08 0 4.6701e-08 0.0007 4.6704e-08 0 4.6898e-08 0 4.6901e-08 0.0007 4.6904e-08 0 4.7098e-08 0 4.7101e-08 0.0007 4.7104e-08 0 4.7298e-08 0 4.7301e-08 0.0007 4.7304e-08 0 4.7498e-08 0 4.7501e-08 0.0007 4.7504e-08 0 4.7698e-08 0 4.7701e-08 0.0007 4.7704e-08 0 4.7898e-08 0 4.7901e-08 0.0007 4.7904e-08 0)
IB2|F 0 B2  PWL(0 0 1.14e-10 0 1.17e-10 0.0007 1.2e-10 0 3.14e-10 0 3.17e-10 0.0007 3.2e-10 0 5.14e-10 0 5.17e-10 0.0007 5.2e-10 0 7.14e-10 0 7.17e-10 0.0007 7.2e-10 0 9.14e-10 0 9.17e-10 0.0007 9.2e-10 0 1.114e-09 0 1.117e-09 0.0007 1.12e-09 0 1.314e-09 0 1.317e-09 0.0007 1.32e-09 0 1.514e-09 0 1.517e-09 0.0007 1.52e-09 0 1.714e-09 0 1.717e-09 0.0007 1.72e-09 0 1.914e-09 0 1.917e-09 0.0007 1.92e-09 0 2.114e-09 0 2.117e-09 0.0007 2.12e-09 0 2.314e-09 0 2.317e-09 0.0007 2.32e-09 0 2.514e-09 0 2.517e-09 0.0007 2.52e-09 0 2.714e-09 0 2.717e-09 0.0007 2.72e-09 0 2.914e-09 0 2.917e-09 0.0007 2.92e-09 0 3.114e-09 0 3.117e-09 0.0007 3.12e-09 0 3.314e-09 0 3.317e-09 0.0007 3.32e-09 0 3.514e-09 0 3.517e-09 0.0007 3.52e-09 0 3.714e-09 0 3.717e-09 0.0007 3.72e-09 0 3.914e-09 0 3.917e-09 0.0007 3.92e-09 0 4.114e-09 0 4.117e-09 0.0007 4.12e-09 0 4.314e-09 0 4.317e-09 0.0007 4.32e-09 0 4.514e-09 0 4.517e-09 0.0007 4.52e-09 0 4.714e-09 0 4.717e-09 0.0007 4.72e-09 0 4.914e-09 0 4.917e-09 0.0007 4.92e-09 0 5.114e-09 0 5.117e-09 0.0007 5.12e-09 0 5.314e-09 0 5.317e-09 0.0007 5.32e-09 0 5.514e-09 0 5.517e-09 0.0007 5.52e-09 0 5.714e-09 0 5.717e-09 0.0007 5.72e-09 0 5.914e-09 0 5.917e-09 0.0007 5.92e-09 0 6.114e-09 0 6.117e-09 0.0007 6.12e-09 0 6.314e-09 0 6.317e-09 0.0007 6.32e-09 0 1.2914e-08 0 1.2917e-08 0.0007 1.292e-08 0 1.3114e-08 0 1.3117e-08 0.0007 1.312e-08 0 1.3314e-08 0 1.3317e-08 0.0007 1.332e-08 0 1.3514e-08 0 1.3517e-08 0.0007 1.352e-08 0 1.3714e-08 0 1.3717e-08 0.0007 1.372e-08 0 1.3914e-08 0 1.3917e-08 0.0007 1.392e-08 0 1.4114e-08 0 1.4117e-08 0.0007 1.412e-08 0 1.4314e-08 0 1.4317e-08 0.0007 1.432e-08 0 1.4514e-08 0 1.4517e-08 0.0007 1.452e-08 0 1.4714e-08 0 1.4717e-08 0.0007 1.472e-08 0 1.4914e-08 0 1.4917e-08 0.0007 1.492e-08 0 1.5114e-08 0 1.5117e-08 0.0007 1.512e-08 0 1.5314e-08 0 1.5317e-08 0.0007 1.532e-08 0 1.5514e-08 0 1.5517e-08 0.0007 1.552e-08 0 1.5714e-08 0 1.5717e-08 0.0007 1.572e-08 0 1.5914e-08 0 1.5917e-08 0.0007 1.592e-08 0 1.6114e-08 0 1.6117e-08 0.0007 1.612e-08 0 1.6314e-08 0 1.6317e-08 0.0007 1.632e-08 0 1.6514e-08 0 1.6517e-08 0.0007 1.652e-08 0 1.6714e-08 0 1.6717e-08 0.0007 1.672e-08 0 1.6914e-08 0 1.6917e-08 0.0007 1.692e-08 0 1.7114e-08 0 1.7117e-08 0.0007 1.712e-08 0 1.7314e-08 0 1.7317e-08 0.0007 1.732e-08 0 1.7514e-08 0 1.7517e-08 0.0007 1.752e-08 0 1.7714e-08 0 1.7717e-08 0.0007 1.772e-08 0 1.7914e-08 0 1.7917e-08 0.0007 1.792e-08 0 1.8114e-08 0 1.8117e-08 0.0007 1.812e-08 0 1.8314e-08 0 1.8317e-08 0.0007 1.832e-08 0 1.8514e-08 0 1.8517e-08 0.0007 1.852e-08 0 1.8714e-08 0 1.8717e-08 0.0007 1.872e-08 0 1.8914e-08 0 1.8917e-08 0.0007 1.892e-08 0 1.9114e-08 0 1.9117e-08 0.0007 1.912e-08 0 2.5714e-08 0 2.5717e-08 0.0007 2.572e-08 0 2.5914e-08 0 2.5917e-08 0.0007 2.592e-08 0 2.6114e-08 0 2.6117e-08 0.0007 2.612e-08 0 2.6314e-08 0 2.6317e-08 0.0007 2.632e-08 0 2.6514e-08 0 2.6517e-08 0.0007 2.652e-08 0 2.6714e-08 0 2.6717e-08 0.0007 2.672e-08 0 2.6914e-08 0 2.6917e-08 0.0007 2.692e-08 0 2.7114e-08 0 2.7117e-08 0.0007 2.712e-08 0 2.7314e-08 0 2.7317e-08 0.0007 2.732e-08 0 2.7514e-08 0 2.7517e-08 0.0007 2.752e-08 0 2.7714e-08 0 2.7717e-08 0.0007 2.772e-08 0 2.7914e-08 0 2.7917e-08 0.0007 2.792e-08 0 2.8114e-08 0 2.8117e-08 0.0007 2.812e-08 0 2.8314e-08 0 2.8317e-08 0.0007 2.832e-08 0 2.8514e-08 0 2.8517e-08 0.0007 2.852e-08 0 2.8714e-08 0 2.8717e-08 0.0007 2.872e-08 0 2.8914e-08 0 2.8917e-08 0.0007 2.892e-08 0 2.9114e-08 0 2.9117e-08 0.0007 2.912e-08 0 2.9314e-08 0 2.9317e-08 0.0007 2.932e-08 0 2.9514e-08 0 2.9517e-08 0.0007 2.952e-08 0 2.9714e-08 0 2.9717e-08 0.0007 2.972e-08 0 2.9914e-08 0 2.9917e-08 0.0007 2.992e-08 0 3.0114e-08 0 3.0117e-08 0.0007 3.012e-08 0 3.0314e-08 0 3.0317e-08 0.0007 3.032e-08 0 3.0514e-08 0 3.0517e-08 0.0007 3.052e-08 0 3.0714e-08 0 3.0717e-08 0.0007 3.072e-08 0 3.0914e-08 0 3.0917e-08 0.0007 3.092e-08 0 3.1114e-08 0 3.1117e-08 0.0007 3.112e-08 0 3.1314e-08 0 3.1317e-08 0.0007 3.132e-08 0 3.1514e-08 0 3.1517e-08 0.0007 3.152e-08 0 3.1714e-08 0 3.1717e-08 0.0007 3.172e-08 0 3.1914e-08 0 3.1917e-08 0.0007 3.192e-08 0 3.8514e-08 0 3.8517e-08 0.0007 3.852e-08 0 3.8714e-08 0 3.8717e-08 0.0007 3.872e-08 0 3.8914e-08 0 3.8917e-08 0.0007 3.892e-08 0 3.9114e-08 0 3.9117e-08 0.0007 3.912e-08 0 3.9314e-08 0 3.9317e-08 0.0007 3.932e-08 0 3.9514e-08 0 3.9517e-08 0.0007 3.952e-08 0 3.9714e-08 0 3.9717e-08 0.0007 3.972e-08 0 3.9914e-08 0 3.9917e-08 0.0007 3.992e-08 0 4.0114e-08 0 4.0117e-08 0.0007 4.012e-08 0 4.0314e-08 0 4.0317e-08 0.0007 4.032e-08 0 4.0514e-08 0 4.0517e-08 0.0007 4.052e-08 0 4.0714e-08 0 4.0717e-08 0.0007 4.072e-08 0 4.0914e-08 0 4.0917e-08 0.0007 4.092e-08 0 4.1114e-08 0 4.1117e-08 0.0007 4.112e-08 0 4.1314e-08 0 4.1317e-08 0.0007 4.132e-08 0 4.1514e-08 0 4.1517e-08 0.0007 4.152e-08 0 4.1714e-08 0 4.1717e-08 0.0007 4.172e-08 0 4.1914e-08 0 4.1917e-08 0.0007 4.192e-08 0 4.2114e-08 0 4.2117e-08 0.0007 4.212e-08 0 4.2314e-08 0 4.2317e-08 0.0007 4.232e-08 0 4.2514e-08 0 4.2517e-08 0.0007 4.252e-08 0 4.2714e-08 0 4.2717e-08 0.0007 4.272e-08 0 4.2914e-08 0 4.2917e-08 0.0007 4.292e-08 0 4.3114e-08 0 4.3117e-08 0.0007 4.312e-08 0 4.3314e-08 0 4.3317e-08 0.0007 4.332e-08 0 4.3514e-08 0 4.3517e-08 0.0007 4.352e-08 0 4.3714e-08 0 4.3717e-08 0.0007 4.372e-08 0 4.3914e-08 0 4.3917e-08 0.0007 4.392e-08 0 4.4114e-08 0 4.4117e-08 0.0007 4.412e-08 0 4.4314e-08 0 4.4317e-08 0.0007 4.432e-08 0 4.4514e-08 0 4.4517e-08 0.0007 4.452e-08 0 4.4714e-08 0 4.4717e-08 0.0007 4.472e-08 0)
IA3|G 0 A3  PWL(0 0 1.3e-10 0 1.33e-10 0.0007 1.36e-10 0 3.3e-10 0 3.33e-10 0.0007 3.36e-10 0 5.3e-10 0 5.33e-10 0.0007 5.36e-10 0 7.3e-10 0 7.33e-10 0.0007 7.36e-10 0 9.3e-10 0 9.33e-10 0.0007 9.36e-10 0 1.13e-09 0 1.133e-09 0.0007 1.136e-09 0 1.33e-09 0 1.333e-09 0.0007 1.336e-09 0 1.53e-09 0 1.533e-09 0.0007 1.536e-09 0 1.73e-09 0 1.733e-09 0.0007 1.736e-09 0 1.93e-09 0 1.933e-09 0.0007 1.936e-09 0 2.13e-09 0 2.133e-09 0.0007 2.136e-09 0 2.33e-09 0 2.333e-09 0.0007 2.336e-09 0 2.53e-09 0 2.533e-09 0.0007 2.536e-09 0 2.73e-09 0 2.733e-09 0.0007 2.736e-09 0 2.93e-09 0 2.933e-09 0.0007 2.936e-09 0 3.13e-09 0 3.133e-09 0.0007 3.136e-09 0 3.33e-09 0 3.333e-09 0.0007 3.336e-09 0 3.53e-09 0 3.533e-09 0.0007 3.536e-09 0 3.73e-09 0 3.733e-09 0.0007 3.736e-09 0 3.93e-09 0 3.933e-09 0.0007 3.936e-09 0 4.13e-09 0 4.133e-09 0.0007 4.136e-09 0 4.33e-09 0 4.333e-09 0.0007 4.336e-09 0 4.53e-09 0 4.533e-09 0.0007 4.536e-09 0 4.73e-09 0 4.733e-09 0.0007 4.736e-09 0 4.93e-09 0 4.933e-09 0.0007 4.936e-09 0 5.13e-09 0 5.133e-09 0.0007 5.136e-09 0 5.33e-09 0 5.333e-09 0.0007 5.336e-09 0 5.53e-09 0 5.533e-09 0.0007 5.536e-09 0 5.73e-09 0 5.733e-09 0.0007 5.736e-09 0 5.93e-09 0 5.933e-09 0.0007 5.936e-09 0 6.13e-09 0 6.133e-09 0.0007 6.136e-09 0 6.33e-09 0 6.333e-09 0.0007 6.336e-09 0 6.53e-09 0 6.533e-09 0.0007 6.536e-09 0 6.73e-09 0 6.733e-09 0.0007 6.736e-09 0 6.93e-09 0 6.933e-09 0.0007 6.936e-09 0 7.13e-09 0 7.133e-09 0.0007 7.136e-09 0 7.33e-09 0 7.333e-09 0.0007 7.336e-09 0 7.53e-09 0 7.533e-09 0.0007 7.536e-09 0 7.73e-09 0 7.733e-09 0.0007 7.736e-09 0 7.93e-09 0 7.933e-09 0.0007 7.936e-09 0 8.13e-09 0 8.133e-09 0.0007 8.136e-09 0 8.33e-09 0 8.333e-09 0.0007 8.336e-09 0 8.53e-09 0 8.533e-09 0.0007 8.536e-09 0 8.73e-09 0 8.733e-09 0.0007 8.736e-09 0 8.93e-09 0 8.933e-09 0.0007 8.936e-09 0 9.13e-09 0 9.133e-09 0.0007 9.136e-09 0 9.33e-09 0 9.333e-09 0.0007 9.336e-09 0 9.53e-09 0 9.533e-09 0.0007 9.536e-09 0 9.73e-09 0 9.733e-09 0.0007 9.736e-09 0 9.93e-09 0 9.933e-09 0.0007 9.936e-09 0 1.013e-08 0 1.0133e-08 0.0007 1.0136e-08 0 1.033e-08 0 1.0333e-08 0.0007 1.0336e-08 0 1.053e-08 0 1.0533e-08 0.0007 1.0536e-08 0 1.073e-08 0 1.0733e-08 0.0007 1.0736e-08 0 1.093e-08 0 1.0933e-08 0.0007 1.0936e-08 0 1.113e-08 0 1.1133e-08 0.0007 1.1136e-08 0 1.133e-08 0 1.1333e-08 0.0007 1.1336e-08 0 1.153e-08 0 1.1533e-08 0.0007 1.1536e-08 0 1.173e-08 0 1.1733e-08 0.0007 1.1736e-08 0 1.193e-08 0 1.1933e-08 0.0007 1.1936e-08 0 1.213e-08 0 1.2133e-08 0.0007 1.2136e-08 0 1.233e-08 0 1.2333e-08 0.0007 1.2336e-08 0 1.253e-08 0 1.2533e-08 0.0007 1.2536e-08 0 1.273e-08 0 1.2733e-08 0.0007 1.2736e-08 0 2.573e-08 0 2.5733e-08 0.0007 2.5736e-08 0 2.593e-08 0 2.5933e-08 0.0007 2.5936e-08 0 2.613e-08 0 2.6133e-08 0.0007 2.6136e-08 0 2.633e-08 0 2.6333e-08 0.0007 2.6336e-08 0 2.653e-08 0 2.6533e-08 0.0007 2.6536e-08 0 2.673e-08 0 2.6733e-08 0.0007 2.6736e-08 0 2.693e-08 0 2.6933e-08 0.0007 2.6936e-08 0 2.713e-08 0 2.7133e-08 0.0007 2.7136e-08 0 2.733e-08 0 2.7333e-08 0.0007 2.7336e-08 0 2.753e-08 0 2.7533e-08 0.0007 2.7536e-08 0 2.773e-08 0 2.7733e-08 0.0007 2.7736e-08 0 2.793e-08 0 2.7933e-08 0.0007 2.7936e-08 0 2.813e-08 0 2.8133e-08 0.0007 2.8136e-08 0 2.833e-08 0 2.8333e-08 0.0007 2.8336e-08 0 2.853e-08 0 2.8533e-08 0.0007 2.8536e-08 0 2.873e-08 0 2.8733e-08 0.0007 2.8736e-08 0 2.893e-08 0 2.8933e-08 0.0007 2.8936e-08 0 2.913e-08 0 2.9133e-08 0.0007 2.9136e-08 0 2.933e-08 0 2.9333e-08 0.0007 2.9336e-08 0 2.953e-08 0 2.9533e-08 0.0007 2.9536e-08 0 2.973e-08 0 2.9733e-08 0.0007 2.9736e-08 0 2.993e-08 0 2.9933e-08 0.0007 2.9936e-08 0 3.013e-08 0 3.0133e-08 0.0007 3.0136e-08 0 3.033e-08 0 3.0333e-08 0.0007 3.0336e-08 0 3.053e-08 0 3.0533e-08 0.0007 3.0536e-08 0 3.073e-08 0 3.0733e-08 0.0007 3.0736e-08 0 3.093e-08 0 3.0933e-08 0.0007 3.0936e-08 0 3.113e-08 0 3.1133e-08 0.0007 3.1136e-08 0 3.133e-08 0 3.1333e-08 0.0007 3.1336e-08 0 3.153e-08 0 3.1533e-08 0.0007 3.1536e-08 0 3.173e-08 0 3.1733e-08 0.0007 3.1736e-08 0 3.193e-08 0 3.1933e-08 0.0007 3.1936e-08 0 3.213e-08 0 3.2133e-08 0.0007 3.2136e-08 0 3.233e-08 0 3.2333e-08 0.0007 3.2336e-08 0 3.253e-08 0 3.2533e-08 0.0007 3.2536e-08 0 3.273e-08 0 3.2733e-08 0.0007 3.2736e-08 0 3.293e-08 0 3.2933e-08 0.0007 3.2936e-08 0 3.313e-08 0 3.3133e-08 0.0007 3.3136e-08 0 3.333e-08 0 3.3333e-08 0.0007 3.3336e-08 0 3.353e-08 0 3.3533e-08 0.0007 3.3536e-08 0 3.373e-08 0 3.3733e-08 0.0007 3.3736e-08 0 3.393e-08 0 3.3933e-08 0.0007 3.3936e-08 0 3.413e-08 0 3.4133e-08 0.0007 3.4136e-08 0 3.433e-08 0 3.4333e-08 0.0007 3.4336e-08 0 3.453e-08 0 3.4533e-08 0.0007 3.4536e-08 0 3.473e-08 0 3.4733e-08 0.0007 3.4736e-08 0 3.493e-08 0 3.4933e-08 0.0007 3.4936e-08 0 3.513e-08 0 3.5133e-08 0.0007 3.5136e-08 0 3.533e-08 0 3.5333e-08 0.0007 3.5336e-08 0 3.553e-08 0 3.5533e-08 0.0007 3.5536e-08 0 3.573e-08 0 3.5733e-08 0.0007 3.5736e-08 0 3.593e-08 0 3.5933e-08 0.0007 3.5936e-08 0 3.613e-08 0 3.6133e-08 0.0007 3.6136e-08 0 3.633e-08 0 3.6333e-08 0.0007 3.6336e-08 0 3.653e-08 0 3.6533e-08 0.0007 3.6536e-08 0 3.673e-08 0 3.6733e-08 0.0007 3.6736e-08 0 3.693e-08 0 3.6933e-08 0.0007 3.6936e-08 0 3.713e-08 0 3.7133e-08 0.0007 3.7136e-08 0 3.733e-08 0 3.7333e-08 0.0007 3.7336e-08 0 3.753e-08 0 3.7533e-08 0.0007 3.7536e-08 0 3.773e-08 0 3.7733e-08 0.0007 3.7736e-08 0 3.793e-08 0 3.7933e-08 0.0007 3.7936e-08 0 3.813e-08 0 3.8133e-08 0.0007 3.8136e-08 0 3.833e-08 0 3.8333e-08 0.0007 3.8336e-08 0)
IB3|H 0 B3  PWL(0 0 1.46e-10 0 1.49e-10 0.0007 1.52e-10 0 3.46e-10 0 3.49e-10 0.0007 3.52e-10 0 5.46e-10 0 5.49e-10 0.0007 5.52e-10 0 7.46e-10 0 7.49e-10 0.0007 7.52e-10 0 9.46e-10 0 9.49e-10 0.0007 9.52e-10 0 1.146e-09 0 1.149e-09 0.0007 1.152e-09 0 1.346e-09 0 1.349e-09 0.0007 1.352e-09 0 1.546e-09 0 1.549e-09 0.0007 1.552e-09 0 1.746e-09 0 1.749e-09 0.0007 1.752e-09 0 1.946e-09 0 1.949e-09 0.0007 1.952e-09 0 2.146e-09 0 2.149e-09 0.0007 2.152e-09 0 2.346e-09 0 2.349e-09 0.0007 2.352e-09 0 2.546e-09 0 2.549e-09 0.0007 2.552e-09 0 2.746e-09 0 2.749e-09 0.0007 2.752e-09 0 2.946e-09 0 2.949e-09 0.0007 2.952e-09 0 3.146e-09 0 3.149e-09 0.0007 3.152e-09 0 3.346e-09 0 3.349e-09 0.0007 3.352e-09 0 3.546e-09 0 3.549e-09 0.0007 3.552e-09 0 3.746e-09 0 3.749e-09 0.0007 3.752e-09 0 3.946e-09 0 3.949e-09 0.0007 3.952e-09 0 4.146e-09 0 4.149e-09 0.0007 4.152e-09 0 4.346e-09 0 4.349e-09 0.0007 4.352e-09 0 4.546e-09 0 4.549e-09 0.0007 4.552e-09 0 4.746e-09 0 4.749e-09 0.0007 4.752e-09 0 4.946e-09 0 4.949e-09 0.0007 4.952e-09 0 5.146e-09 0 5.149e-09 0.0007 5.152e-09 0 5.346e-09 0 5.349e-09 0.0007 5.352e-09 0 5.546e-09 0 5.549e-09 0.0007 5.552e-09 0 5.746e-09 0 5.749e-09 0.0007 5.752e-09 0 5.946e-09 0 5.949e-09 0.0007 5.952e-09 0 6.146e-09 0 6.149e-09 0.0007 6.152e-09 0 6.346e-09 0 6.349e-09 0.0007 6.352e-09 0 6.546e-09 0 6.549e-09 0.0007 6.552e-09 0 6.746e-09 0 6.749e-09 0.0007 6.752e-09 0 6.946e-09 0 6.949e-09 0.0007 6.952e-09 0 7.146e-09 0 7.149e-09 0.0007 7.152e-09 0 7.346e-09 0 7.349e-09 0.0007 7.352e-09 0 7.546e-09 0 7.549e-09 0.0007 7.552e-09 0 7.746e-09 0 7.749e-09 0.0007 7.752e-09 0 7.946e-09 0 7.949e-09 0.0007 7.952e-09 0 8.146e-09 0 8.149e-09 0.0007 8.152e-09 0 8.346e-09 0 8.349e-09 0.0007 8.352e-09 0 8.546e-09 0 8.549e-09 0.0007 8.552e-09 0 8.746e-09 0 8.749e-09 0.0007 8.752e-09 0 8.946e-09 0 8.949e-09 0.0007 8.952e-09 0 9.146e-09 0 9.149e-09 0.0007 9.152e-09 0 9.346e-09 0 9.349e-09 0.0007 9.352e-09 0 9.546e-09 0 9.549e-09 0.0007 9.552e-09 0 9.746e-09 0 9.749e-09 0.0007 9.752e-09 0 9.946e-09 0 9.949e-09 0.0007 9.952e-09 0 1.0146e-08 0 1.0149e-08 0.0007 1.0152e-08 0 1.0346e-08 0 1.0349e-08 0.0007 1.0352e-08 0 1.0546e-08 0 1.0549e-08 0.0007 1.0552e-08 0 1.0746e-08 0 1.0749e-08 0.0007 1.0752e-08 0 1.0946e-08 0 1.0949e-08 0.0007 1.0952e-08 0 1.1146e-08 0 1.1149e-08 0.0007 1.1152e-08 0 1.1346e-08 0 1.1349e-08 0.0007 1.1352e-08 0 1.1546e-08 0 1.1549e-08 0.0007 1.1552e-08 0 1.1746e-08 0 1.1749e-08 0.0007 1.1752e-08 0 1.1946e-08 0 1.1949e-08 0.0007 1.1952e-08 0 1.2146e-08 0 1.2149e-08 0.0007 1.2152e-08 0 1.2346e-08 0 1.2349e-08 0.0007 1.2352e-08 0 1.2546e-08 0 1.2549e-08 0.0007 1.2552e-08 0 1.2746e-08 0 1.2749e-08 0.0007 1.2752e-08 0 1.2946e-08 0 1.2949e-08 0.0007 1.2952e-08 0 1.3146e-08 0 1.3149e-08 0.0007 1.3152e-08 0 1.3346e-08 0 1.3349e-08 0.0007 1.3352e-08 0 1.3546e-08 0 1.3549e-08 0.0007 1.3552e-08 0 1.3746e-08 0 1.3749e-08 0.0007 1.3752e-08 0 1.3946e-08 0 1.3949e-08 0.0007 1.3952e-08 0 1.4146e-08 0 1.4149e-08 0.0007 1.4152e-08 0 1.4346e-08 0 1.4349e-08 0.0007 1.4352e-08 0 1.4546e-08 0 1.4549e-08 0.0007 1.4552e-08 0 1.4746e-08 0 1.4749e-08 0.0007 1.4752e-08 0 1.4946e-08 0 1.4949e-08 0.0007 1.4952e-08 0 1.5146e-08 0 1.5149e-08 0.0007 1.5152e-08 0 1.5346e-08 0 1.5349e-08 0.0007 1.5352e-08 0 1.5546e-08 0 1.5549e-08 0.0007 1.5552e-08 0 1.5746e-08 0 1.5749e-08 0.0007 1.5752e-08 0 1.5946e-08 0 1.5949e-08 0.0007 1.5952e-08 0 1.6146e-08 0 1.6149e-08 0.0007 1.6152e-08 0 1.6346e-08 0 1.6349e-08 0.0007 1.6352e-08 0 1.6546e-08 0 1.6549e-08 0.0007 1.6552e-08 0 1.6746e-08 0 1.6749e-08 0.0007 1.6752e-08 0 1.6946e-08 0 1.6949e-08 0.0007 1.6952e-08 0 1.7146e-08 0 1.7149e-08 0.0007 1.7152e-08 0 1.7346e-08 0 1.7349e-08 0.0007 1.7352e-08 0 1.7546e-08 0 1.7549e-08 0.0007 1.7552e-08 0 1.7746e-08 0 1.7749e-08 0.0007 1.7752e-08 0 1.7946e-08 0 1.7949e-08 0.0007 1.7952e-08 0 1.8146e-08 0 1.8149e-08 0.0007 1.8152e-08 0 1.8346e-08 0 1.8349e-08 0.0007 1.8352e-08 0 1.8546e-08 0 1.8549e-08 0.0007 1.8552e-08 0 1.8746e-08 0 1.8749e-08 0.0007 1.8752e-08 0 1.8946e-08 0 1.8949e-08 0.0007 1.8952e-08 0 1.9146e-08 0 1.9149e-08 0.0007 1.9152e-08 0 1.9346e-08 0 1.9349e-08 0.0007 1.9352e-08 0 1.9546e-08 0 1.9549e-08 0.0007 1.9552e-08 0 1.9746e-08 0 1.9749e-08 0.0007 1.9752e-08 0 1.9946e-08 0 1.9949e-08 0.0007 1.9952e-08 0 2.0146e-08 0 2.0149e-08 0.0007 2.0152e-08 0 2.0346e-08 0 2.0349e-08 0.0007 2.0352e-08 0 2.0546e-08 0 2.0549e-08 0.0007 2.0552e-08 0 2.0746e-08 0 2.0749e-08 0.0007 2.0752e-08 0 2.0946e-08 0 2.0949e-08 0.0007 2.0952e-08 0 2.1146e-08 0 2.1149e-08 0.0007 2.1152e-08 0 2.1346e-08 0 2.1349e-08 0.0007 2.1352e-08 0 2.1546e-08 0 2.1549e-08 0.0007 2.1552e-08 0 2.1746e-08 0 2.1749e-08 0.0007 2.1752e-08 0 2.1946e-08 0 2.1949e-08 0.0007 2.1952e-08 0 2.2146e-08 0 2.2149e-08 0.0007 2.2152e-08 0 2.2346e-08 0 2.2349e-08 0.0007 2.2352e-08 0 2.2546e-08 0 2.2549e-08 0.0007 2.2552e-08 0 2.2746e-08 0 2.2749e-08 0.0007 2.2752e-08 0 2.2946e-08 0 2.2949e-08 0.0007 2.2952e-08 0 2.3146e-08 0 2.3149e-08 0.0007 2.3152e-08 0 2.3346e-08 0 2.3349e-08 0.0007 2.3352e-08 0 2.3546e-08 0 2.3549e-08 0.0007 2.3552e-08 0 2.3746e-08 0 2.3749e-08 0.0007 2.3752e-08 0 2.3946e-08 0 2.3949e-08 0.0007 2.3952e-08 0 2.4146e-08 0 2.4149e-08 0.0007 2.4152e-08 0 2.4346e-08 0 2.4349e-08 0.0007 2.4352e-08 0 2.4546e-08 0 2.4549e-08 0.0007 2.4552e-08 0 2.4746e-08 0 2.4749e-08 0.0007 2.4752e-08 0 2.4946e-08 0 2.4949e-08 0.0007 2.4952e-08 0 2.5146e-08 0 2.5149e-08 0.0007 2.5152e-08 0 2.5346e-08 0 2.5349e-08 0.0007 2.5352e-08 0 2.5546e-08 0 2.5549e-08 0.0007 2.5552e-08 0)
IT00|T 0 T00  PWL(0 0 1.7e-11 0 2e-11 0.0021 2.3e-11 0 2.17e-10 0 2.2e-10 0.0021 2.23e-10 0 4.17e-10 0 4.2e-10 0.0021 4.23e-10 0 6.17e-10 0 6.2e-10 0.0021 6.23e-10 0 8.17e-10 0 8.2e-10 0.0021 8.23e-10 0 1.017e-09 0 1.02e-09 0.0021 1.023e-09 0 1.217e-09 0 1.22e-09 0.0021 1.223e-09 0 1.417e-09 0 1.42e-09 0.0021 1.423e-09 0 1.617e-09 0 1.62e-09 0.0021 1.623e-09 0 1.817e-09 0 1.82e-09 0.0021 1.823e-09 0 2.017e-09 0 2.02e-09 0.0021 2.023e-09 0 2.217e-09 0 2.22e-09 0.0021 2.223e-09 0 2.417e-09 0 2.42e-09 0.0021 2.423e-09 0 2.617e-09 0 2.62e-09 0.0021 2.623e-09 0 2.817e-09 0 2.82e-09 0.0021 2.823e-09 0 3.017e-09 0 3.02e-09 0.0021 3.023e-09 0 3.217e-09 0 3.22e-09 0.0021 3.223e-09 0 3.417e-09 0 3.42e-09 0.0021 3.423e-09 0 3.617e-09 0 3.62e-09 0.0021 3.623e-09 0 3.817e-09 0 3.82e-09 0.0021 3.823e-09 0 4.017e-09 0 4.02e-09 0.0021 4.023e-09 0 4.217e-09 0 4.22e-09 0.0021 4.223e-09 0 4.417e-09 0 4.42e-09 0.0021 4.423e-09 0 4.617e-09 0 4.62e-09 0.0021 4.623e-09 0 4.817e-09 0 4.82e-09 0.0021 4.823e-09 0 5.017e-09 0 5.02e-09 0.0021 5.023e-09 0 5.217e-09 0 5.22e-09 0.0021 5.223e-09 0 5.417e-09 0 5.42e-09 0.0021 5.423e-09 0 5.617e-09 0 5.62e-09 0.0021 5.623e-09 0 5.817e-09 0 5.82e-09 0.0021 5.823e-09 0 6.017e-09 0 6.02e-09 0.0021 6.023e-09 0 6.217e-09 0 6.22e-09 0.0021 6.223e-09 0 6.417e-09 0 6.42e-09 0.0021 6.423e-09 0 6.617e-09 0 6.62e-09 0.0021 6.623e-09 0 6.817e-09 0 6.82e-09 0.0021 6.823e-09 0 7.017e-09 0 7.02e-09 0.0021 7.023e-09 0 7.217e-09 0 7.22e-09 0.0021 7.223e-09 0 7.417e-09 0 7.42e-09 0.0021 7.423e-09 0 7.617e-09 0 7.62e-09 0.0021 7.623e-09 0 7.817e-09 0 7.82e-09 0.0021 7.823e-09 0 8.017e-09 0 8.02e-09 0.0021 8.023e-09 0 8.217e-09 0 8.22e-09 0.0021 8.223e-09 0 8.417e-09 0 8.42e-09 0.0021 8.423e-09 0 8.617e-09 0 8.62e-09 0.0021 8.623e-09 0 8.817e-09 0 8.82e-09 0.0021 8.823e-09 0 9.017e-09 0 9.02e-09 0.0021 9.023e-09 0 9.217e-09 0 9.22e-09 0.0021 9.223e-09 0 9.417e-09 0 9.42e-09 0.0021 9.423e-09 0 9.617e-09 0 9.62e-09 0.0021 9.623e-09 0 9.817e-09 0 9.82e-09 0.0021 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0021 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0021 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0021 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0021 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0021 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0021 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0021 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0021 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0021 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0021 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0021 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0021 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0021 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0021 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0021 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0021 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0021 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0021 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0021 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0021 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0021 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0021 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0021 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0021 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0021 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0021 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0021 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0021 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0021 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0021 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0021 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0021 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0021 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0021 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0021 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0021 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0021 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0021 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0021 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0021 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0021 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0021 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0021 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0021 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0021 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0021 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0021 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0021 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0021 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0021 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0021 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0021 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0021 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0021 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0021 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0021 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0021 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0021 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0021 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0021 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0021 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0021 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0021 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0021 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0021 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0021 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0021 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0021 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0021 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0021 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0021 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0021 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0021 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0021 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0021 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0021 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0021 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0021 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0021 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0021 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0021 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0021 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0021 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0021 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0021 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0021 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0021 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0021 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0021 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0021 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0021 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0021 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0021 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0021 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0021 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0021 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0021 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0021 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0021 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0021 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0021 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0021 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0021 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0021 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0021 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0021 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0021 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0021 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0021 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0021 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0021 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0021 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0021 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0021 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0021 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0021 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0021 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0021 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0021 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0021 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0021 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0021 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0021 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0021 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0021 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0021 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0021 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0021 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0021 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0021 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0021 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0021 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0021 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0021 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0021 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0021 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0021 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0021 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0021 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0021 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0021 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0021 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0021 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0021 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0021 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0021 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0021 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0021 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0021 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0021 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0021 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0021 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0021 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0021 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0021 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0021 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0021 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0021 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0021 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0021 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0021 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0021 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0021 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0021 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0021 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0021 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0021 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0021 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0021 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0021 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0021 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0021 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0021 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0021 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0021 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0021 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0021 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0021 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0021 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0021 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0021 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0021 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0021 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0021 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0021 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0021 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0021 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0021 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0021 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0021 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0021 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0021 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0021 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0021 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0021 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0021 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0021 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0021 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0021 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0021 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0021 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0021 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0021 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0021 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0021 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0021 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0021 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0021 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0021 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0021 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0021 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0021 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0021 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0021 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0021 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0021 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0021 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0021 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0021 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0021 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0021 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0021 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0021 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0021 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0021 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0021 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0021 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0021 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0021 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0021 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0021 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0021 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0021 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0021 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0021 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0021 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0021 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0021 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0021 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0021 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0021 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0021 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0021 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0021 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0021 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0021 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0021 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0021 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0021 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0021 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0021 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0021 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0021 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0021 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0021 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0021 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0021 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0021 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0021 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0021 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0021 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0021 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0021 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0021 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0021 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0021 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0021 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0021 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0021 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0021 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0021 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0021 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0021 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0021 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0021 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0021 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0021 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0021 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0021 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0021 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0021 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0021 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0021 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0021 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0021 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0021 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0021 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0021 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0021 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0021 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0021 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0021 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0021 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0021 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0021 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0021 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0021 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0021 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0021 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0021 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0021 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0021 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0021 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0021 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0021 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0021 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0021 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0021 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0021 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0021 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0021 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0021 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0021 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0021 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0021 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0021 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0021 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0021 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0021 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0021 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0021 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0021 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0021 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0021 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0021 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0021 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0021 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0021 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0021 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0021 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0021 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0021 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0021 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0021 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0021 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0021 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0021 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0021 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0021 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0021 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0021 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0021 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0021 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0021 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0021 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0021 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0021 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0021 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0021 7.9623e-08 0)
IT01|T 0 T01  PWL(0 0 1.7e-11 0 2e-11 0.0021 2.3e-11 0 2.17e-10 0 2.2e-10 0.0021 2.23e-10 0 4.17e-10 0 4.2e-10 0.0021 4.23e-10 0 6.17e-10 0 6.2e-10 0.0021 6.23e-10 0 8.17e-10 0 8.2e-10 0.0021 8.23e-10 0 1.017e-09 0 1.02e-09 0.0021 1.023e-09 0 1.217e-09 0 1.22e-09 0.0021 1.223e-09 0 1.417e-09 0 1.42e-09 0.0021 1.423e-09 0 1.617e-09 0 1.62e-09 0.0021 1.623e-09 0 1.817e-09 0 1.82e-09 0.0021 1.823e-09 0 2.017e-09 0 2.02e-09 0.0021 2.023e-09 0 2.217e-09 0 2.22e-09 0.0021 2.223e-09 0 2.417e-09 0 2.42e-09 0.0021 2.423e-09 0 2.617e-09 0 2.62e-09 0.0021 2.623e-09 0 2.817e-09 0 2.82e-09 0.0021 2.823e-09 0 3.017e-09 0 3.02e-09 0.0021 3.023e-09 0 3.217e-09 0 3.22e-09 0.0021 3.223e-09 0 3.417e-09 0 3.42e-09 0.0021 3.423e-09 0 3.617e-09 0 3.62e-09 0.0021 3.623e-09 0 3.817e-09 0 3.82e-09 0.0021 3.823e-09 0 4.017e-09 0 4.02e-09 0.0021 4.023e-09 0 4.217e-09 0 4.22e-09 0.0021 4.223e-09 0 4.417e-09 0 4.42e-09 0.0021 4.423e-09 0 4.617e-09 0 4.62e-09 0.0021 4.623e-09 0 4.817e-09 0 4.82e-09 0.0021 4.823e-09 0 5.017e-09 0 5.02e-09 0.0021 5.023e-09 0 5.217e-09 0 5.22e-09 0.0021 5.223e-09 0 5.417e-09 0 5.42e-09 0.0021 5.423e-09 0 5.617e-09 0 5.62e-09 0.0021 5.623e-09 0 5.817e-09 0 5.82e-09 0.0021 5.823e-09 0 6.017e-09 0 6.02e-09 0.0021 6.023e-09 0 6.217e-09 0 6.22e-09 0.0021 6.223e-09 0 6.417e-09 0 6.42e-09 0.0021 6.423e-09 0 6.617e-09 0 6.62e-09 0.0021 6.623e-09 0 6.817e-09 0 6.82e-09 0.0021 6.823e-09 0 7.017e-09 0 7.02e-09 0.0021 7.023e-09 0 7.217e-09 0 7.22e-09 0.0021 7.223e-09 0 7.417e-09 0 7.42e-09 0.0021 7.423e-09 0 7.617e-09 0 7.62e-09 0.0021 7.623e-09 0 7.817e-09 0 7.82e-09 0.0021 7.823e-09 0 8.017e-09 0 8.02e-09 0.0021 8.023e-09 0 8.217e-09 0 8.22e-09 0.0021 8.223e-09 0 8.417e-09 0 8.42e-09 0.0021 8.423e-09 0 8.617e-09 0 8.62e-09 0.0021 8.623e-09 0 8.817e-09 0 8.82e-09 0.0021 8.823e-09 0 9.017e-09 0 9.02e-09 0.0021 9.023e-09 0 9.217e-09 0 9.22e-09 0.0021 9.223e-09 0 9.417e-09 0 9.42e-09 0.0021 9.423e-09 0 9.617e-09 0 9.62e-09 0.0021 9.623e-09 0 9.817e-09 0 9.82e-09 0.0021 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0021 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0021 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0021 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0021 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0021 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0021 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0021 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0021 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0021 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0021 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0021 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0021 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0021 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0021 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0021 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0021 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0021 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0021 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0021 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0021 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0021 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0021 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0021 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0021 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0021 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0021 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0021 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0021 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0021 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0021 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0021 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0021 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0021 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0021 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0021 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0021 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0021 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0021 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0021 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0021 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0021 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0021 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0021 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0021 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0021 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0021 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0021 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0021 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0021 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0021 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0021 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0021 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0021 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0021 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0021 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0021 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0021 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0021 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0021 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0021 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0021 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0021 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0021 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0021 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0021 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0021 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0021 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0021 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0021 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0021 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0021 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0021 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0021 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0021 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0021 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0021 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0021 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0021 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0021 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0021 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0021 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0021 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0021 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0021 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0021 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0021 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0021 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0021 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0021 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0021 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0021 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0021 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0021 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0021 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0021 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0021 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0021 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0021 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0021 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0021 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0021 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0021 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0021 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0021 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0021 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0021 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0021 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0021 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0021 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0021 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0021 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0021 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0021 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0021 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0021 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0021 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0021 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0021 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0021 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0021 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0021 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0021 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0021 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0021 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0021 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0021 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0021 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0021 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0021 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0021 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0021 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0021 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0021 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0021 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0021 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0021 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0021 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0021 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0021 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0021 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0021 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0021 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0021 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0021 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0021 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0021 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0021 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0021 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0021 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0021 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0021 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0021 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0021 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0021 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0021 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0021 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0021 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0021 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0021 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0021 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0021 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0021 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0021 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0021 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0021 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0021 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0021 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0021 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0021 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0021 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0021 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0021 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0021 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0021 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0021 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0021 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0021 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0021 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0021 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0021 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0021 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0021 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0021 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0021 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0021 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0021 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0021 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0021 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0021 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0021 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0021 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0021 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0021 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0021 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0021 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0021 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0021 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0021 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0021 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0021 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0021 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0021 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0021 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0021 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0021 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0021 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0021 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0021 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0021 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0021 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0021 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0021 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0021 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0021 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0021 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0021 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0021 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0021 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0021 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0021 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0021 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0021 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0021 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0021 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0021 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0021 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0021 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0021 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0021 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0021 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0021 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0021 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0021 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0021 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0021 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0021 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0021 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0021 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0021 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0021 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0021 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0021 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0021 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0021 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0021 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0021 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0021 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0021 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0021 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0021 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0021 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0021 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0021 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0021 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0021 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0021 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0021 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0021 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0021 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0021 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0021 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0021 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0021 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0021 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0021 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0021 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0021 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0021 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0021 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0021 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0021 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0021 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0021 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0021 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0021 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0021 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0021 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0021 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0021 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0021 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0021 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0021 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0021 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0021 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0021 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0021 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0021 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0021 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0021 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0021 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0021 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0021 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0021 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0021 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0021 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0021 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0021 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0021 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0021 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0021 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0021 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0021 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0021 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0021 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0021 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0021 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0021 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0021 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0021 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0021 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0021 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0021 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0021 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0021 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0021 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0021 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0021 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0021 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0021 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0021 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0021 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0021 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0021 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0021 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0021 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0021 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0021 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0021 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0021 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0021 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0021 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0021 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0021 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0021 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0021 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0021 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0021 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0021 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0021 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0021 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0021 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0021 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0021 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0021 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0021 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0021 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0021 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0021 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0021 7.9623e-08 0)
IT02|T 0 T02  PWL(0 0 1.7e-11 0 2e-11 0.0021 2.3e-11 0 2.17e-10 0 2.2e-10 0.0021 2.23e-10 0 4.17e-10 0 4.2e-10 0.0021 4.23e-10 0 6.17e-10 0 6.2e-10 0.0021 6.23e-10 0 8.17e-10 0 8.2e-10 0.0021 8.23e-10 0 1.017e-09 0 1.02e-09 0.0021 1.023e-09 0 1.217e-09 0 1.22e-09 0.0021 1.223e-09 0 1.417e-09 0 1.42e-09 0.0021 1.423e-09 0 1.617e-09 0 1.62e-09 0.0021 1.623e-09 0 1.817e-09 0 1.82e-09 0.0021 1.823e-09 0 2.017e-09 0 2.02e-09 0.0021 2.023e-09 0 2.217e-09 0 2.22e-09 0.0021 2.223e-09 0 2.417e-09 0 2.42e-09 0.0021 2.423e-09 0 2.617e-09 0 2.62e-09 0.0021 2.623e-09 0 2.817e-09 0 2.82e-09 0.0021 2.823e-09 0 3.017e-09 0 3.02e-09 0.0021 3.023e-09 0 3.217e-09 0 3.22e-09 0.0021 3.223e-09 0 3.417e-09 0 3.42e-09 0.0021 3.423e-09 0 3.617e-09 0 3.62e-09 0.0021 3.623e-09 0 3.817e-09 0 3.82e-09 0.0021 3.823e-09 0 4.017e-09 0 4.02e-09 0.0021 4.023e-09 0 4.217e-09 0 4.22e-09 0.0021 4.223e-09 0 4.417e-09 0 4.42e-09 0.0021 4.423e-09 0 4.617e-09 0 4.62e-09 0.0021 4.623e-09 0 4.817e-09 0 4.82e-09 0.0021 4.823e-09 0 5.017e-09 0 5.02e-09 0.0021 5.023e-09 0 5.217e-09 0 5.22e-09 0.0021 5.223e-09 0 5.417e-09 0 5.42e-09 0.0021 5.423e-09 0 5.617e-09 0 5.62e-09 0.0021 5.623e-09 0 5.817e-09 0 5.82e-09 0.0021 5.823e-09 0 6.017e-09 0 6.02e-09 0.0021 6.023e-09 0 6.217e-09 0 6.22e-09 0.0021 6.223e-09 0 6.417e-09 0 6.42e-09 0.0021 6.423e-09 0 6.617e-09 0 6.62e-09 0.0021 6.623e-09 0 6.817e-09 0 6.82e-09 0.0021 6.823e-09 0 7.017e-09 0 7.02e-09 0.0021 7.023e-09 0 7.217e-09 0 7.22e-09 0.0021 7.223e-09 0 7.417e-09 0 7.42e-09 0.0021 7.423e-09 0 7.617e-09 0 7.62e-09 0.0021 7.623e-09 0 7.817e-09 0 7.82e-09 0.0021 7.823e-09 0 8.017e-09 0 8.02e-09 0.0021 8.023e-09 0 8.217e-09 0 8.22e-09 0.0021 8.223e-09 0 8.417e-09 0 8.42e-09 0.0021 8.423e-09 0 8.617e-09 0 8.62e-09 0.0021 8.623e-09 0 8.817e-09 0 8.82e-09 0.0021 8.823e-09 0 9.017e-09 0 9.02e-09 0.0021 9.023e-09 0 9.217e-09 0 9.22e-09 0.0021 9.223e-09 0 9.417e-09 0 9.42e-09 0.0021 9.423e-09 0 9.617e-09 0 9.62e-09 0.0021 9.623e-09 0 9.817e-09 0 9.82e-09 0.0021 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0021 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0021 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0021 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0021 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0021 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0021 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0021 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0021 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0021 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0021 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0021 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0021 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0021 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0021 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0021 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0021 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0021 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0021 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0021 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0021 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0021 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0021 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0021 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0021 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0021 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0021 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0021 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0021 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0021 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0021 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0021 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0021 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0021 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0021 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0021 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0021 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0021 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0021 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0021 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0021 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0021 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0021 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0021 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0021 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0021 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0021 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0021 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0021 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0021 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0021 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0021 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0021 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0021 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0021 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0021 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0021 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0021 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0021 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0021 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0021 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0021 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0021 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0021 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0021 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0021 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0021 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0021 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0021 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0021 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0021 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0021 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0021 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0021 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0021 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0021 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0021 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0021 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0021 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0021 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0021 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0021 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0021 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0021 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0021 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0021 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0021 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0021 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0021 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0021 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0021 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0021 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0021 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0021 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0021 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0021 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0021 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0021 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0021 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0021 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0021 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0021 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0021 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0021 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0021 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0021 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0021 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0021 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0021 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0021 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0021 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0021 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0021 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0021 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0021 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0021 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0021 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0021 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0021 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0021 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0021 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0021 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0021 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0021 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0021 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0021 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0021 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0021 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0021 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0021 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0021 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0021 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0021 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0021 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0021 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0021 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0021 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0021 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0021 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0021 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0021 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0021 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0021 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0021 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0021 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0021 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0021 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0021 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0021 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0021 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0021 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0021 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0021 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0021 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0021 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0021 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0021 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0021 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0021 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0021 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0021 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0021 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0021 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0021 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0021 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0021 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0021 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0021 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0021 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0021 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0021 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0021 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0021 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0021 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0021 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0021 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0021 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0021 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0021 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0021 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0021 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0021 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0021 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0021 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0021 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0021 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0021 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0021 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0021 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0021 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0021 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0021 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0021 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0021 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0021 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0021 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0021 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0021 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0021 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0021 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0021 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0021 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0021 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0021 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0021 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0021 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0021 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0021 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0021 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0021 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0021 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0021 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0021 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0021 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0021 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0021 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0021 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0021 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0021 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0021 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0021 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0021 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0021 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0021 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0021 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0021 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0021 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0021 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0021 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0021 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0021 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0021 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0021 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0021 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0021 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0021 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0021 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0021 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0021 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0021 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0021 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0021 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0021 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0021 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0021 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0021 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0021 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0021 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0021 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0021 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0021 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0021 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0021 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0021 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0021 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0021 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0021 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0021 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0021 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0021 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0021 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0021 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0021 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0021 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0021 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0021 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0021 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0021 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0021 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0021 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0021 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0021 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0021 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0021 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0021 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0021 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0021 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0021 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0021 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0021 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0021 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0021 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0021 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0021 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0021 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0021 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0021 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0021 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0021 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0021 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0021 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0021 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0021 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0021 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0021 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0021 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0021 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0021 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0021 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0021 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0021 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0021 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0021 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0021 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0021 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0021 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0021 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0021 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0021 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0021 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0021 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0021 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0021 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0021 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0021 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0021 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0021 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0021 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0021 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0021 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0021 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0021 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0021 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0021 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0021 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0021 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0021 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0021 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0021 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0021 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0021 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0021 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0021 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0021 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0021 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0021 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0021 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0021 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0021 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0021 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0021 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0021 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0021 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0021 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0021 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0021 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0021 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0021 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0021 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0021 7.9623e-08 0)
IT03|T 0 T03  PWL(0 0 1.7e-11 0 2e-11 0.0021 2.3e-11 0 2.17e-10 0 2.2e-10 0.0021 2.23e-10 0 4.17e-10 0 4.2e-10 0.0021 4.23e-10 0 6.17e-10 0 6.2e-10 0.0021 6.23e-10 0 8.17e-10 0 8.2e-10 0.0021 8.23e-10 0 1.017e-09 0 1.02e-09 0.0021 1.023e-09 0 1.217e-09 0 1.22e-09 0.0021 1.223e-09 0 1.417e-09 0 1.42e-09 0.0021 1.423e-09 0 1.617e-09 0 1.62e-09 0.0021 1.623e-09 0 1.817e-09 0 1.82e-09 0.0021 1.823e-09 0 2.017e-09 0 2.02e-09 0.0021 2.023e-09 0 2.217e-09 0 2.22e-09 0.0021 2.223e-09 0 2.417e-09 0 2.42e-09 0.0021 2.423e-09 0 2.617e-09 0 2.62e-09 0.0021 2.623e-09 0 2.817e-09 0 2.82e-09 0.0021 2.823e-09 0 3.017e-09 0 3.02e-09 0.0021 3.023e-09 0 3.217e-09 0 3.22e-09 0.0021 3.223e-09 0 3.417e-09 0 3.42e-09 0.0021 3.423e-09 0 3.617e-09 0 3.62e-09 0.0021 3.623e-09 0 3.817e-09 0 3.82e-09 0.0021 3.823e-09 0 4.017e-09 0 4.02e-09 0.0021 4.023e-09 0 4.217e-09 0 4.22e-09 0.0021 4.223e-09 0 4.417e-09 0 4.42e-09 0.0021 4.423e-09 0 4.617e-09 0 4.62e-09 0.0021 4.623e-09 0 4.817e-09 0 4.82e-09 0.0021 4.823e-09 0 5.017e-09 0 5.02e-09 0.0021 5.023e-09 0 5.217e-09 0 5.22e-09 0.0021 5.223e-09 0 5.417e-09 0 5.42e-09 0.0021 5.423e-09 0 5.617e-09 0 5.62e-09 0.0021 5.623e-09 0 5.817e-09 0 5.82e-09 0.0021 5.823e-09 0 6.017e-09 0 6.02e-09 0.0021 6.023e-09 0 6.217e-09 0 6.22e-09 0.0021 6.223e-09 0 6.417e-09 0 6.42e-09 0.0021 6.423e-09 0 6.617e-09 0 6.62e-09 0.0021 6.623e-09 0 6.817e-09 0 6.82e-09 0.0021 6.823e-09 0 7.017e-09 0 7.02e-09 0.0021 7.023e-09 0 7.217e-09 0 7.22e-09 0.0021 7.223e-09 0 7.417e-09 0 7.42e-09 0.0021 7.423e-09 0 7.617e-09 0 7.62e-09 0.0021 7.623e-09 0 7.817e-09 0 7.82e-09 0.0021 7.823e-09 0 8.017e-09 0 8.02e-09 0.0021 8.023e-09 0 8.217e-09 0 8.22e-09 0.0021 8.223e-09 0 8.417e-09 0 8.42e-09 0.0021 8.423e-09 0 8.617e-09 0 8.62e-09 0.0021 8.623e-09 0 8.817e-09 0 8.82e-09 0.0021 8.823e-09 0 9.017e-09 0 9.02e-09 0.0021 9.023e-09 0 9.217e-09 0 9.22e-09 0.0021 9.223e-09 0 9.417e-09 0 9.42e-09 0.0021 9.423e-09 0 9.617e-09 0 9.62e-09 0.0021 9.623e-09 0 9.817e-09 0 9.82e-09 0.0021 9.823e-09 0 1.0017e-08 0 1.002e-08 0.0021 1.0023e-08 0 1.0217e-08 0 1.022e-08 0.0021 1.0223e-08 0 1.0417e-08 0 1.042e-08 0.0021 1.0423e-08 0 1.0617e-08 0 1.062e-08 0.0021 1.0623e-08 0 1.0817e-08 0 1.082e-08 0.0021 1.0823e-08 0 1.1017e-08 0 1.102e-08 0.0021 1.1023e-08 0 1.1217e-08 0 1.122e-08 0.0021 1.1223e-08 0 1.1417e-08 0 1.142e-08 0.0021 1.1423e-08 0 1.1617e-08 0 1.162e-08 0.0021 1.1623e-08 0 1.1817e-08 0 1.182e-08 0.0021 1.1823e-08 0 1.2017e-08 0 1.202e-08 0.0021 1.2023e-08 0 1.2217e-08 0 1.222e-08 0.0021 1.2223e-08 0 1.2417e-08 0 1.242e-08 0.0021 1.2423e-08 0 1.2617e-08 0 1.262e-08 0.0021 1.2623e-08 0 1.2817e-08 0 1.282e-08 0.0021 1.2823e-08 0 1.3017e-08 0 1.302e-08 0.0021 1.3023e-08 0 1.3217e-08 0 1.322e-08 0.0021 1.3223e-08 0 1.3417e-08 0 1.342e-08 0.0021 1.3423e-08 0 1.3617e-08 0 1.362e-08 0.0021 1.3623e-08 0 1.3817e-08 0 1.382e-08 0.0021 1.3823e-08 0 1.4017e-08 0 1.402e-08 0.0021 1.4023e-08 0 1.4217e-08 0 1.422e-08 0.0021 1.4223e-08 0 1.4417e-08 0 1.442e-08 0.0021 1.4423e-08 0 1.4617e-08 0 1.462e-08 0.0021 1.4623e-08 0 1.4817e-08 0 1.482e-08 0.0021 1.4823e-08 0 1.5017e-08 0 1.502e-08 0.0021 1.5023e-08 0 1.5217e-08 0 1.522e-08 0.0021 1.5223e-08 0 1.5417e-08 0 1.542e-08 0.0021 1.5423e-08 0 1.5617e-08 0 1.562e-08 0.0021 1.5623e-08 0 1.5817e-08 0 1.582e-08 0.0021 1.5823e-08 0 1.6017e-08 0 1.602e-08 0.0021 1.6023e-08 0 1.6217e-08 0 1.622e-08 0.0021 1.6223e-08 0 1.6417e-08 0 1.642e-08 0.0021 1.6423e-08 0 1.6617e-08 0 1.662e-08 0.0021 1.6623e-08 0 1.6817e-08 0 1.682e-08 0.0021 1.6823e-08 0 1.7017e-08 0 1.702e-08 0.0021 1.7023e-08 0 1.7217e-08 0 1.722e-08 0.0021 1.7223e-08 0 1.7417e-08 0 1.742e-08 0.0021 1.7423e-08 0 1.7617e-08 0 1.762e-08 0.0021 1.7623e-08 0 1.7817e-08 0 1.782e-08 0.0021 1.7823e-08 0 1.8017e-08 0 1.802e-08 0.0021 1.8023e-08 0 1.8217e-08 0 1.822e-08 0.0021 1.8223e-08 0 1.8417e-08 0 1.842e-08 0.0021 1.8423e-08 0 1.8617e-08 0 1.862e-08 0.0021 1.8623e-08 0 1.8817e-08 0 1.882e-08 0.0021 1.8823e-08 0 1.9017e-08 0 1.902e-08 0.0021 1.9023e-08 0 1.9217e-08 0 1.922e-08 0.0021 1.9223e-08 0 1.9417e-08 0 1.942e-08 0.0021 1.9423e-08 0 1.9617e-08 0 1.962e-08 0.0021 1.9623e-08 0 1.9817e-08 0 1.982e-08 0.0021 1.9823e-08 0 2.0017e-08 0 2.002e-08 0.0021 2.0023e-08 0 2.0217e-08 0 2.022e-08 0.0021 2.0223e-08 0 2.0417e-08 0 2.042e-08 0.0021 2.0423e-08 0 2.0617e-08 0 2.062e-08 0.0021 2.0623e-08 0 2.0817e-08 0 2.082e-08 0.0021 2.0823e-08 0 2.1017e-08 0 2.102e-08 0.0021 2.1023e-08 0 2.1217e-08 0 2.122e-08 0.0021 2.1223e-08 0 2.1417e-08 0 2.142e-08 0.0021 2.1423e-08 0 2.1617e-08 0 2.162e-08 0.0021 2.1623e-08 0 2.1817e-08 0 2.182e-08 0.0021 2.1823e-08 0 2.2017e-08 0 2.202e-08 0.0021 2.2023e-08 0 2.2217e-08 0 2.222e-08 0.0021 2.2223e-08 0 2.2417e-08 0 2.242e-08 0.0021 2.2423e-08 0 2.2617e-08 0 2.262e-08 0.0021 2.2623e-08 0 2.2817e-08 0 2.282e-08 0.0021 2.2823e-08 0 2.3017e-08 0 2.302e-08 0.0021 2.3023e-08 0 2.3217e-08 0 2.322e-08 0.0021 2.3223e-08 0 2.3417e-08 0 2.342e-08 0.0021 2.3423e-08 0 2.3617e-08 0 2.362e-08 0.0021 2.3623e-08 0 2.3817e-08 0 2.382e-08 0.0021 2.3823e-08 0 2.4017e-08 0 2.402e-08 0.0021 2.4023e-08 0 2.4217e-08 0 2.422e-08 0.0021 2.4223e-08 0 2.4417e-08 0 2.442e-08 0.0021 2.4423e-08 0 2.4617e-08 0 2.462e-08 0.0021 2.4623e-08 0 2.4817e-08 0 2.482e-08 0.0021 2.4823e-08 0 2.5017e-08 0 2.502e-08 0.0021 2.5023e-08 0 2.5217e-08 0 2.522e-08 0.0021 2.5223e-08 0 2.5417e-08 0 2.542e-08 0.0021 2.5423e-08 0 2.5617e-08 0 2.562e-08 0.0021 2.5623e-08 0 2.5817e-08 0 2.582e-08 0.0021 2.5823e-08 0 2.6017e-08 0 2.602e-08 0.0021 2.6023e-08 0 2.6217e-08 0 2.622e-08 0.0021 2.6223e-08 0 2.6417e-08 0 2.642e-08 0.0021 2.6423e-08 0 2.6617e-08 0 2.662e-08 0.0021 2.6623e-08 0 2.6817e-08 0 2.682e-08 0.0021 2.6823e-08 0 2.7017e-08 0 2.702e-08 0.0021 2.7023e-08 0 2.7217e-08 0 2.722e-08 0.0021 2.7223e-08 0 2.7417e-08 0 2.742e-08 0.0021 2.7423e-08 0 2.7617e-08 0 2.762e-08 0.0021 2.7623e-08 0 2.7817e-08 0 2.782e-08 0.0021 2.7823e-08 0 2.8017e-08 0 2.802e-08 0.0021 2.8023e-08 0 2.8217e-08 0 2.822e-08 0.0021 2.8223e-08 0 2.8417e-08 0 2.842e-08 0.0021 2.8423e-08 0 2.8617e-08 0 2.862e-08 0.0021 2.8623e-08 0 2.8817e-08 0 2.882e-08 0.0021 2.8823e-08 0 2.9017e-08 0 2.902e-08 0.0021 2.9023e-08 0 2.9217e-08 0 2.922e-08 0.0021 2.9223e-08 0 2.9417e-08 0 2.942e-08 0.0021 2.9423e-08 0 2.9617e-08 0 2.962e-08 0.0021 2.9623e-08 0 2.9817e-08 0 2.982e-08 0.0021 2.9823e-08 0 3.0017e-08 0 3.002e-08 0.0021 3.0023e-08 0 3.0217e-08 0 3.022e-08 0.0021 3.0223e-08 0 3.0417e-08 0 3.042e-08 0.0021 3.0423e-08 0 3.0617e-08 0 3.062e-08 0.0021 3.0623e-08 0 3.0817e-08 0 3.082e-08 0.0021 3.0823e-08 0 3.1017e-08 0 3.102e-08 0.0021 3.1023e-08 0 3.1217e-08 0 3.122e-08 0.0021 3.1223e-08 0 3.1417e-08 0 3.142e-08 0.0021 3.1423e-08 0 3.1617e-08 0 3.162e-08 0.0021 3.1623e-08 0 3.1817e-08 0 3.182e-08 0.0021 3.1823e-08 0 3.2017e-08 0 3.202e-08 0.0021 3.2023e-08 0 3.2217e-08 0 3.222e-08 0.0021 3.2223e-08 0 3.2417e-08 0 3.242e-08 0.0021 3.2423e-08 0 3.2617e-08 0 3.262e-08 0.0021 3.2623e-08 0 3.2817e-08 0 3.282e-08 0.0021 3.2823e-08 0 3.3017e-08 0 3.302e-08 0.0021 3.3023e-08 0 3.3217e-08 0 3.322e-08 0.0021 3.3223e-08 0 3.3417e-08 0 3.342e-08 0.0021 3.3423e-08 0 3.3617e-08 0 3.362e-08 0.0021 3.3623e-08 0 3.3817e-08 0 3.382e-08 0.0021 3.3823e-08 0 3.4017e-08 0 3.402e-08 0.0021 3.4023e-08 0 3.4217e-08 0 3.422e-08 0.0021 3.4223e-08 0 3.4417e-08 0 3.442e-08 0.0021 3.4423e-08 0 3.4617e-08 0 3.462e-08 0.0021 3.4623e-08 0 3.4817e-08 0 3.482e-08 0.0021 3.4823e-08 0 3.5017e-08 0 3.502e-08 0.0021 3.5023e-08 0 3.5217e-08 0 3.522e-08 0.0021 3.5223e-08 0 3.5417e-08 0 3.542e-08 0.0021 3.5423e-08 0 3.5617e-08 0 3.562e-08 0.0021 3.5623e-08 0 3.5817e-08 0 3.582e-08 0.0021 3.5823e-08 0 3.6017e-08 0 3.602e-08 0.0021 3.6023e-08 0 3.6217e-08 0 3.622e-08 0.0021 3.6223e-08 0 3.6417e-08 0 3.642e-08 0.0021 3.6423e-08 0 3.6617e-08 0 3.662e-08 0.0021 3.6623e-08 0 3.6817e-08 0 3.682e-08 0.0021 3.6823e-08 0 3.7017e-08 0 3.702e-08 0.0021 3.7023e-08 0 3.7217e-08 0 3.722e-08 0.0021 3.7223e-08 0 3.7417e-08 0 3.742e-08 0.0021 3.7423e-08 0 3.7617e-08 0 3.762e-08 0.0021 3.7623e-08 0 3.7817e-08 0 3.782e-08 0.0021 3.7823e-08 0 3.8017e-08 0 3.802e-08 0.0021 3.8023e-08 0 3.8217e-08 0 3.822e-08 0.0021 3.8223e-08 0 3.8417e-08 0 3.842e-08 0.0021 3.8423e-08 0 3.8617e-08 0 3.862e-08 0.0021 3.8623e-08 0 3.8817e-08 0 3.882e-08 0.0021 3.8823e-08 0 3.9017e-08 0 3.902e-08 0.0021 3.9023e-08 0 3.9217e-08 0 3.922e-08 0.0021 3.9223e-08 0 3.9417e-08 0 3.942e-08 0.0021 3.9423e-08 0 3.9617e-08 0 3.962e-08 0.0021 3.9623e-08 0 3.9817e-08 0 3.982e-08 0.0021 3.9823e-08 0 4.0017e-08 0 4.002e-08 0.0021 4.0023e-08 0 4.0217e-08 0 4.022e-08 0.0021 4.0223e-08 0 4.0417e-08 0 4.042e-08 0.0021 4.0423e-08 0 4.0617e-08 0 4.062e-08 0.0021 4.0623e-08 0 4.0817e-08 0 4.082e-08 0.0021 4.0823e-08 0 4.1017e-08 0 4.102e-08 0.0021 4.1023e-08 0 4.1217e-08 0 4.122e-08 0.0021 4.1223e-08 0 4.1417e-08 0 4.142e-08 0.0021 4.1423e-08 0 4.1617e-08 0 4.162e-08 0.0021 4.1623e-08 0 4.1817e-08 0 4.182e-08 0.0021 4.1823e-08 0 4.2017e-08 0 4.202e-08 0.0021 4.2023e-08 0 4.2217e-08 0 4.222e-08 0.0021 4.2223e-08 0 4.2417e-08 0 4.242e-08 0.0021 4.2423e-08 0 4.2617e-08 0 4.262e-08 0.0021 4.2623e-08 0 4.2817e-08 0 4.282e-08 0.0021 4.2823e-08 0 4.3017e-08 0 4.302e-08 0.0021 4.3023e-08 0 4.3217e-08 0 4.322e-08 0.0021 4.3223e-08 0 4.3417e-08 0 4.342e-08 0.0021 4.3423e-08 0 4.3617e-08 0 4.362e-08 0.0021 4.3623e-08 0 4.3817e-08 0 4.382e-08 0.0021 4.3823e-08 0 4.4017e-08 0 4.402e-08 0.0021 4.4023e-08 0 4.4217e-08 0 4.422e-08 0.0021 4.4223e-08 0 4.4417e-08 0 4.442e-08 0.0021 4.4423e-08 0 4.4617e-08 0 4.462e-08 0.0021 4.4623e-08 0 4.4817e-08 0 4.482e-08 0.0021 4.4823e-08 0 4.5017e-08 0 4.502e-08 0.0021 4.5023e-08 0 4.5217e-08 0 4.522e-08 0.0021 4.5223e-08 0 4.5417e-08 0 4.542e-08 0.0021 4.5423e-08 0 4.5617e-08 0 4.562e-08 0.0021 4.5623e-08 0 4.5817e-08 0 4.582e-08 0.0021 4.5823e-08 0 4.6017e-08 0 4.602e-08 0.0021 4.6023e-08 0 4.6217e-08 0 4.622e-08 0.0021 4.6223e-08 0 4.6417e-08 0 4.642e-08 0.0021 4.6423e-08 0 4.6617e-08 0 4.662e-08 0.0021 4.6623e-08 0 4.6817e-08 0 4.682e-08 0.0021 4.6823e-08 0 4.7017e-08 0 4.702e-08 0.0021 4.7023e-08 0 4.7217e-08 0 4.722e-08 0.0021 4.7223e-08 0 4.7417e-08 0 4.742e-08 0.0021 4.7423e-08 0 4.7617e-08 0 4.762e-08 0.0021 4.7623e-08 0 4.7817e-08 0 4.782e-08 0.0021 4.7823e-08 0 4.8017e-08 0 4.802e-08 0.0021 4.8023e-08 0 4.8217e-08 0 4.822e-08 0.0021 4.8223e-08 0 4.8417e-08 0 4.842e-08 0.0021 4.8423e-08 0 4.8617e-08 0 4.862e-08 0.0021 4.8623e-08 0 4.8817e-08 0 4.882e-08 0.0021 4.8823e-08 0 4.9017e-08 0 4.902e-08 0.0021 4.9023e-08 0 4.9217e-08 0 4.922e-08 0.0021 4.9223e-08 0 4.9417e-08 0 4.942e-08 0.0021 4.9423e-08 0 4.9617e-08 0 4.962e-08 0.0021 4.9623e-08 0 4.9817e-08 0 4.982e-08 0.0021 4.9823e-08 0 5.0017e-08 0 5.002e-08 0.0021 5.0023e-08 0 5.0217e-08 0 5.022e-08 0.0021 5.0223e-08 0 5.0417e-08 0 5.042e-08 0.0021 5.0423e-08 0 5.0617e-08 0 5.062e-08 0.0021 5.0623e-08 0 5.0817e-08 0 5.082e-08 0.0021 5.0823e-08 0 5.1017e-08 0 5.102e-08 0.0021 5.1023e-08 0 5.1217e-08 0 5.122e-08 0.0021 5.1223e-08 0 5.1417e-08 0 5.142e-08 0.0021 5.1423e-08 0 5.1617e-08 0 5.162e-08 0.0021 5.1623e-08 0 5.1817e-08 0 5.182e-08 0.0021 5.1823e-08 0 5.2017e-08 0 5.202e-08 0.0021 5.2023e-08 0 5.2217e-08 0 5.222e-08 0.0021 5.2223e-08 0 5.2417e-08 0 5.242e-08 0.0021 5.2423e-08 0 5.2617e-08 0 5.262e-08 0.0021 5.2623e-08 0 5.2817e-08 0 5.282e-08 0.0021 5.2823e-08 0 5.3017e-08 0 5.302e-08 0.0021 5.3023e-08 0 5.3217e-08 0 5.322e-08 0.0021 5.3223e-08 0 5.3417e-08 0 5.342e-08 0.0021 5.3423e-08 0 5.3617e-08 0 5.362e-08 0.0021 5.3623e-08 0 5.3817e-08 0 5.382e-08 0.0021 5.3823e-08 0 5.4017e-08 0 5.402e-08 0.0021 5.4023e-08 0 5.4217e-08 0 5.422e-08 0.0021 5.4223e-08 0 5.4417e-08 0 5.442e-08 0.0021 5.4423e-08 0 5.4617e-08 0 5.462e-08 0.0021 5.4623e-08 0 5.4817e-08 0 5.482e-08 0.0021 5.4823e-08 0 5.5017e-08 0 5.502e-08 0.0021 5.5023e-08 0 5.5217e-08 0 5.522e-08 0.0021 5.5223e-08 0 5.5417e-08 0 5.542e-08 0.0021 5.5423e-08 0 5.5617e-08 0 5.562e-08 0.0021 5.5623e-08 0 5.5817e-08 0 5.582e-08 0.0021 5.5823e-08 0 5.6017e-08 0 5.602e-08 0.0021 5.6023e-08 0 5.6217e-08 0 5.622e-08 0.0021 5.6223e-08 0 5.6417e-08 0 5.642e-08 0.0021 5.6423e-08 0 5.6617e-08 0 5.662e-08 0.0021 5.6623e-08 0 5.6817e-08 0 5.682e-08 0.0021 5.6823e-08 0 5.7017e-08 0 5.702e-08 0.0021 5.7023e-08 0 5.7217e-08 0 5.722e-08 0.0021 5.7223e-08 0 5.7417e-08 0 5.742e-08 0.0021 5.7423e-08 0 5.7617e-08 0 5.762e-08 0.0021 5.7623e-08 0 5.7817e-08 0 5.782e-08 0.0021 5.7823e-08 0 5.8017e-08 0 5.802e-08 0.0021 5.8023e-08 0 5.8217e-08 0 5.822e-08 0.0021 5.8223e-08 0 5.8417e-08 0 5.842e-08 0.0021 5.8423e-08 0 5.8617e-08 0 5.862e-08 0.0021 5.8623e-08 0 5.8817e-08 0 5.882e-08 0.0021 5.8823e-08 0 5.9017e-08 0 5.902e-08 0.0021 5.9023e-08 0 5.9217e-08 0 5.922e-08 0.0021 5.9223e-08 0 5.9417e-08 0 5.942e-08 0.0021 5.9423e-08 0 5.9617e-08 0 5.962e-08 0.0021 5.9623e-08 0 5.9817e-08 0 5.982e-08 0.0021 5.9823e-08 0 6.0017e-08 0 6.002e-08 0.0021 6.0023e-08 0 6.0217e-08 0 6.022e-08 0.0021 6.0223e-08 0 6.0417e-08 0 6.042e-08 0.0021 6.0423e-08 0 6.0617e-08 0 6.062e-08 0.0021 6.0623e-08 0 6.0817e-08 0 6.082e-08 0.0021 6.0823e-08 0 6.1017e-08 0 6.102e-08 0.0021 6.1023e-08 0 6.1217e-08 0 6.122e-08 0.0021 6.1223e-08 0 6.1417e-08 0 6.142e-08 0.0021 6.1423e-08 0 6.1617e-08 0 6.162e-08 0.0021 6.1623e-08 0 6.1817e-08 0 6.182e-08 0.0021 6.1823e-08 0 6.2017e-08 0 6.202e-08 0.0021 6.2023e-08 0 6.2217e-08 0 6.222e-08 0.0021 6.2223e-08 0 6.2417e-08 0 6.242e-08 0.0021 6.2423e-08 0 6.2617e-08 0 6.262e-08 0.0021 6.2623e-08 0 6.2817e-08 0 6.282e-08 0.0021 6.2823e-08 0 6.3017e-08 0 6.302e-08 0.0021 6.3023e-08 0 6.3217e-08 0 6.322e-08 0.0021 6.3223e-08 0 6.3417e-08 0 6.342e-08 0.0021 6.3423e-08 0 6.3617e-08 0 6.362e-08 0.0021 6.3623e-08 0 6.3817e-08 0 6.382e-08 0.0021 6.3823e-08 0 6.4017e-08 0 6.402e-08 0.0021 6.4023e-08 0 6.4217e-08 0 6.422e-08 0.0021 6.4223e-08 0 6.4417e-08 0 6.442e-08 0.0021 6.4423e-08 0 6.4617e-08 0 6.462e-08 0.0021 6.4623e-08 0 6.4817e-08 0 6.482e-08 0.0021 6.4823e-08 0 6.5017e-08 0 6.502e-08 0.0021 6.5023e-08 0 6.5217e-08 0 6.522e-08 0.0021 6.5223e-08 0 6.5417e-08 0 6.542e-08 0.0021 6.5423e-08 0 6.5617e-08 0 6.562e-08 0.0021 6.5623e-08 0 6.5817e-08 0 6.582e-08 0.0021 6.5823e-08 0 6.6017e-08 0 6.602e-08 0.0021 6.6023e-08 0 6.6217e-08 0 6.622e-08 0.0021 6.6223e-08 0 6.6417e-08 0 6.642e-08 0.0021 6.6423e-08 0 6.6617e-08 0 6.662e-08 0.0021 6.6623e-08 0 6.6817e-08 0 6.682e-08 0.0021 6.6823e-08 0 6.7017e-08 0 6.702e-08 0.0021 6.7023e-08 0 6.7217e-08 0 6.722e-08 0.0021 6.7223e-08 0 6.7417e-08 0 6.742e-08 0.0021 6.7423e-08 0 6.7617e-08 0 6.762e-08 0.0021 6.7623e-08 0 6.7817e-08 0 6.782e-08 0.0021 6.7823e-08 0 6.8017e-08 0 6.802e-08 0.0021 6.8023e-08 0 6.8217e-08 0 6.822e-08 0.0021 6.8223e-08 0 6.8417e-08 0 6.842e-08 0.0021 6.8423e-08 0 6.8617e-08 0 6.862e-08 0.0021 6.8623e-08 0 6.8817e-08 0 6.882e-08 0.0021 6.8823e-08 0 6.9017e-08 0 6.902e-08 0.0021 6.9023e-08 0 6.9217e-08 0 6.922e-08 0.0021 6.9223e-08 0 6.9417e-08 0 6.942e-08 0.0021 6.9423e-08 0 6.9617e-08 0 6.962e-08 0.0021 6.9623e-08 0 6.9817e-08 0 6.982e-08 0.0021 6.9823e-08 0 7.0017e-08 0 7.002e-08 0.0021 7.0023e-08 0 7.0217e-08 0 7.022e-08 0.0021 7.0223e-08 0 7.0417e-08 0 7.042e-08 0.0021 7.0423e-08 0 7.0617e-08 0 7.062e-08 0.0021 7.0623e-08 0 7.0817e-08 0 7.082e-08 0.0021 7.0823e-08 0 7.1017e-08 0 7.102e-08 0.0021 7.1023e-08 0 7.1217e-08 0 7.122e-08 0.0021 7.1223e-08 0 7.1417e-08 0 7.142e-08 0.0021 7.1423e-08 0 7.1617e-08 0 7.162e-08 0.0021 7.1623e-08 0 7.1817e-08 0 7.182e-08 0.0021 7.1823e-08 0 7.2017e-08 0 7.202e-08 0.0021 7.2023e-08 0 7.2217e-08 0 7.222e-08 0.0021 7.2223e-08 0 7.2417e-08 0 7.242e-08 0.0021 7.2423e-08 0 7.2617e-08 0 7.262e-08 0.0021 7.2623e-08 0 7.2817e-08 0 7.282e-08 0.0021 7.2823e-08 0 7.3017e-08 0 7.302e-08 0.0021 7.3023e-08 0 7.3217e-08 0 7.322e-08 0.0021 7.3223e-08 0 7.3417e-08 0 7.342e-08 0.0021 7.3423e-08 0 7.3617e-08 0 7.362e-08 0.0021 7.3623e-08 0 7.3817e-08 0 7.382e-08 0.0021 7.3823e-08 0 7.4017e-08 0 7.402e-08 0.0021 7.4023e-08 0 7.4217e-08 0 7.422e-08 0.0021 7.4223e-08 0 7.4417e-08 0 7.442e-08 0.0021 7.4423e-08 0 7.4617e-08 0 7.462e-08 0.0021 7.4623e-08 0 7.4817e-08 0 7.482e-08 0.0021 7.4823e-08 0 7.5017e-08 0 7.502e-08 0.0021 7.5023e-08 0 7.5217e-08 0 7.522e-08 0.0021 7.5223e-08 0 7.5417e-08 0 7.542e-08 0.0021 7.5423e-08 0 7.5617e-08 0 7.562e-08 0.0021 7.5623e-08 0 7.5817e-08 0 7.582e-08 0.0021 7.5823e-08 0 7.6017e-08 0 7.602e-08 0.0021 7.6023e-08 0 7.6217e-08 0 7.622e-08 0.0021 7.6223e-08 0 7.6417e-08 0 7.642e-08 0.0021 7.6423e-08 0 7.6617e-08 0 7.662e-08 0.0021 7.6623e-08 0 7.6817e-08 0 7.682e-08 0.0021 7.6823e-08 0 7.7017e-08 0 7.702e-08 0.0021 7.7023e-08 0 7.7217e-08 0 7.722e-08 0.0021 7.7223e-08 0 7.7417e-08 0 7.742e-08 0.0021 7.7423e-08 0 7.7617e-08 0 7.762e-08 0.0021 7.7623e-08 0 7.7817e-08 0 7.782e-08 0.0021 7.7823e-08 0 7.8017e-08 0 7.802e-08 0.0021 7.8023e-08 0 7.8217e-08 0 7.822e-08 0.0021 7.8223e-08 0 7.8417e-08 0 7.842e-08 0.0021 7.8423e-08 0 7.8617e-08 0 7.862e-08 0.0021 7.8623e-08 0 7.8817e-08 0 7.882e-08 0.0021 7.8823e-08 0 7.9017e-08 0 7.902e-08 0.0021 7.9023e-08 0 7.9217e-08 0 7.922e-08 0.0021 7.9223e-08 0 7.9417e-08 0 7.942e-08 0.0021 7.9423e-08 0 7.9617e-08 0 7.962e-08 0.0021 7.9623e-08 0)
LSPL_IG0_0|1 IG0_0 SPL_IG0_0|D1  2e-12
LSPL_IG0_0|2 SPL_IG0_0|D1 SPL_IG0_0|D2  4.135667696e-12
LSPL_IG0_0|3 SPL_IG0_0|D2 SPL_IG0_0|JCT  9.84682784761905e-13
LSPL_IG0_0|4 SPL_IG0_0|JCT SPL_IG0_0|QA1  9.84682784761905e-13
LSPL_IG0_0|5 SPL_IG0_0|QA1 IG0_0_TO0  2e-12
LSPL_IG0_0|6 SPL_IG0_0|JCT SPL_IG0_0|QB1  9.84682784761905e-13
LSPL_IG0_0|7 SPL_IG0_0|QB1 IG0_0_TO1  2e-12
LSPL_IP1_0|1 IP1_0 SPL_IP1_0|D1  2e-12
LSPL_IP1_0|2 SPL_IP1_0|D1 SPL_IP1_0|D2  4.135667696e-12
LSPL_IP1_0|3 SPL_IP1_0|D2 SPL_IP1_0|JCT  9.84682784761905e-13
LSPL_IP1_0|4 SPL_IP1_0|JCT SPL_IP1_0|QA1  9.84682784761905e-13
LSPL_IP1_0|5 SPL_IP1_0|QA1 IP1_0_TO1  2e-12
LSPL_IP1_0|6 SPL_IP1_0|JCT SPL_IP1_0|QB1  9.84682784761905e-13
LSPL_IP1_0|7 SPL_IP1_0|QB1 IP1_0_OUT  2e-12
LSPL_IG2_0|1 IG2_0 SPL_IG2_0|D1  2e-12
LSPL_IG2_0|2 SPL_IG2_0|D1 SPL_IG2_0|D2  4.135667696e-12
LSPL_IG2_0|3 SPL_IG2_0|D2 SPL_IG2_0|JCT  9.84682784761905e-13
LSPL_IG2_0|4 SPL_IG2_0|JCT SPL_IG2_0|QA1  9.84682784761905e-13
LSPL_IG2_0|5 SPL_IG2_0|QA1 IG2_0_TO2  2e-12
LSPL_IG2_0|6 SPL_IG2_0|JCT SPL_IG2_0|QB1  9.84682784761905e-13
LSPL_IG2_0|7 SPL_IG2_0|QB1 IG2_0_TO3  2e-12
LSPL_IP3_0|1 IP3_0 SPL_IP3_0|D1  2e-12
LSPL_IP3_0|2 SPL_IP3_0|D1 SPL_IP3_0|D2  4.135667696e-12
LSPL_IP3_0|3 SPL_IP3_0|D2 SPL_IP3_0|JCT  9.84682784761905e-13
LSPL_IP3_0|4 SPL_IP3_0|JCT SPL_IP3_0|QA1  9.84682784761905e-13
LSPL_IP3_0|5 SPL_IP3_0|QA1 IP3_0_TO1  2e-12
LSPL_IP3_0|6 SPL_IP3_0|JCT SPL_IP3_0|QB1  9.84682784761905e-13
LSPL_IP3_0|7 SPL_IP3_0|QB1 IP3_0_OUT  2e-12
IT04|T 0 T04  PWL(0 0 1.2e-11 0 1.5e-11 0.0014 1.8e-11 0 2.12e-10 0 2.15e-10 0.0014 2.18e-10 0 4.12e-10 0 4.15e-10 0.0014 4.18e-10 0 6.12e-10 0 6.15e-10 0.0014 6.18e-10 0 8.12e-10 0 8.15e-10 0.0014 8.18e-10 0 1.012e-09 0 1.015e-09 0.0014 1.018e-09 0 1.212e-09 0 1.215e-09 0.0014 1.218e-09 0 1.412e-09 0 1.415e-09 0.0014 1.418e-09 0 1.612e-09 0 1.615e-09 0.0014 1.618e-09 0 1.812e-09 0 1.815e-09 0.0014 1.818e-09 0 2.012e-09 0 2.015e-09 0.0014 2.018e-09 0 2.212e-09 0 2.215e-09 0.0014 2.218e-09 0 2.412e-09 0 2.415e-09 0.0014 2.418e-09 0 2.612e-09 0 2.615e-09 0.0014 2.618e-09 0 2.812e-09 0 2.815e-09 0.0014 2.818e-09 0 3.012e-09 0 3.015e-09 0.0014 3.018e-09 0 3.212e-09 0 3.215e-09 0.0014 3.218e-09 0 3.412e-09 0 3.415e-09 0.0014 3.418e-09 0 3.612e-09 0 3.615e-09 0.0014 3.618e-09 0 3.812e-09 0 3.815e-09 0.0014 3.818e-09 0 4.012e-09 0 4.015e-09 0.0014 4.018e-09 0 4.212e-09 0 4.215e-09 0.0014 4.218e-09 0 4.412e-09 0 4.415e-09 0.0014 4.418e-09 0 4.612e-09 0 4.615e-09 0.0014 4.618e-09 0 4.812e-09 0 4.815e-09 0.0014 4.818e-09 0 5.012e-09 0 5.015e-09 0.0014 5.018e-09 0 5.212e-09 0 5.215e-09 0.0014 5.218e-09 0 5.412e-09 0 5.415e-09 0.0014 5.418e-09 0 5.612e-09 0 5.615e-09 0.0014 5.618e-09 0 5.812e-09 0 5.815e-09 0.0014 5.818e-09 0 6.012e-09 0 6.015e-09 0.0014 6.018e-09 0 6.212e-09 0 6.215e-09 0.0014 6.218e-09 0 6.412e-09 0 6.415e-09 0.0014 6.418e-09 0 6.612e-09 0 6.615e-09 0.0014 6.618e-09 0 6.812e-09 0 6.815e-09 0.0014 6.818e-09 0 7.012e-09 0 7.015e-09 0.0014 7.018e-09 0 7.212e-09 0 7.215e-09 0.0014 7.218e-09 0 7.412e-09 0 7.415e-09 0.0014 7.418e-09 0 7.612e-09 0 7.615e-09 0.0014 7.618e-09 0 7.812e-09 0 7.815e-09 0.0014 7.818e-09 0 8.012e-09 0 8.015e-09 0.0014 8.018e-09 0 8.212e-09 0 8.215e-09 0.0014 8.218e-09 0 8.412e-09 0 8.415e-09 0.0014 8.418e-09 0 8.612e-09 0 8.615e-09 0.0014 8.618e-09 0 8.812e-09 0 8.815e-09 0.0014 8.818e-09 0 9.012e-09 0 9.015e-09 0.0014 9.018e-09 0 9.212e-09 0 9.215e-09 0.0014 9.218e-09 0 9.412e-09 0 9.415e-09 0.0014 9.418e-09 0 9.612e-09 0 9.615e-09 0.0014 9.618e-09 0 9.812e-09 0 9.815e-09 0.0014 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0014 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0014 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0014 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0014 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0014 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0014 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0014 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0014 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0014 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0014 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0014 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0014 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0014 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0014 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0014 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0014 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0014 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0014 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0014 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0014 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0014 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0014 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0014 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0014 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0014 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0014 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0014 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0014 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0014 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0014 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0014 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0014 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0014 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0014 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0014 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0014 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0014 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0014 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0014 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0014 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0014 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0014 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0014 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0014 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0014 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0014 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0014 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0014 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0014 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0014 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0014 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0014 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0014 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0014 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0014 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0014 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0014 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0014 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0014 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0014 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0014 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0014 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0014 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0014 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0014 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0014 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0014 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0014 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0014 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0014 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0014 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0014 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0014 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0014 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0014 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0014 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0014 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0014 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0014 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0014 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0014 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0014 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0014 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0014 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0014 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0014 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0014 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0014 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0014 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0014 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0014 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0014 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0014 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0014 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0014 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0014 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0014 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0014 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0014 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0014 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0014 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0014 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0014 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0014 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0014 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0014 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0014 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0014 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0014 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0014 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0014 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0014 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0014 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0014 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0014 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0014 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0014 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0014 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0014 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0014 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0014 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0014 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0014 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0014 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0014 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0014 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0014 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0014 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0014 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0014 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0014 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0014 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0014 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0014 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0014 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0014 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0014 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0014 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0014 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0014 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0014 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0014 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0014 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0014 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0014 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0014 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0014 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0014 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0014 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0014 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0014 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0014 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0014 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0014 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0014 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0014 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0014 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0014 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0014 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0014 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0014 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0014 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0014 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0014 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0014 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0014 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0014 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0014 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0014 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0014 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0014 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0014 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0014 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0014 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0014 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0014 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0014 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0014 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0014 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0014 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0014 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0014 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0014 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0014 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0014 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0014 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0014 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0014 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0014 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0014 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0014 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0014 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0014 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0014 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0014 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0014 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0014 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0014 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0014 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0014 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0014 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0014 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0014 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0014 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0014 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0014 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0014 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0014 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0014 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0014 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0014 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0014 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0014 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0014 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0014 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0014 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0014 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0014 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0014 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0014 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0014 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0014 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0014 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0014 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0014 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0014 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0014 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0014 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0014 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0014 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0014 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0014 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0014 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0014 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0014 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0014 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0014 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0014 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0014 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0014 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0014 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0014 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0014 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0014 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0014 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0014 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0014 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0014 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0014 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0014 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0014 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0014 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0014 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0014 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0014 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0014 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0014 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0014 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0014 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0014 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0014 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0014 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0014 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0014 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0014 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0014 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0014 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0014 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0014 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0014 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0014 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0014 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0014 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0014 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0014 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0014 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0014 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0014 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0014 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0014 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0014 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0014 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0014 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0014 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0014 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0014 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0014 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0014 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0014 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0014 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0014 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0014 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0014 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0014 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0014 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0014 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0014 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0014 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0014 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0014 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0014 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0014 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0014 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0014 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0014 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0014 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0014 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0014 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0014 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0014 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0014 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0014 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0014 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0014 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0014 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0014 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0014 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0014 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0014 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0014 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0014 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0014 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0014 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0014 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0014 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0014 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0014 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0014 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0014 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0014 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0014 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0014 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0014 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0014 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0014 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0014 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0014 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0014 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0014 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0014 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0014 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0014 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0014 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0014 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0014 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0014 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0014 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0014 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0014 7.9618e-08 0)
IT05|T 0 T05  PWL(0 0 1.2e-11 0 1.5e-11 0.0014 1.8e-11 0 2.12e-10 0 2.15e-10 0.0014 2.18e-10 0 4.12e-10 0 4.15e-10 0.0014 4.18e-10 0 6.12e-10 0 6.15e-10 0.0014 6.18e-10 0 8.12e-10 0 8.15e-10 0.0014 8.18e-10 0 1.012e-09 0 1.015e-09 0.0014 1.018e-09 0 1.212e-09 0 1.215e-09 0.0014 1.218e-09 0 1.412e-09 0 1.415e-09 0.0014 1.418e-09 0 1.612e-09 0 1.615e-09 0.0014 1.618e-09 0 1.812e-09 0 1.815e-09 0.0014 1.818e-09 0 2.012e-09 0 2.015e-09 0.0014 2.018e-09 0 2.212e-09 0 2.215e-09 0.0014 2.218e-09 0 2.412e-09 0 2.415e-09 0.0014 2.418e-09 0 2.612e-09 0 2.615e-09 0.0014 2.618e-09 0 2.812e-09 0 2.815e-09 0.0014 2.818e-09 0 3.012e-09 0 3.015e-09 0.0014 3.018e-09 0 3.212e-09 0 3.215e-09 0.0014 3.218e-09 0 3.412e-09 0 3.415e-09 0.0014 3.418e-09 0 3.612e-09 0 3.615e-09 0.0014 3.618e-09 0 3.812e-09 0 3.815e-09 0.0014 3.818e-09 0 4.012e-09 0 4.015e-09 0.0014 4.018e-09 0 4.212e-09 0 4.215e-09 0.0014 4.218e-09 0 4.412e-09 0 4.415e-09 0.0014 4.418e-09 0 4.612e-09 0 4.615e-09 0.0014 4.618e-09 0 4.812e-09 0 4.815e-09 0.0014 4.818e-09 0 5.012e-09 0 5.015e-09 0.0014 5.018e-09 0 5.212e-09 0 5.215e-09 0.0014 5.218e-09 0 5.412e-09 0 5.415e-09 0.0014 5.418e-09 0 5.612e-09 0 5.615e-09 0.0014 5.618e-09 0 5.812e-09 0 5.815e-09 0.0014 5.818e-09 0 6.012e-09 0 6.015e-09 0.0014 6.018e-09 0 6.212e-09 0 6.215e-09 0.0014 6.218e-09 0 6.412e-09 0 6.415e-09 0.0014 6.418e-09 0 6.612e-09 0 6.615e-09 0.0014 6.618e-09 0 6.812e-09 0 6.815e-09 0.0014 6.818e-09 0 7.012e-09 0 7.015e-09 0.0014 7.018e-09 0 7.212e-09 0 7.215e-09 0.0014 7.218e-09 0 7.412e-09 0 7.415e-09 0.0014 7.418e-09 0 7.612e-09 0 7.615e-09 0.0014 7.618e-09 0 7.812e-09 0 7.815e-09 0.0014 7.818e-09 0 8.012e-09 0 8.015e-09 0.0014 8.018e-09 0 8.212e-09 0 8.215e-09 0.0014 8.218e-09 0 8.412e-09 0 8.415e-09 0.0014 8.418e-09 0 8.612e-09 0 8.615e-09 0.0014 8.618e-09 0 8.812e-09 0 8.815e-09 0.0014 8.818e-09 0 9.012e-09 0 9.015e-09 0.0014 9.018e-09 0 9.212e-09 0 9.215e-09 0.0014 9.218e-09 0 9.412e-09 0 9.415e-09 0.0014 9.418e-09 0 9.612e-09 0 9.615e-09 0.0014 9.618e-09 0 9.812e-09 0 9.815e-09 0.0014 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0014 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0014 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0014 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0014 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0014 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0014 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0014 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0014 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0014 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0014 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0014 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0014 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0014 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0014 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0014 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0014 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0014 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0014 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0014 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0014 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0014 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0014 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0014 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0014 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0014 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0014 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0014 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0014 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0014 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0014 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0014 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0014 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0014 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0014 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0014 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0014 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0014 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0014 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0014 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0014 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0014 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0014 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0014 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0014 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0014 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0014 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0014 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0014 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0014 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0014 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0014 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0014 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0014 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0014 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0014 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0014 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0014 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0014 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0014 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0014 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0014 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0014 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0014 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0014 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0014 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0014 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0014 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0014 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0014 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0014 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0014 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0014 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0014 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0014 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0014 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0014 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0014 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0014 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0014 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0014 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0014 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0014 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0014 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0014 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0014 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0014 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0014 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0014 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0014 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0014 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0014 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0014 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0014 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0014 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0014 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0014 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0014 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0014 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0014 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0014 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0014 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0014 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0014 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0014 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0014 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0014 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0014 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0014 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0014 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0014 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0014 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0014 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0014 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0014 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0014 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0014 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0014 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0014 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0014 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0014 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0014 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0014 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0014 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0014 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0014 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0014 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0014 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0014 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0014 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0014 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0014 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0014 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0014 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0014 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0014 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0014 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0014 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0014 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0014 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0014 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0014 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0014 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0014 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0014 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0014 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0014 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0014 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0014 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0014 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0014 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0014 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0014 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0014 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0014 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0014 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0014 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0014 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0014 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0014 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0014 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0014 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0014 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0014 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0014 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0014 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0014 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0014 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0014 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0014 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0014 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0014 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0014 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0014 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0014 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0014 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0014 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0014 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0014 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0014 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0014 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0014 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0014 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0014 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0014 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0014 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0014 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0014 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0014 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0014 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0014 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0014 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0014 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0014 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0014 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0014 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0014 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0014 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0014 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0014 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0014 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0014 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0014 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0014 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0014 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0014 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0014 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0014 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0014 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0014 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0014 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0014 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0014 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0014 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0014 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0014 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0014 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0014 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0014 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0014 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0014 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0014 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0014 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0014 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0014 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0014 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0014 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0014 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0014 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0014 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0014 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0014 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0014 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0014 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0014 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0014 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0014 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0014 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0014 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0014 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0014 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0014 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0014 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0014 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0014 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0014 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0014 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0014 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0014 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0014 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0014 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0014 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0014 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0014 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0014 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0014 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0014 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0014 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0014 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0014 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0014 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0014 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0014 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0014 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0014 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0014 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0014 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0014 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0014 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0014 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0014 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0014 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0014 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0014 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0014 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0014 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0014 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0014 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0014 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0014 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0014 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0014 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0014 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0014 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0014 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0014 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0014 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0014 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0014 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0014 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0014 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0014 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0014 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0014 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0014 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0014 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0014 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0014 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0014 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0014 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0014 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0014 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0014 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0014 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0014 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0014 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0014 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0014 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0014 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0014 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0014 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0014 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0014 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0014 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0014 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0014 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0014 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0014 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0014 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0014 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0014 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0014 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0014 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0014 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0014 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0014 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0014 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0014 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0014 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0014 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0014 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0014 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0014 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0014 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0014 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0014 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0014 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0014 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0014 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0014 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0014 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0014 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0014 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0014 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0014 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0014 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0014 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0014 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0014 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0014 7.9618e-08 0)
IT06|T 0 T06  PWL(0 0 1.2e-11 0 1.5e-11 0.0014 1.8e-11 0 2.12e-10 0 2.15e-10 0.0014 2.18e-10 0 4.12e-10 0 4.15e-10 0.0014 4.18e-10 0 6.12e-10 0 6.15e-10 0.0014 6.18e-10 0 8.12e-10 0 8.15e-10 0.0014 8.18e-10 0 1.012e-09 0 1.015e-09 0.0014 1.018e-09 0 1.212e-09 0 1.215e-09 0.0014 1.218e-09 0 1.412e-09 0 1.415e-09 0.0014 1.418e-09 0 1.612e-09 0 1.615e-09 0.0014 1.618e-09 0 1.812e-09 0 1.815e-09 0.0014 1.818e-09 0 2.012e-09 0 2.015e-09 0.0014 2.018e-09 0 2.212e-09 0 2.215e-09 0.0014 2.218e-09 0 2.412e-09 0 2.415e-09 0.0014 2.418e-09 0 2.612e-09 0 2.615e-09 0.0014 2.618e-09 0 2.812e-09 0 2.815e-09 0.0014 2.818e-09 0 3.012e-09 0 3.015e-09 0.0014 3.018e-09 0 3.212e-09 0 3.215e-09 0.0014 3.218e-09 0 3.412e-09 0 3.415e-09 0.0014 3.418e-09 0 3.612e-09 0 3.615e-09 0.0014 3.618e-09 0 3.812e-09 0 3.815e-09 0.0014 3.818e-09 0 4.012e-09 0 4.015e-09 0.0014 4.018e-09 0 4.212e-09 0 4.215e-09 0.0014 4.218e-09 0 4.412e-09 0 4.415e-09 0.0014 4.418e-09 0 4.612e-09 0 4.615e-09 0.0014 4.618e-09 0 4.812e-09 0 4.815e-09 0.0014 4.818e-09 0 5.012e-09 0 5.015e-09 0.0014 5.018e-09 0 5.212e-09 0 5.215e-09 0.0014 5.218e-09 0 5.412e-09 0 5.415e-09 0.0014 5.418e-09 0 5.612e-09 0 5.615e-09 0.0014 5.618e-09 0 5.812e-09 0 5.815e-09 0.0014 5.818e-09 0 6.012e-09 0 6.015e-09 0.0014 6.018e-09 0 6.212e-09 0 6.215e-09 0.0014 6.218e-09 0 6.412e-09 0 6.415e-09 0.0014 6.418e-09 0 6.612e-09 0 6.615e-09 0.0014 6.618e-09 0 6.812e-09 0 6.815e-09 0.0014 6.818e-09 0 7.012e-09 0 7.015e-09 0.0014 7.018e-09 0 7.212e-09 0 7.215e-09 0.0014 7.218e-09 0 7.412e-09 0 7.415e-09 0.0014 7.418e-09 0 7.612e-09 0 7.615e-09 0.0014 7.618e-09 0 7.812e-09 0 7.815e-09 0.0014 7.818e-09 0 8.012e-09 0 8.015e-09 0.0014 8.018e-09 0 8.212e-09 0 8.215e-09 0.0014 8.218e-09 0 8.412e-09 0 8.415e-09 0.0014 8.418e-09 0 8.612e-09 0 8.615e-09 0.0014 8.618e-09 0 8.812e-09 0 8.815e-09 0.0014 8.818e-09 0 9.012e-09 0 9.015e-09 0.0014 9.018e-09 0 9.212e-09 0 9.215e-09 0.0014 9.218e-09 0 9.412e-09 0 9.415e-09 0.0014 9.418e-09 0 9.612e-09 0 9.615e-09 0.0014 9.618e-09 0 9.812e-09 0 9.815e-09 0.0014 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0014 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0014 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0014 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0014 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0014 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0014 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0014 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0014 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0014 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0014 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0014 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0014 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0014 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0014 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0014 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0014 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0014 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0014 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0014 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0014 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0014 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0014 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0014 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0014 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0014 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0014 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0014 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0014 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0014 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0014 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0014 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0014 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0014 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0014 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0014 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0014 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0014 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0014 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0014 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0014 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0014 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0014 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0014 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0014 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0014 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0014 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0014 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0014 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0014 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0014 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0014 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0014 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0014 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0014 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0014 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0014 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0014 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0014 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0014 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0014 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0014 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0014 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0014 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0014 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0014 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0014 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0014 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0014 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0014 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0014 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0014 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0014 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0014 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0014 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0014 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0014 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0014 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0014 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0014 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0014 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0014 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0014 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0014 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0014 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0014 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0014 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0014 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0014 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0014 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0014 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0014 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0014 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0014 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0014 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0014 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0014 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0014 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0014 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0014 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0014 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0014 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0014 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0014 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0014 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0014 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0014 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0014 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0014 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0014 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0014 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0014 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0014 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0014 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0014 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0014 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0014 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0014 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0014 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0014 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0014 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0014 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0014 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0014 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0014 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0014 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0014 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0014 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0014 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0014 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0014 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0014 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0014 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0014 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0014 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0014 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0014 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0014 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0014 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0014 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0014 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0014 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0014 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0014 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0014 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0014 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0014 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0014 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0014 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0014 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0014 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0014 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0014 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0014 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0014 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0014 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0014 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0014 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0014 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0014 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0014 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0014 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0014 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0014 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0014 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0014 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0014 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0014 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0014 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0014 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0014 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0014 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0014 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0014 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0014 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0014 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0014 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0014 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0014 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0014 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0014 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0014 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0014 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0014 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0014 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0014 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0014 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0014 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0014 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0014 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0014 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0014 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0014 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0014 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0014 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0014 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0014 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0014 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0014 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0014 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0014 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0014 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0014 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0014 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0014 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0014 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0014 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0014 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0014 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0014 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0014 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0014 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0014 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0014 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0014 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0014 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0014 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0014 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0014 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0014 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0014 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0014 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0014 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0014 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0014 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0014 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0014 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0014 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0014 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0014 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0014 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0014 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0014 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0014 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0014 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0014 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0014 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0014 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0014 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0014 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0014 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0014 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0014 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0014 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0014 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0014 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0014 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0014 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0014 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0014 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0014 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0014 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0014 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0014 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0014 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0014 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0014 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0014 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0014 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0014 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0014 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0014 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0014 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0014 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0014 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0014 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0014 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0014 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0014 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0014 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0014 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0014 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0014 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0014 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0014 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0014 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0014 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0014 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0014 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0014 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0014 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0014 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0014 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0014 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0014 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0014 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0014 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0014 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0014 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0014 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0014 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0014 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0014 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0014 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0014 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0014 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0014 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0014 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0014 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0014 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0014 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0014 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0014 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0014 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0014 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0014 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0014 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0014 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0014 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0014 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0014 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0014 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0014 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0014 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0014 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0014 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0014 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0014 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0014 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0014 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0014 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0014 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0014 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0014 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0014 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0014 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0014 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0014 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0014 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0014 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0014 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0014 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0014 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0014 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0014 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0014 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0014 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0014 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0014 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0014 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0014 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0014 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0014 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0014 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0014 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0014 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0014 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0014 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0014 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0014 7.9618e-08 0)
IT07|T 0 T07  PWL(0 0 1.2e-11 0 1.5e-11 0.0028 1.8e-11 0 2.12e-10 0 2.15e-10 0.0028 2.18e-10 0 4.12e-10 0 4.15e-10 0.0028 4.18e-10 0 6.12e-10 0 6.15e-10 0.0028 6.18e-10 0 8.12e-10 0 8.15e-10 0.0028 8.18e-10 0 1.012e-09 0 1.015e-09 0.0028 1.018e-09 0 1.212e-09 0 1.215e-09 0.0028 1.218e-09 0 1.412e-09 0 1.415e-09 0.0028 1.418e-09 0 1.612e-09 0 1.615e-09 0.0028 1.618e-09 0 1.812e-09 0 1.815e-09 0.0028 1.818e-09 0 2.012e-09 0 2.015e-09 0.0028 2.018e-09 0 2.212e-09 0 2.215e-09 0.0028 2.218e-09 0 2.412e-09 0 2.415e-09 0.0028 2.418e-09 0 2.612e-09 0 2.615e-09 0.0028 2.618e-09 0 2.812e-09 0 2.815e-09 0.0028 2.818e-09 0 3.012e-09 0 3.015e-09 0.0028 3.018e-09 0 3.212e-09 0 3.215e-09 0.0028 3.218e-09 0 3.412e-09 0 3.415e-09 0.0028 3.418e-09 0 3.612e-09 0 3.615e-09 0.0028 3.618e-09 0 3.812e-09 0 3.815e-09 0.0028 3.818e-09 0 4.012e-09 0 4.015e-09 0.0028 4.018e-09 0 4.212e-09 0 4.215e-09 0.0028 4.218e-09 0 4.412e-09 0 4.415e-09 0.0028 4.418e-09 0 4.612e-09 0 4.615e-09 0.0028 4.618e-09 0 4.812e-09 0 4.815e-09 0.0028 4.818e-09 0 5.012e-09 0 5.015e-09 0.0028 5.018e-09 0 5.212e-09 0 5.215e-09 0.0028 5.218e-09 0 5.412e-09 0 5.415e-09 0.0028 5.418e-09 0 5.612e-09 0 5.615e-09 0.0028 5.618e-09 0 5.812e-09 0 5.815e-09 0.0028 5.818e-09 0 6.012e-09 0 6.015e-09 0.0028 6.018e-09 0 6.212e-09 0 6.215e-09 0.0028 6.218e-09 0 6.412e-09 0 6.415e-09 0.0028 6.418e-09 0 6.612e-09 0 6.615e-09 0.0028 6.618e-09 0 6.812e-09 0 6.815e-09 0.0028 6.818e-09 0 7.012e-09 0 7.015e-09 0.0028 7.018e-09 0 7.212e-09 0 7.215e-09 0.0028 7.218e-09 0 7.412e-09 0 7.415e-09 0.0028 7.418e-09 0 7.612e-09 0 7.615e-09 0.0028 7.618e-09 0 7.812e-09 0 7.815e-09 0.0028 7.818e-09 0 8.012e-09 0 8.015e-09 0.0028 8.018e-09 0 8.212e-09 0 8.215e-09 0.0028 8.218e-09 0 8.412e-09 0 8.415e-09 0.0028 8.418e-09 0 8.612e-09 0 8.615e-09 0.0028 8.618e-09 0 8.812e-09 0 8.815e-09 0.0028 8.818e-09 0 9.012e-09 0 9.015e-09 0.0028 9.018e-09 0 9.212e-09 0 9.215e-09 0.0028 9.218e-09 0 9.412e-09 0 9.415e-09 0.0028 9.418e-09 0 9.612e-09 0 9.615e-09 0.0028 9.618e-09 0 9.812e-09 0 9.815e-09 0.0028 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0028 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0028 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0028 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0028 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0028 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0028 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0028 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0028 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0028 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0028 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0028 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0028 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0028 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0028 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0028 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0028 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0028 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0028 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0028 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0028 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0028 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0028 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0028 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0028 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0028 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0028 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0028 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0028 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0028 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0028 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0028 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0028 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0028 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0028 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0028 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0028 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0028 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0028 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0028 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0028 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0028 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0028 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0028 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0028 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0028 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0028 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0028 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0028 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0028 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0028 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0028 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0028 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0028 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0028 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0028 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0028 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0028 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0028 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0028 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0028 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0028 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0028 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0028 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0028 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0028 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0028 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0028 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0028 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0028 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0028 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0028 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0028 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0028 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0028 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0028 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0028 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0028 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0028 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0028 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0028 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0028 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0028 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0028 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0028 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0028 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0028 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0028 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0028 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0028 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0028 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0028 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0028 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0028 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0028 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0028 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0028 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0028 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0028 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0028 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0028 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0028 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0028 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0028 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0028 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0028 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0028 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0028 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0028 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0028 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0028 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0028 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0028 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0028 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0028 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0028 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0028 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0028 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0028 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0028 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0028 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0028 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0028 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0028 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0028 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0028 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0028 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0028 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0028 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0028 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0028 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0028 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0028 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0028 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0028 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0028 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0028 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0028 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0028 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0028 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0028 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0028 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0028 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0028 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0028 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0028 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0028 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0028 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0028 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0028 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0028 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0028 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0028 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0028 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0028 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0028 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0028 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0028 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0028 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0028 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0028 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0028 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0028 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0028 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0028 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0028 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0028 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0028 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0028 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0028 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0028 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0028 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0028 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0028 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0028 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0028 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0028 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0028 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0028 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0028 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0028 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0028 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0028 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0028 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0028 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0028 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0028 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0028 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0028 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0028 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0028 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0028 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0028 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0028 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0028 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0028 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0028 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0028 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0028 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0028 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0028 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0028 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0028 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0028 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0028 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0028 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0028 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0028 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0028 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0028 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0028 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0028 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0028 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0028 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0028 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0028 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0028 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0028 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0028 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0028 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0028 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0028 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0028 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0028 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0028 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0028 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0028 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0028 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0028 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0028 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0028 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0028 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0028 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0028 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0028 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0028 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0028 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0028 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0028 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0028 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0028 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0028 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0028 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0028 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0028 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0028 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0028 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0028 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0028 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0028 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0028 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0028 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0028 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0028 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0028 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0028 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0028 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0028 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0028 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0028 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0028 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0028 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0028 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0028 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0028 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0028 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0028 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0028 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0028 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0028 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0028 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0028 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0028 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0028 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0028 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0028 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0028 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0028 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0028 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0028 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0028 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0028 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0028 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0028 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0028 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0028 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0028 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0028 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0028 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0028 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0028 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0028 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0028 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0028 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0028 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0028 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0028 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0028 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0028 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0028 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0028 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0028 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0028 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0028 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0028 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0028 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0028 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0028 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0028 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0028 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0028 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0028 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0028 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0028 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0028 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0028 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0028 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0028 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0028 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0028 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0028 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0028 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0028 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0028 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0028 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0028 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0028 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0028 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0028 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0028 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0028 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0028 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0028 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0028 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0028 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0028 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0028 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0028 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0028 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0028 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0028 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0028 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0028 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0028 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0028 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0028 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0028 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0028 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0028 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0028 7.9618e-08 0)
ID01|T 0 D01  PWL(0 0 1.2e-11 0 1.5e-11 0.0007 1.8e-11 0 2.12e-10 0 2.15e-10 0.0007 2.18e-10 0 4.12e-10 0 4.15e-10 0.0007 4.18e-10 0 6.12e-10 0 6.15e-10 0.0007 6.18e-10 0 8.12e-10 0 8.15e-10 0.0007 8.18e-10 0 1.012e-09 0 1.015e-09 0.0007 1.018e-09 0 1.212e-09 0 1.215e-09 0.0007 1.218e-09 0 1.412e-09 0 1.415e-09 0.0007 1.418e-09 0 1.612e-09 0 1.615e-09 0.0007 1.618e-09 0 1.812e-09 0 1.815e-09 0.0007 1.818e-09 0 2.012e-09 0 2.015e-09 0.0007 2.018e-09 0 2.212e-09 0 2.215e-09 0.0007 2.218e-09 0 2.412e-09 0 2.415e-09 0.0007 2.418e-09 0 2.612e-09 0 2.615e-09 0.0007 2.618e-09 0 2.812e-09 0 2.815e-09 0.0007 2.818e-09 0 3.012e-09 0 3.015e-09 0.0007 3.018e-09 0 3.212e-09 0 3.215e-09 0.0007 3.218e-09 0 3.412e-09 0 3.415e-09 0.0007 3.418e-09 0 3.612e-09 0 3.615e-09 0.0007 3.618e-09 0 3.812e-09 0 3.815e-09 0.0007 3.818e-09 0 4.012e-09 0 4.015e-09 0.0007 4.018e-09 0 4.212e-09 0 4.215e-09 0.0007 4.218e-09 0 4.412e-09 0 4.415e-09 0.0007 4.418e-09 0 4.612e-09 0 4.615e-09 0.0007 4.618e-09 0 4.812e-09 0 4.815e-09 0.0007 4.818e-09 0 5.012e-09 0 5.015e-09 0.0007 5.018e-09 0 5.212e-09 0 5.215e-09 0.0007 5.218e-09 0 5.412e-09 0 5.415e-09 0.0007 5.418e-09 0 5.612e-09 0 5.615e-09 0.0007 5.618e-09 0 5.812e-09 0 5.815e-09 0.0007 5.818e-09 0 6.012e-09 0 6.015e-09 0.0007 6.018e-09 0 6.212e-09 0 6.215e-09 0.0007 6.218e-09 0 6.412e-09 0 6.415e-09 0.0007 6.418e-09 0 6.612e-09 0 6.615e-09 0.0007 6.618e-09 0 6.812e-09 0 6.815e-09 0.0007 6.818e-09 0 7.012e-09 0 7.015e-09 0.0007 7.018e-09 0 7.212e-09 0 7.215e-09 0.0007 7.218e-09 0 7.412e-09 0 7.415e-09 0.0007 7.418e-09 0 7.612e-09 0 7.615e-09 0.0007 7.618e-09 0 7.812e-09 0 7.815e-09 0.0007 7.818e-09 0 8.012e-09 0 8.015e-09 0.0007 8.018e-09 0 8.212e-09 0 8.215e-09 0.0007 8.218e-09 0 8.412e-09 0 8.415e-09 0.0007 8.418e-09 0 8.612e-09 0 8.615e-09 0.0007 8.618e-09 0 8.812e-09 0 8.815e-09 0.0007 8.818e-09 0 9.012e-09 0 9.015e-09 0.0007 9.018e-09 0 9.212e-09 0 9.215e-09 0.0007 9.218e-09 0 9.412e-09 0 9.415e-09 0.0007 9.418e-09 0 9.612e-09 0 9.615e-09 0.0007 9.618e-09 0 9.812e-09 0 9.815e-09 0.0007 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0007 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0007 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0007 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0007 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0007 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0007 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0007 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0007 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0007 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0007 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0007 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0007 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0007 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0007 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0007 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0007 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0007 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0007 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0007 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0007 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0007 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0007 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0007 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0007 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0007 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0007 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0007 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0007 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0007 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0007 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0007 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0007 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0007 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0007 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0007 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0007 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0007 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0007 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0007 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0007 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0007 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0007 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0007 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0007 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0007 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0007 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0007 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0007 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0007 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0007 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0007 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0007 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0007 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0007 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0007 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0007 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0007 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0007 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0007 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0007 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0007 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0007 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0007 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0007 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0007 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0007 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0007 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0007 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0007 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0007 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0007 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0007 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0007 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0007 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0007 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0007 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0007 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0007 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0007 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0007 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0007 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0007 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0007 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0007 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0007 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0007 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0007 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0007 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0007 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0007 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0007 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0007 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0007 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0007 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0007 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0007 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0007 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0007 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0007 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0007 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0007 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0007 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0007 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0007 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0007 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0007 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0007 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0007 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0007 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0007 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0007 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0007 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0007 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0007 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0007 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0007 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0007 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0007 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0007 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0007 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0007 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0007 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0007 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0007 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0007 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0007 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0007 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0007 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0007 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0007 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0007 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0007 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0007 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0007 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0007 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0007 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0007 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0007 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0007 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0007 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0007 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0007 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0007 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0007 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0007 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0007 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0007 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0007 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0007 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0007 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0007 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0007 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0007 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0007 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0007 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0007 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0007 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0007 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0007 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0007 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0007 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0007 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0007 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0007 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0007 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0007 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0007 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0007 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0007 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0007 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0007 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0007 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0007 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0007 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0007 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0007 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0007 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0007 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0007 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0007 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0007 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0007 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0007 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0007 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0007 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0007 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0007 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0007 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0007 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0007 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0007 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0007 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0007 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0007 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0007 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0007 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0007 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0007 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0007 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0007 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0007 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0007 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0007 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0007 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0007 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0007 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0007 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0007 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0007 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0007 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0007 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0007 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0007 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0007 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0007 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0007 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0007 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0007 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0007 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0007 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0007 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0007 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0007 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0007 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0007 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0007 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0007 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0007 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0007 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0007 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0007 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0007 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0007 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0007 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0007 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0007 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0007 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0007 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0007 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0007 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0007 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0007 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0007 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0007 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0007 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0007 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0007 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0007 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0007 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0007 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0007 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0007 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0007 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0007 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0007 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0007 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0007 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0007 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0007 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0007 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0007 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0007 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0007 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0007 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0007 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0007 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0007 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0007 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0007 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0007 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0007 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0007 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0007 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0007 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0007 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0007 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0007 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0007 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0007 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0007 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0007 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0007 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0007 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0007 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0007 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0007 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0007 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0007 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0007 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0007 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0007 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0007 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0007 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0007 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0007 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0007 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0007 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0007 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0007 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0007 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0007 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0007 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0007 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0007 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0007 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0007 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0007 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0007 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0007 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0007 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0007 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0007 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0007 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0007 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0007 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0007 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0007 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0007 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0007 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0007 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0007 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0007 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0007 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0007 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0007 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0007 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0007 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0007 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0007 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0007 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0007 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0007 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0007 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0007 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0007 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0007 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0007 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0007 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0007 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0007 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0007 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0007 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0007 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0007 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0007 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0007 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0007 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0007 7.9618e-08 0)
L_DFF_IP1_01|1 IP1_0_OUT _DFF_IP1_01|A1  2.067833848e-12
L_DFF_IP1_01|2 _DFF_IP1_01|A1 _DFF_IP1_01|A2  4.135667696e-12
L_DFF_IP1_01|3 _DFF_IP1_01|A3 _DFF_IP1_01|A4  8.271335392e-12
L_DFF_IP1_01|T D01 _DFF_IP1_01|T1  2.067833848e-12
L_DFF_IP1_01|4 _DFF_IP1_01|T1 _DFF_IP1_01|T2  4.135667696e-12
L_DFF_IP1_01|5 _DFF_IP1_01|A4 _DFF_IP1_01|Q1  4.135667696e-12
L_DFF_IP1_01|6 _DFF_IP1_01|Q1 IP1_1_OUT  2.067833848e-12
ID02|T 0 D02  PWL(0 0 1.2e-11 0 1.5e-11 0.0007 1.8e-11 0 2.12e-10 0 2.15e-10 0.0007 2.18e-10 0 4.12e-10 0 4.15e-10 0.0007 4.18e-10 0 6.12e-10 0 6.15e-10 0.0007 6.18e-10 0 8.12e-10 0 8.15e-10 0.0007 8.18e-10 0 1.012e-09 0 1.015e-09 0.0007 1.018e-09 0 1.212e-09 0 1.215e-09 0.0007 1.218e-09 0 1.412e-09 0 1.415e-09 0.0007 1.418e-09 0 1.612e-09 0 1.615e-09 0.0007 1.618e-09 0 1.812e-09 0 1.815e-09 0.0007 1.818e-09 0 2.012e-09 0 2.015e-09 0.0007 2.018e-09 0 2.212e-09 0 2.215e-09 0.0007 2.218e-09 0 2.412e-09 0 2.415e-09 0.0007 2.418e-09 0 2.612e-09 0 2.615e-09 0.0007 2.618e-09 0 2.812e-09 0 2.815e-09 0.0007 2.818e-09 0 3.012e-09 0 3.015e-09 0.0007 3.018e-09 0 3.212e-09 0 3.215e-09 0.0007 3.218e-09 0 3.412e-09 0 3.415e-09 0.0007 3.418e-09 0 3.612e-09 0 3.615e-09 0.0007 3.618e-09 0 3.812e-09 0 3.815e-09 0.0007 3.818e-09 0 4.012e-09 0 4.015e-09 0.0007 4.018e-09 0 4.212e-09 0 4.215e-09 0.0007 4.218e-09 0 4.412e-09 0 4.415e-09 0.0007 4.418e-09 0 4.612e-09 0 4.615e-09 0.0007 4.618e-09 0 4.812e-09 0 4.815e-09 0.0007 4.818e-09 0 5.012e-09 0 5.015e-09 0.0007 5.018e-09 0 5.212e-09 0 5.215e-09 0.0007 5.218e-09 0 5.412e-09 0 5.415e-09 0.0007 5.418e-09 0 5.612e-09 0 5.615e-09 0.0007 5.618e-09 0 5.812e-09 0 5.815e-09 0.0007 5.818e-09 0 6.012e-09 0 6.015e-09 0.0007 6.018e-09 0 6.212e-09 0 6.215e-09 0.0007 6.218e-09 0 6.412e-09 0 6.415e-09 0.0007 6.418e-09 0 6.612e-09 0 6.615e-09 0.0007 6.618e-09 0 6.812e-09 0 6.815e-09 0.0007 6.818e-09 0 7.012e-09 0 7.015e-09 0.0007 7.018e-09 0 7.212e-09 0 7.215e-09 0.0007 7.218e-09 0 7.412e-09 0 7.415e-09 0.0007 7.418e-09 0 7.612e-09 0 7.615e-09 0.0007 7.618e-09 0 7.812e-09 0 7.815e-09 0.0007 7.818e-09 0 8.012e-09 0 8.015e-09 0.0007 8.018e-09 0 8.212e-09 0 8.215e-09 0.0007 8.218e-09 0 8.412e-09 0 8.415e-09 0.0007 8.418e-09 0 8.612e-09 0 8.615e-09 0.0007 8.618e-09 0 8.812e-09 0 8.815e-09 0.0007 8.818e-09 0 9.012e-09 0 9.015e-09 0.0007 9.018e-09 0 9.212e-09 0 9.215e-09 0.0007 9.218e-09 0 9.412e-09 0 9.415e-09 0.0007 9.418e-09 0 9.612e-09 0 9.615e-09 0.0007 9.618e-09 0 9.812e-09 0 9.815e-09 0.0007 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0007 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0007 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0007 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0007 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0007 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0007 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0007 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0007 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0007 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0007 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0007 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0007 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0007 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0007 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0007 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0007 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0007 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0007 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0007 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0007 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0007 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0007 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0007 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0007 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0007 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0007 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0007 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0007 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0007 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0007 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0007 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0007 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0007 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0007 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0007 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0007 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0007 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0007 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0007 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0007 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0007 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0007 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0007 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0007 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0007 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0007 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0007 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0007 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0007 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0007 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0007 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0007 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0007 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0007 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0007 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0007 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0007 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0007 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0007 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0007 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0007 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0007 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0007 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0007 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0007 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0007 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0007 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0007 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0007 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0007 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0007 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0007 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0007 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0007 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0007 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0007 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0007 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0007 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0007 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0007 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0007 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0007 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0007 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0007 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0007 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0007 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0007 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0007 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0007 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0007 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0007 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0007 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0007 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0007 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0007 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0007 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0007 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0007 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0007 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0007 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0007 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0007 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0007 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0007 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0007 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0007 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0007 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0007 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0007 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0007 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0007 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0007 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0007 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0007 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0007 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0007 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0007 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0007 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0007 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0007 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0007 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0007 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0007 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0007 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0007 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0007 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0007 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0007 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0007 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0007 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0007 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0007 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0007 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0007 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0007 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0007 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0007 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0007 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0007 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0007 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0007 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0007 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0007 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0007 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0007 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0007 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0007 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0007 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0007 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0007 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0007 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0007 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0007 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0007 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0007 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0007 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0007 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0007 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0007 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0007 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0007 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0007 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0007 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0007 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0007 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0007 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0007 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0007 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0007 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0007 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0007 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0007 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0007 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0007 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0007 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0007 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0007 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0007 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0007 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0007 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0007 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0007 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0007 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0007 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0007 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0007 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0007 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0007 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0007 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0007 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0007 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0007 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0007 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0007 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0007 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0007 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0007 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0007 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0007 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0007 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0007 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0007 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0007 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0007 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0007 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0007 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0007 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0007 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0007 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0007 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0007 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0007 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0007 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0007 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0007 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0007 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0007 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0007 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0007 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0007 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0007 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0007 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0007 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0007 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0007 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0007 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0007 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0007 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0007 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0007 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0007 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0007 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0007 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0007 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0007 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0007 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0007 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0007 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0007 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0007 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0007 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0007 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0007 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0007 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0007 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0007 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0007 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0007 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0007 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0007 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0007 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0007 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0007 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0007 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0007 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0007 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0007 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0007 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0007 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0007 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0007 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0007 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0007 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0007 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0007 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0007 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0007 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0007 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0007 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0007 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0007 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0007 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0007 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0007 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0007 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0007 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0007 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0007 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0007 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0007 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0007 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0007 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0007 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0007 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0007 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0007 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0007 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0007 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0007 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0007 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0007 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0007 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0007 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0007 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0007 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0007 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0007 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0007 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0007 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0007 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0007 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0007 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0007 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0007 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0007 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0007 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0007 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0007 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0007 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0007 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0007 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0007 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0007 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0007 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0007 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0007 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0007 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0007 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0007 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0007 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0007 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0007 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0007 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0007 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0007 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0007 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0007 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0007 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0007 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0007 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0007 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0007 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0007 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0007 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0007 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0007 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0007 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0007 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0007 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0007 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0007 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0007 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0007 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0007 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0007 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0007 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0007 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0007 7.9618e-08 0)
L_DFF_IP2_01|1 IP2_0_OUT _DFF_IP2_01|A1  2.067833848e-12
L_DFF_IP2_01|2 _DFF_IP2_01|A1 _DFF_IP2_01|A2  4.135667696e-12
L_DFF_IP2_01|3 _DFF_IP2_01|A3 _DFF_IP2_01|A4  8.271335392e-12
L_DFF_IP2_01|T D02 _DFF_IP2_01|T1  2.067833848e-12
L_DFF_IP2_01|4 _DFF_IP2_01|T1 _DFF_IP2_01|T2  4.135667696e-12
L_DFF_IP2_01|5 _DFF_IP2_01|A4 _DFF_IP2_01|Q1  4.135667696e-12
L_DFF_IP2_01|6 _DFF_IP2_01|Q1 IP2_1_OUT  2.067833848e-12
ID03|T 0 D03  PWL(0 0 1.2e-11 0 1.5e-11 0.0007 1.8e-11 0 2.12e-10 0 2.15e-10 0.0007 2.18e-10 0 4.12e-10 0 4.15e-10 0.0007 4.18e-10 0 6.12e-10 0 6.15e-10 0.0007 6.18e-10 0 8.12e-10 0 8.15e-10 0.0007 8.18e-10 0 1.012e-09 0 1.015e-09 0.0007 1.018e-09 0 1.212e-09 0 1.215e-09 0.0007 1.218e-09 0 1.412e-09 0 1.415e-09 0.0007 1.418e-09 0 1.612e-09 0 1.615e-09 0.0007 1.618e-09 0 1.812e-09 0 1.815e-09 0.0007 1.818e-09 0 2.012e-09 0 2.015e-09 0.0007 2.018e-09 0 2.212e-09 0 2.215e-09 0.0007 2.218e-09 0 2.412e-09 0 2.415e-09 0.0007 2.418e-09 0 2.612e-09 0 2.615e-09 0.0007 2.618e-09 0 2.812e-09 0 2.815e-09 0.0007 2.818e-09 0 3.012e-09 0 3.015e-09 0.0007 3.018e-09 0 3.212e-09 0 3.215e-09 0.0007 3.218e-09 0 3.412e-09 0 3.415e-09 0.0007 3.418e-09 0 3.612e-09 0 3.615e-09 0.0007 3.618e-09 0 3.812e-09 0 3.815e-09 0.0007 3.818e-09 0 4.012e-09 0 4.015e-09 0.0007 4.018e-09 0 4.212e-09 0 4.215e-09 0.0007 4.218e-09 0 4.412e-09 0 4.415e-09 0.0007 4.418e-09 0 4.612e-09 0 4.615e-09 0.0007 4.618e-09 0 4.812e-09 0 4.815e-09 0.0007 4.818e-09 0 5.012e-09 0 5.015e-09 0.0007 5.018e-09 0 5.212e-09 0 5.215e-09 0.0007 5.218e-09 0 5.412e-09 0 5.415e-09 0.0007 5.418e-09 0 5.612e-09 0 5.615e-09 0.0007 5.618e-09 0 5.812e-09 0 5.815e-09 0.0007 5.818e-09 0 6.012e-09 0 6.015e-09 0.0007 6.018e-09 0 6.212e-09 0 6.215e-09 0.0007 6.218e-09 0 6.412e-09 0 6.415e-09 0.0007 6.418e-09 0 6.612e-09 0 6.615e-09 0.0007 6.618e-09 0 6.812e-09 0 6.815e-09 0.0007 6.818e-09 0 7.012e-09 0 7.015e-09 0.0007 7.018e-09 0 7.212e-09 0 7.215e-09 0.0007 7.218e-09 0 7.412e-09 0 7.415e-09 0.0007 7.418e-09 0 7.612e-09 0 7.615e-09 0.0007 7.618e-09 0 7.812e-09 0 7.815e-09 0.0007 7.818e-09 0 8.012e-09 0 8.015e-09 0.0007 8.018e-09 0 8.212e-09 0 8.215e-09 0.0007 8.218e-09 0 8.412e-09 0 8.415e-09 0.0007 8.418e-09 0 8.612e-09 0 8.615e-09 0.0007 8.618e-09 0 8.812e-09 0 8.815e-09 0.0007 8.818e-09 0 9.012e-09 0 9.015e-09 0.0007 9.018e-09 0 9.212e-09 0 9.215e-09 0.0007 9.218e-09 0 9.412e-09 0 9.415e-09 0.0007 9.418e-09 0 9.612e-09 0 9.615e-09 0.0007 9.618e-09 0 9.812e-09 0 9.815e-09 0.0007 9.818e-09 0 1.0012e-08 0 1.0015e-08 0.0007 1.0018e-08 0 1.0212e-08 0 1.0215e-08 0.0007 1.0218e-08 0 1.0412e-08 0 1.0415e-08 0.0007 1.0418e-08 0 1.0612e-08 0 1.0615e-08 0.0007 1.0618e-08 0 1.0812e-08 0 1.0815e-08 0.0007 1.0818e-08 0 1.1012e-08 0 1.1015e-08 0.0007 1.1018e-08 0 1.1212e-08 0 1.1215e-08 0.0007 1.1218e-08 0 1.1412e-08 0 1.1415e-08 0.0007 1.1418e-08 0 1.1612e-08 0 1.1615e-08 0.0007 1.1618e-08 0 1.1812e-08 0 1.1815e-08 0.0007 1.1818e-08 0 1.2012e-08 0 1.2015e-08 0.0007 1.2018e-08 0 1.2212e-08 0 1.2215e-08 0.0007 1.2218e-08 0 1.2412e-08 0 1.2415e-08 0.0007 1.2418e-08 0 1.2612e-08 0 1.2615e-08 0.0007 1.2618e-08 0 1.2812e-08 0 1.2815e-08 0.0007 1.2818e-08 0 1.3012e-08 0 1.3015e-08 0.0007 1.3018e-08 0 1.3212e-08 0 1.3215e-08 0.0007 1.3218e-08 0 1.3412e-08 0 1.3415e-08 0.0007 1.3418e-08 0 1.3612e-08 0 1.3615e-08 0.0007 1.3618e-08 0 1.3812e-08 0 1.3815e-08 0.0007 1.3818e-08 0 1.4012e-08 0 1.4015e-08 0.0007 1.4018e-08 0 1.4212e-08 0 1.4215e-08 0.0007 1.4218e-08 0 1.4412e-08 0 1.4415e-08 0.0007 1.4418e-08 0 1.4612e-08 0 1.4615e-08 0.0007 1.4618e-08 0 1.4812e-08 0 1.4815e-08 0.0007 1.4818e-08 0 1.5012e-08 0 1.5015e-08 0.0007 1.5018e-08 0 1.5212e-08 0 1.5215e-08 0.0007 1.5218e-08 0 1.5412e-08 0 1.5415e-08 0.0007 1.5418e-08 0 1.5612e-08 0 1.5615e-08 0.0007 1.5618e-08 0 1.5812e-08 0 1.5815e-08 0.0007 1.5818e-08 0 1.6012e-08 0 1.6015e-08 0.0007 1.6018e-08 0 1.6212e-08 0 1.6215e-08 0.0007 1.6218e-08 0 1.6412e-08 0 1.6415e-08 0.0007 1.6418e-08 0 1.6612e-08 0 1.6615e-08 0.0007 1.6618e-08 0 1.6812e-08 0 1.6815e-08 0.0007 1.6818e-08 0 1.7012e-08 0 1.7015e-08 0.0007 1.7018e-08 0 1.7212e-08 0 1.7215e-08 0.0007 1.7218e-08 0 1.7412e-08 0 1.7415e-08 0.0007 1.7418e-08 0 1.7612e-08 0 1.7615e-08 0.0007 1.7618e-08 0 1.7812e-08 0 1.7815e-08 0.0007 1.7818e-08 0 1.8012e-08 0 1.8015e-08 0.0007 1.8018e-08 0 1.8212e-08 0 1.8215e-08 0.0007 1.8218e-08 0 1.8412e-08 0 1.8415e-08 0.0007 1.8418e-08 0 1.8612e-08 0 1.8615e-08 0.0007 1.8618e-08 0 1.8812e-08 0 1.8815e-08 0.0007 1.8818e-08 0 1.9012e-08 0 1.9015e-08 0.0007 1.9018e-08 0 1.9212e-08 0 1.9215e-08 0.0007 1.9218e-08 0 1.9412e-08 0 1.9415e-08 0.0007 1.9418e-08 0 1.9612e-08 0 1.9615e-08 0.0007 1.9618e-08 0 1.9812e-08 0 1.9815e-08 0.0007 1.9818e-08 0 2.0012e-08 0 2.0015e-08 0.0007 2.0018e-08 0 2.0212e-08 0 2.0215e-08 0.0007 2.0218e-08 0 2.0412e-08 0 2.0415e-08 0.0007 2.0418e-08 0 2.0612e-08 0 2.0615e-08 0.0007 2.0618e-08 0 2.0812e-08 0 2.0815e-08 0.0007 2.0818e-08 0 2.1012e-08 0 2.1015e-08 0.0007 2.1018e-08 0 2.1212e-08 0 2.1215e-08 0.0007 2.1218e-08 0 2.1412e-08 0 2.1415e-08 0.0007 2.1418e-08 0 2.1612e-08 0 2.1615e-08 0.0007 2.1618e-08 0 2.1812e-08 0 2.1815e-08 0.0007 2.1818e-08 0 2.2012e-08 0 2.2015e-08 0.0007 2.2018e-08 0 2.2212e-08 0 2.2215e-08 0.0007 2.2218e-08 0 2.2412e-08 0 2.2415e-08 0.0007 2.2418e-08 0 2.2612e-08 0 2.2615e-08 0.0007 2.2618e-08 0 2.2812e-08 0 2.2815e-08 0.0007 2.2818e-08 0 2.3012e-08 0 2.3015e-08 0.0007 2.3018e-08 0 2.3212e-08 0 2.3215e-08 0.0007 2.3218e-08 0 2.3412e-08 0 2.3415e-08 0.0007 2.3418e-08 0 2.3612e-08 0 2.3615e-08 0.0007 2.3618e-08 0 2.3812e-08 0 2.3815e-08 0.0007 2.3818e-08 0 2.4012e-08 0 2.4015e-08 0.0007 2.4018e-08 0 2.4212e-08 0 2.4215e-08 0.0007 2.4218e-08 0 2.4412e-08 0 2.4415e-08 0.0007 2.4418e-08 0 2.4612e-08 0 2.4615e-08 0.0007 2.4618e-08 0 2.4812e-08 0 2.4815e-08 0.0007 2.4818e-08 0 2.5012e-08 0 2.5015e-08 0.0007 2.5018e-08 0 2.5212e-08 0 2.5215e-08 0.0007 2.5218e-08 0 2.5412e-08 0 2.5415e-08 0.0007 2.5418e-08 0 2.5612e-08 0 2.5615e-08 0.0007 2.5618e-08 0 2.5812e-08 0 2.5815e-08 0.0007 2.5818e-08 0 2.6012e-08 0 2.6015e-08 0.0007 2.6018e-08 0 2.6212e-08 0 2.6215e-08 0.0007 2.6218e-08 0 2.6412e-08 0 2.6415e-08 0.0007 2.6418e-08 0 2.6612e-08 0 2.6615e-08 0.0007 2.6618e-08 0 2.6812e-08 0 2.6815e-08 0.0007 2.6818e-08 0 2.7012e-08 0 2.7015e-08 0.0007 2.7018e-08 0 2.7212e-08 0 2.7215e-08 0.0007 2.7218e-08 0 2.7412e-08 0 2.7415e-08 0.0007 2.7418e-08 0 2.7612e-08 0 2.7615e-08 0.0007 2.7618e-08 0 2.7812e-08 0 2.7815e-08 0.0007 2.7818e-08 0 2.8012e-08 0 2.8015e-08 0.0007 2.8018e-08 0 2.8212e-08 0 2.8215e-08 0.0007 2.8218e-08 0 2.8412e-08 0 2.8415e-08 0.0007 2.8418e-08 0 2.8612e-08 0 2.8615e-08 0.0007 2.8618e-08 0 2.8812e-08 0 2.8815e-08 0.0007 2.8818e-08 0 2.9012e-08 0 2.9015e-08 0.0007 2.9018e-08 0 2.9212e-08 0 2.9215e-08 0.0007 2.9218e-08 0 2.9412e-08 0 2.9415e-08 0.0007 2.9418e-08 0 2.9612e-08 0 2.9615e-08 0.0007 2.9618e-08 0 2.9812e-08 0 2.9815e-08 0.0007 2.9818e-08 0 3.0012e-08 0 3.0015e-08 0.0007 3.0018e-08 0 3.0212e-08 0 3.0215e-08 0.0007 3.0218e-08 0 3.0412e-08 0 3.0415e-08 0.0007 3.0418e-08 0 3.0612e-08 0 3.0615e-08 0.0007 3.0618e-08 0 3.0812e-08 0 3.0815e-08 0.0007 3.0818e-08 0 3.1012e-08 0 3.1015e-08 0.0007 3.1018e-08 0 3.1212e-08 0 3.1215e-08 0.0007 3.1218e-08 0 3.1412e-08 0 3.1415e-08 0.0007 3.1418e-08 0 3.1612e-08 0 3.1615e-08 0.0007 3.1618e-08 0 3.1812e-08 0 3.1815e-08 0.0007 3.1818e-08 0 3.2012e-08 0 3.2015e-08 0.0007 3.2018e-08 0 3.2212e-08 0 3.2215e-08 0.0007 3.2218e-08 0 3.2412e-08 0 3.2415e-08 0.0007 3.2418e-08 0 3.2612e-08 0 3.2615e-08 0.0007 3.2618e-08 0 3.2812e-08 0 3.2815e-08 0.0007 3.2818e-08 0 3.3012e-08 0 3.3015e-08 0.0007 3.3018e-08 0 3.3212e-08 0 3.3215e-08 0.0007 3.3218e-08 0 3.3412e-08 0 3.3415e-08 0.0007 3.3418e-08 0 3.3612e-08 0 3.3615e-08 0.0007 3.3618e-08 0 3.3812e-08 0 3.3815e-08 0.0007 3.3818e-08 0 3.4012e-08 0 3.4015e-08 0.0007 3.4018e-08 0 3.4212e-08 0 3.4215e-08 0.0007 3.4218e-08 0 3.4412e-08 0 3.4415e-08 0.0007 3.4418e-08 0 3.4612e-08 0 3.4615e-08 0.0007 3.4618e-08 0 3.4812e-08 0 3.4815e-08 0.0007 3.4818e-08 0 3.5012e-08 0 3.5015e-08 0.0007 3.5018e-08 0 3.5212e-08 0 3.5215e-08 0.0007 3.5218e-08 0 3.5412e-08 0 3.5415e-08 0.0007 3.5418e-08 0 3.5612e-08 0 3.5615e-08 0.0007 3.5618e-08 0 3.5812e-08 0 3.5815e-08 0.0007 3.5818e-08 0 3.6012e-08 0 3.6015e-08 0.0007 3.6018e-08 0 3.6212e-08 0 3.6215e-08 0.0007 3.6218e-08 0 3.6412e-08 0 3.6415e-08 0.0007 3.6418e-08 0 3.6612e-08 0 3.6615e-08 0.0007 3.6618e-08 0 3.6812e-08 0 3.6815e-08 0.0007 3.6818e-08 0 3.7012e-08 0 3.7015e-08 0.0007 3.7018e-08 0 3.7212e-08 0 3.7215e-08 0.0007 3.7218e-08 0 3.7412e-08 0 3.7415e-08 0.0007 3.7418e-08 0 3.7612e-08 0 3.7615e-08 0.0007 3.7618e-08 0 3.7812e-08 0 3.7815e-08 0.0007 3.7818e-08 0 3.8012e-08 0 3.8015e-08 0.0007 3.8018e-08 0 3.8212e-08 0 3.8215e-08 0.0007 3.8218e-08 0 3.8412e-08 0 3.8415e-08 0.0007 3.8418e-08 0 3.8612e-08 0 3.8615e-08 0.0007 3.8618e-08 0 3.8812e-08 0 3.8815e-08 0.0007 3.8818e-08 0 3.9012e-08 0 3.9015e-08 0.0007 3.9018e-08 0 3.9212e-08 0 3.9215e-08 0.0007 3.9218e-08 0 3.9412e-08 0 3.9415e-08 0.0007 3.9418e-08 0 3.9612e-08 0 3.9615e-08 0.0007 3.9618e-08 0 3.9812e-08 0 3.9815e-08 0.0007 3.9818e-08 0 4.0012e-08 0 4.0015e-08 0.0007 4.0018e-08 0 4.0212e-08 0 4.0215e-08 0.0007 4.0218e-08 0 4.0412e-08 0 4.0415e-08 0.0007 4.0418e-08 0 4.0612e-08 0 4.0615e-08 0.0007 4.0618e-08 0 4.0812e-08 0 4.0815e-08 0.0007 4.0818e-08 0 4.1012e-08 0 4.1015e-08 0.0007 4.1018e-08 0 4.1212e-08 0 4.1215e-08 0.0007 4.1218e-08 0 4.1412e-08 0 4.1415e-08 0.0007 4.1418e-08 0 4.1612e-08 0 4.1615e-08 0.0007 4.1618e-08 0 4.1812e-08 0 4.1815e-08 0.0007 4.1818e-08 0 4.2012e-08 0 4.2015e-08 0.0007 4.2018e-08 0 4.2212e-08 0 4.2215e-08 0.0007 4.2218e-08 0 4.2412e-08 0 4.2415e-08 0.0007 4.2418e-08 0 4.2612e-08 0 4.2615e-08 0.0007 4.2618e-08 0 4.2812e-08 0 4.2815e-08 0.0007 4.2818e-08 0 4.3012e-08 0 4.3015e-08 0.0007 4.3018e-08 0 4.3212e-08 0 4.3215e-08 0.0007 4.3218e-08 0 4.3412e-08 0 4.3415e-08 0.0007 4.3418e-08 0 4.3612e-08 0 4.3615e-08 0.0007 4.3618e-08 0 4.3812e-08 0 4.3815e-08 0.0007 4.3818e-08 0 4.4012e-08 0 4.4015e-08 0.0007 4.4018e-08 0 4.4212e-08 0 4.4215e-08 0.0007 4.4218e-08 0 4.4412e-08 0 4.4415e-08 0.0007 4.4418e-08 0 4.4612e-08 0 4.4615e-08 0.0007 4.4618e-08 0 4.4812e-08 0 4.4815e-08 0.0007 4.4818e-08 0 4.5012e-08 0 4.5015e-08 0.0007 4.5018e-08 0 4.5212e-08 0 4.5215e-08 0.0007 4.5218e-08 0 4.5412e-08 0 4.5415e-08 0.0007 4.5418e-08 0 4.5612e-08 0 4.5615e-08 0.0007 4.5618e-08 0 4.5812e-08 0 4.5815e-08 0.0007 4.5818e-08 0 4.6012e-08 0 4.6015e-08 0.0007 4.6018e-08 0 4.6212e-08 0 4.6215e-08 0.0007 4.6218e-08 0 4.6412e-08 0 4.6415e-08 0.0007 4.6418e-08 0 4.6612e-08 0 4.6615e-08 0.0007 4.6618e-08 0 4.6812e-08 0 4.6815e-08 0.0007 4.6818e-08 0 4.7012e-08 0 4.7015e-08 0.0007 4.7018e-08 0 4.7212e-08 0 4.7215e-08 0.0007 4.7218e-08 0 4.7412e-08 0 4.7415e-08 0.0007 4.7418e-08 0 4.7612e-08 0 4.7615e-08 0.0007 4.7618e-08 0 4.7812e-08 0 4.7815e-08 0.0007 4.7818e-08 0 4.8012e-08 0 4.8015e-08 0.0007 4.8018e-08 0 4.8212e-08 0 4.8215e-08 0.0007 4.8218e-08 0 4.8412e-08 0 4.8415e-08 0.0007 4.8418e-08 0 4.8612e-08 0 4.8615e-08 0.0007 4.8618e-08 0 4.8812e-08 0 4.8815e-08 0.0007 4.8818e-08 0 4.9012e-08 0 4.9015e-08 0.0007 4.9018e-08 0 4.9212e-08 0 4.9215e-08 0.0007 4.9218e-08 0 4.9412e-08 0 4.9415e-08 0.0007 4.9418e-08 0 4.9612e-08 0 4.9615e-08 0.0007 4.9618e-08 0 4.9812e-08 0 4.9815e-08 0.0007 4.9818e-08 0 5.0012e-08 0 5.0015e-08 0.0007 5.0018e-08 0 5.0212e-08 0 5.0215e-08 0.0007 5.0218e-08 0 5.0412e-08 0 5.0415e-08 0.0007 5.0418e-08 0 5.0612e-08 0 5.0615e-08 0.0007 5.0618e-08 0 5.0812e-08 0 5.0815e-08 0.0007 5.0818e-08 0 5.1012e-08 0 5.1015e-08 0.0007 5.1018e-08 0 5.1212e-08 0 5.1215e-08 0.0007 5.1218e-08 0 5.1412e-08 0 5.1415e-08 0.0007 5.1418e-08 0 5.1612e-08 0 5.1615e-08 0.0007 5.1618e-08 0 5.1812e-08 0 5.1815e-08 0.0007 5.1818e-08 0 5.2012e-08 0 5.2015e-08 0.0007 5.2018e-08 0 5.2212e-08 0 5.2215e-08 0.0007 5.2218e-08 0 5.2412e-08 0 5.2415e-08 0.0007 5.2418e-08 0 5.2612e-08 0 5.2615e-08 0.0007 5.2618e-08 0 5.2812e-08 0 5.2815e-08 0.0007 5.2818e-08 0 5.3012e-08 0 5.3015e-08 0.0007 5.3018e-08 0 5.3212e-08 0 5.3215e-08 0.0007 5.3218e-08 0 5.3412e-08 0 5.3415e-08 0.0007 5.3418e-08 0 5.3612e-08 0 5.3615e-08 0.0007 5.3618e-08 0 5.3812e-08 0 5.3815e-08 0.0007 5.3818e-08 0 5.4012e-08 0 5.4015e-08 0.0007 5.4018e-08 0 5.4212e-08 0 5.4215e-08 0.0007 5.4218e-08 0 5.4412e-08 0 5.4415e-08 0.0007 5.4418e-08 0 5.4612e-08 0 5.4615e-08 0.0007 5.4618e-08 0 5.4812e-08 0 5.4815e-08 0.0007 5.4818e-08 0 5.5012e-08 0 5.5015e-08 0.0007 5.5018e-08 0 5.5212e-08 0 5.5215e-08 0.0007 5.5218e-08 0 5.5412e-08 0 5.5415e-08 0.0007 5.5418e-08 0 5.5612e-08 0 5.5615e-08 0.0007 5.5618e-08 0 5.5812e-08 0 5.5815e-08 0.0007 5.5818e-08 0 5.6012e-08 0 5.6015e-08 0.0007 5.6018e-08 0 5.6212e-08 0 5.6215e-08 0.0007 5.6218e-08 0 5.6412e-08 0 5.6415e-08 0.0007 5.6418e-08 0 5.6612e-08 0 5.6615e-08 0.0007 5.6618e-08 0 5.6812e-08 0 5.6815e-08 0.0007 5.6818e-08 0 5.7012e-08 0 5.7015e-08 0.0007 5.7018e-08 0 5.7212e-08 0 5.7215e-08 0.0007 5.7218e-08 0 5.7412e-08 0 5.7415e-08 0.0007 5.7418e-08 0 5.7612e-08 0 5.7615e-08 0.0007 5.7618e-08 0 5.7812e-08 0 5.7815e-08 0.0007 5.7818e-08 0 5.8012e-08 0 5.8015e-08 0.0007 5.8018e-08 0 5.8212e-08 0 5.8215e-08 0.0007 5.8218e-08 0 5.8412e-08 0 5.8415e-08 0.0007 5.8418e-08 0 5.8612e-08 0 5.8615e-08 0.0007 5.8618e-08 0 5.8812e-08 0 5.8815e-08 0.0007 5.8818e-08 0 5.9012e-08 0 5.9015e-08 0.0007 5.9018e-08 0 5.9212e-08 0 5.9215e-08 0.0007 5.9218e-08 0 5.9412e-08 0 5.9415e-08 0.0007 5.9418e-08 0 5.9612e-08 0 5.9615e-08 0.0007 5.9618e-08 0 5.9812e-08 0 5.9815e-08 0.0007 5.9818e-08 0 6.0012e-08 0 6.0015e-08 0.0007 6.0018e-08 0 6.0212e-08 0 6.0215e-08 0.0007 6.0218e-08 0 6.0412e-08 0 6.0415e-08 0.0007 6.0418e-08 0 6.0612e-08 0 6.0615e-08 0.0007 6.0618e-08 0 6.0812e-08 0 6.0815e-08 0.0007 6.0818e-08 0 6.1012e-08 0 6.1015e-08 0.0007 6.1018e-08 0 6.1212e-08 0 6.1215e-08 0.0007 6.1218e-08 0 6.1412e-08 0 6.1415e-08 0.0007 6.1418e-08 0 6.1612e-08 0 6.1615e-08 0.0007 6.1618e-08 0 6.1812e-08 0 6.1815e-08 0.0007 6.1818e-08 0 6.2012e-08 0 6.2015e-08 0.0007 6.2018e-08 0 6.2212e-08 0 6.2215e-08 0.0007 6.2218e-08 0 6.2412e-08 0 6.2415e-08 0.0007 6.2418e-08 0 6.2612e-08 0 6.2615e-08 0.0007 6.2618e-08 0 6.2812e-08 0 6.2815e-08 0.0007 6.2818e-08 0 6.3012e-08 0 6.3015e-08 0.0007 6.3018e-08 0 6.3212e-08 0 6.3215e-08 0.0007 6.3218e-08 0 6.3412e-08 0 6.3415e-08 0.0007 6.3418e-08 0 6.3612e-08 0 6.3615e-08 0.0007 6.3618e-08 0 6.3812e-08 0 6.3815e-08 0.0007 6.3818e-08 0 6.4012e-08 0 6.4015e-08 0.0007 6.4018e-08 0 6.4212e-08 0 6.4215e-08 0.0007 6.4218e-08 0 6.4412e-08 0 6.4415e-08 0.0007 6.4418e-08 0 6.4612e-08 0 6.4615e-08 0.0007 6.4618e-08 0 6.4812e-08 0 6.4815e-08 0.0007 6.4818e-08 0 6.5012e-08 0 6.5015e-08 0.0007 6.5018e-08 0 6.5212e-08 0 6.5215e-08 0.0007 6.5218e-08 0 6.5412e-08 0 6.5415e-08 0.0007 6.5418e-08 0 6.5612e-08 0 6.5615e-08 0.0007 6.5618e-08 0 6.5812e-08 0 6.5815e-08 0.0007 6.5818e-08 0 6.6012e-08 0 6.6015e-08 0.0007 6.6018e-08 0 6.6212e-08 0 6.6215e-08 0.0007 6.6218e-08 0 6.6412e-08 0 6.6415e-08 0.0007 6.6418e-08 0 6.6612e-08 0 6.6615e-08 0.0007 6.6618e-08 0 6.6812e-08 0 6.6815e-08 0.0007 6.6818e-08 0 6.7012e-08 0 6.7015e-08 0.0007 6.7018e-08 0 6.7212e-08 0 6.7215e-08 0.0007 6.7218e-08 0 6.7412e-08 0 6.7415e-08 0.0007 6.7418e-08 0 6.7612e-08 0 6.7615e-08 0.0007 6.7618e-08 0 6.7812e-08 0 6.7815e-08 0.0007 6.7818e-08 0 6.8012e-08 0 6.8015e-08 0.0007 6.8018e-08 0 6.8212e-08 0 6.8215e-08 0.0007 6.8218e-08 0 6.8412e-08 0 6.8415e-08 0.0007 6.8418e-08 0 6.8612e-08 0 6.8615e-08 0.0007 6.8618e-08 0 6.8812e-08 0 6.8815e-08 0.0007 6.8818e-08 0 6.9012e-08 0 6.9015e-08 0.0007 6.9018e-08 0 6.9212e-08 0 6.9215e-08 0.0007 6.9218e-08 0 6.9412e-08 0 6.9415e-08 0.0007 6.9418e-08 0 6.9612e-08 0 6.9615e-08 0.0007 6.9618e-08 0 6.9812e-08 0 6.9815e-08 0.0007 6.9818e-08 0 7.0012e-08 0 7.0015e-08 0.0007 7.0018e-08 0 7.0212e-08 0 7.0215e-08 0.0007 7.0218e-08 0 7.0412e-08 0 7.0415e-08 0.0007 7.0418e-08 0 7.0612e-08 0 7.0615e-08 0.0007 7.0618e-08 0 7.0812e-08 0 7.0815e-08 0.0007 7.0818e-08 0 7.1012e-08 0 7.1015e-08 0.0007 7.1018e-08 0 7.1212e-08 0 7.1215e-08 0.0007 7.1218e-08 0 7.1412e-08 0 7.1415e-08 0.0007 7.1418e-08 0 7.1612e-08 0 7.1615e-08 0.0007 7.1618e-08 0 7.1812e-08 0 7.1815e-08 0.0007 7.1818e-08 0 7.2012e-08 0 7.2015e-08 0.0007 7.2018e-08 0 7.2212e-08 0 7.2215e-08 0.0007 7.2218e-08 0 7.2412e-08 0 7.2415e-08 0.0007 7.2418e-08 0 7.2612e-08 0 7.2615e-08 0.0007 7.2618e-08 0 7.2812e-08 0 7.2815e-08 0.0007 7.2818e-08 0 7.3012e-08 0 7.3015e-08 0.0007 7.3018e-08 0 7.3212e-08 0 7.3215e-08 0.0007 7.3218e-08 0 7.3412e-08 0 7.3415e-08 0.0007 7.3418e-08 0 7.3612e-08 0 7.3615e-08 0.0007 7.3618e-08 0 7.3812e-08 0 7.3815e-08 0.0007 7.3818e-08 0 7.4012e-08 0 7.4015e-08 0.0007 7.4018e-08 0 7.4212e-08 0 7.4215e-08 0.0007 7.4218e-08 0 7.4412e-08 0 7.4415e-08 0.0007 7.4418e-08 0 7.4612e-08 0 7.4615e-08 0.0007 7.4618e-08 0 7.4812e-08 0 7.4815e-08 0.0007 7.4818e-08 0 7.5012e-08 0 7.5015e-08 0.0007 7.5018e-08 0 7.5212e-08 0 7.5215e-08 0.0007 7.5218e-08 0 7.5412e-08 0 7.5415e-08 0.0007 7.5418e-08 0 7.5612e-08 0 7.5615e-08 0.0007 7.5618e-08 0 7.5812e-08 0 7.5815e-08 0.0007 7.5818e-08 0 7.6012e-08 0 7.6015e-08 0.0007 7.6018e-08 0 7.6212e-08 0 7.6215e-08 0.0007 7.6218e-08 0 7.6412e-08 0 7.6415e-08 0.0007 7.6418e-08 0 7.6612e-08 0 7.6615e-08 0.0007 7.6618e-08 0 7.6812e-08 0 7.6815e-08 0.0007 7.6818e-08 0 7.7012e-08 0 7.7015e-08 0.0007 7.7018e-08 0 7.7212e-08 0 7.7215e-08 0.0007 7.7218e-08 0 7.7412e-08 0 7.7415e-08 0.0007 7.7418e-08 0 7.7612e-08 0 7.7615e-08 0.0007 7.7618e-08 0 7.7812e-08 0 7.7815e-08 0.0007 7.7818e-08 0 7.8012e-08 0 7.8015e-08 0.0007 7.8018e-08 0 7.8212e-08 0 7.8215e-08 0.0007 7.8218e-08 0 7.8412e-08 0 7.8415e-08 0.0007 7.8418e-08 0 7.8612e-08 0 7.8615e-08 0.0007 7.8618e-08 0 7.8812e-08 0 7.8815e-08 0.0007 7.8818e-08 0 7.9012e-08 0 7.9015e-08 0.0007 7.9018e-08 0 7.9212e-08 0 7.9215e-08 0.0007 7.9218e-08 0 7.9412e-08 0 7.9415e-08 0.0007 7.9418e-08 0 7.9612e-08 0 7.9615e-08 0.0007 7.9618e-08 0)
L_DFF_IP3_01|1 IP3_0_OUT _DFF_IP3_01|A1  2.067833848e-12
L_DFF_IP3_01|2 _DFF_IP3_01|A1 _DFF_IP3_01|A2  4.135667696e-12
L_DFF_IP3_01|3 _DFF_IP3_01|A3 _DFF_IP3_01|A4  8.271335392e-12
L_DFF_IP3_01|T D03 _DFF_IP3_01|T1  2.067833848e-12
L_DFF_IP3_01|4 _DFF_IP3_01|T1 _DFF_IP3_01|T2  4.135667696e-12
L_DFF_IP3_01|5 _DFF_IP3_01|A4 _DFF_IP3_01|Q1  4.135667696e-12
L_DFF_IP3_01|6 _DFF_IP3_01|Q1 IP3_1_OUT  2.067833848e-12
IT08|T 0 T08  PWL(0 0 7e-12 0 1e-11 0.0014 1.3e-11 0 2.07e-10 0 2.1e-10 0.0014 2.13e-10 0 4.07e-10 0 4.1e-10 0.0014 4.13e-10 0 6.07e-10 0 6.1e-10 0.0014 6.13e-10 0 8.07e-10 0 8.1e-10 0.0014 8.13e-10 0 1.007e-09 0 1.01e-09 0.0014 1.013e-09 0 1.207e-09 0 1.21e-09 0.0014 1.213e-09 0 1.407e-09 0 1.41e-09 0.0014 1.413e-09 0 1.607e-09 0 1.61e-09 0.0014 1.613e-09 0 1.807e-09 0 1.81e-09 0.0014 1.813e-09 0 2.007e-09 0 2.01e-09 0.0014 2.013e-09 0 2.207e-09 0 2.21e-09 0.0014 2.213e-09 0 2.407e-09 0 2.41e-09 0.0014 2.413e-09 0 2.607e-09 0 2.61e-09 0.0014 2.613e-09 0 2.807e-09 0 2.81e-09 0.0014 2.813e-09 0 3.007e-09 0 3.01e-09 0.0014 3.013e-09 0 3.207e-09 0 3.21e-09 0.0014 3.213e-09 0 3.407e-09 0 3.41e-09 0.0014 3.413e-09 0 3.607e-09 0 3.61e-09 0.0014 3.613e-09 0 3.807e-09 0 3.81e-09 0.0014 3.813e-09 0 4.007e-09 0 4.01e-09 0.0014 4.013e-09 0 4.207e-09 0 4.21e-09 0.0014 4.213e-09 0 4.407e-09 0 4.41e-09 0.0014 4.413e-09 0 4.607e-09 0 4.61e-09 0.0014 4.613e-09 0 4.807e-09 0 4.81e-09 0.0014 4.813e-09 0 5.007e-09 0 5.01e-09 0.0014 5.013e-09 0 5.207e-09 0 5.21e-09 0.0014 5.213e-09 0 5.407e-09 0 5.41e-09 0.0014 5.413e-09 0 5.607e-09 0 5.61e-09 0.0014 5.613e-09 0 5.807e-09 0 5.81e-09 0.0014 5.813e-09 0 6.007e-09 0 6.01e-09 0.0014 6.013e-09 0 6.207e-09 0 6.21e-09 0.0014 6.213e-09 0 6.407e-09 0 6.41e-09 0.0014 6.413e-09 0 6.607e-09 0 6.61e-09 0.0014 6.613e-09 0 6.807e-09 0 6.81e-09 0.0014 6.813e-09 0 7.007e-09 0 7.01e-09 0.0014 7.013e-09 0 7.207e-09 0 7.21e-09 0.0014 7.213e-09 0 7.407e-09 0 7.41e-09 0.0014 7.413e-09 0 7.607e-09 0 7.61e-09 0.0014 7.613e-09 0 7.807e-09 0 7.81e-09 0.0014 7.813e-09 0 8.007e-09 0 8.01e-09 0.0014 8.013e-09 0 8.207e-09 0 8.21e-09 0.0014 8.213e-09 0 8.407e-09 0 8.41e-09 0.0014 8.413e-09 0 8.607e-09 0 8.61e-09 0.0014 8.613e-09 0 8.807e-09 0 8.81e-09 0.0014 8.813e-09 0 9.007e-09 0 9.01e-09 0.0014 9.013e-09 0 9.207e-09 0 9.21e-09 0.0014 9.213e-09 0 9.407e-09 0 9.41e-09 0.0014 9.413e-09 0 9.607e-09 0 9.61e-09 0.0014 9.613e-09 0 9.807e-09 0 9.81e-09 0.0014 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0014 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0014 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0014 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0014 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0014 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0014 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0014 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0014 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0014 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0014 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0014 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0014 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0014 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0014 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0014 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0014 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0014 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0014 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0014 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0014 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0014 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0014 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0014 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0014 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0014 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0014 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0014 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0014 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0014 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0014 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0014 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0014 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0014 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0014 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0014 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0014 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0014 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0014 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0014 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0014 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0014 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0014 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0014 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0014 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0014 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0014 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0014 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0014 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0014 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0014 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0014 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0014 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0014 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0014 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0014 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0014 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0014 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0014 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0014 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0014 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0014 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0014 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0014 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0014 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0014 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0014 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0014 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0014 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0014 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0014 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0014 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0014 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0014 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0014 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0014 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0014 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0014 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0014 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0014 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0014 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0014 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0014 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0014 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0014 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0014 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0014 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0014 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0014 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0014 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0014 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0014 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0014 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0014 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0014 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0014 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0014 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0014 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0014 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0014 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0014 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0014 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0014 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0014 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0014 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0014 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0014 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0014 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0014 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0014 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0014 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0014 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0014 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0014 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0014 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0014 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0014 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0014 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0014 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0014 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0014 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0014 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0014 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0014 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0014 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0014 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0014 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0014 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0014 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0014 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0014 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0014 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0014 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0014 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0014 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0014 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0014 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0014 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0014 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0014 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0014 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0014 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0014 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0014 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0014 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0014 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0014 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0014 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0014 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0014 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0014 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0014 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0014 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0014 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0014 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0014 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0014 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0014 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0014 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0014 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0014 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0014 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0014 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0014 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0014 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0014 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0014 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0014 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0014 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0014 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0014 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0014 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0014 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0014 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0014 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0014 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0014 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0014 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0014 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0014 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0014 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0014 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0014 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0014 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0014 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0014 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0014 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0014 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0014 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0014 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0014 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0014 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0014 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0014 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0014 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0014 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0014 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0014 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0014 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0014 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0014 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0014 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0014 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0014 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0014 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0014 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0014 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0014 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0014 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0014 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0014 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0014 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0014 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0014 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0014 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0014 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0014 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0014 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0014 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0014 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0014 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0014 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0014 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0014 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0014 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0014 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0014 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0014 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0014 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0014 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0014 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0014 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0014 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0014 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0014 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0014 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0014 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0014 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0014 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0014 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0014 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0014 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0014 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0014 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0014 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0014 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0014 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0014 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0014 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0014 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0014 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0014 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0014 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0014 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0014 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0014 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0014 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0014 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0014 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0014 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0014 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0014 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0014 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0014 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0014 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0014 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0014 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0014 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0014 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0014 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0014 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0014 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0014 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0014 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0014 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0014 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0014 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0014 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0014 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0014 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0014 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0014 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0014 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0014 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0014 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0014 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0014 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0014 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0014 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0014 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0014 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0014 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0014 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0014 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0014 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0014 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0014 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0014 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0014 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0014 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0014 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0014 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0014 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0014 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0014 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0014 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0014 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0014 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0014 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0014 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0014 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0014 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0014 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0014 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0014 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0014 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0014 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0014 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0014 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0014 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0014 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0014 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0014 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0014 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0014 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0014 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0014 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0014 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0014 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0014 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0014 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0014 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0014 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0014 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0014 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0014 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0014 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0014 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0014 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0014 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0014 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0014 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0014 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0014 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0014 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0014 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0014 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0014 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0014 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0014 7.9613e-08 0)
IT09|T 0 T09  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_PG1_12|1 G1_1_TO1 _PG1_12|A1  2.067833848e-12
L_PG1_12|2 _PG1_12|A1 _PG1_12|A2  4.135667696e-12
L_PG1_12|3 _PG1_12|A3 _PG1_12|A4  8.271335392e-12
L_PG1_12|T T09 _PG1_12|T1  2.067833848e-12
L_PG1_12|4 _PG1_12|T1 _PG1_12|T2  4.135667696e-12
L_PG1_12|5 _PG1_12|A4 _PG1_12|Q1  4.135667696e-12
L_PG1_12|6 _PG1_12|Q1 G1_2  2.067833848e-12
IT10|T 0 T10  PWL(0 0 7e-12 0 1e-11 0.0014 1.3e-11 0 2.07e-10 0 2.1e-10 0.0014 2.13e-10 0 4.07e-10 0 4.1e-10 0.0014 4.13e-10 0 6.07e-10 0 6.1e-10 0.0014 6.13e-10 0 8.07e-10 0 8.1e-10 0.0014 8.13e-10 0 1.007e-09 0 1.01e-09 0.0014 1.013e-09 0 1.207e-09 0 1.21e-09 0.0014 1.213e-09 0 1.407e-09 0 1.41e-09 0.0014 1.413e-09 0 1.607e-09 0 1.61e-09 0.0014 1.613e-09 0 1.807e-09 0 1.81e-09 0.0014 1.813e-09 0 2.007e-09 0 2.01e-09 0.0014 2.013e-09 0 2.207e-09 0 2.21e-09 0.0014 2.213e-09 0 2.407e-09 0 2.41e-09 0.0014 2.413e-09 0 2.607e-09 0 2.61e-09 0.0014 2.613e-09 0 2.807e-09 0 2.81e-09 0.0014 2.813e-09 0 3.007e-09 0 3.01e-09 0.0014 3.013e-09 0 3.207e-09 0 3.21e-09 0.0014 3.213e-09 0 3.407e-09 0 3.41e-09 0.0014 3.413e-09 0 3.607e-09 0 3.61e-09 0.0014 3.613e-09 0 3.807e-09 0 3.81e-09 0.0014 3.813e-09 0 4.007e-09 0 4.01e-09 0.0014 4.013e-09 0 4.207e-09 0 4.21e-09 0.0014 4.213e-09 0 4.407e-09 0 4.41e-09 0.0014 4.413e-09 0 4.607e-09 0 4.61e-09 0.0014 4.613e-09 0 4.807e-09 0 4.81e-09 0.0014 4.813e-09 0 5.007e-09 0 5.01e-09 0.0014 5.013e-09 0 5.207e-09 0 5.21e-09 0.0014 5.213e-09 0 5.407e-09 0 5.41e-09 0.0014 5.413e-09 0 5.607e-09 0 5.61e-09 0.0014 5.613e-09 0 5.807e-09 0 5.81e-09 0.0014 5.813e-09 0 6.007e-09 0 6.01e-09 0.0014 6.013e-09 0 6.207e-09 0 6.21e-09 0.0014 6.213e-09 0 6.407e-09 0 6.41e-09 0.0014 6.413e-09 0 6.607e-09 0 6.61e-09 0.0014 6.613e-09 0 6.807e-09 0 6.81e-09 0.0014 6.813e-09 0 7.007e-09 0 7.01e-09 0.0014 7.013e-09 0 7.207e-09 0 7.21e-09 0.0014 7.213e-09 0 7.407e-09 0 7.41e-09 0.0014 7.413e-09 0 7.607e-09 0 7.61e-09 0.0014 7.613e-09 0 7.807e-09 0 7.81e-09 0.0014 7.813e-09 0 8.007e-09 0 8.01e-09 0.0014 8.013e-09 0 8.207e-09 0 8.21e-09 0.0014 8.213e-09 0 8.407e-09 0 8.41e-09 0.0014 8.413e-09 0 8.607e-09 0 8.61e-09 0.0014 8.613e-09 0 8.807e-09 0 8.81e-09 0.0014 8.813e-09 0 9.007e-09 0 9.01e-09 0.0014 9.013e-09 0 9.207e-09 0 9.21e-09 0.0014 9.213e-09 0 9.407e-09 0 9.41e-09 0.0014 9.413e-09 0 9.607e-09 0 9.61e-09 0.0014 9.613e-09 0 9.807e-09 0 9.81e-09 0.0014 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0014 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0014 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0014 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0014 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0014 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0014 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0014 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0014 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0014 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0014 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0014 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0014 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0014 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0014 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0014 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0014 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0014 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0014 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0014 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0014 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0014 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0014 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0014 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0014 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0014 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0014 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0014 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0014 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0014 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0014 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0014 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0014 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0014 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0014 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0014 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0014 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0014 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0014 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0014 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0014 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0014 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0014 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0014 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0014 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0014 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0014 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0014 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0014 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0014 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0014 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0014 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0014 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0014 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0014 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0014 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0014 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0014 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0014 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0014 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0014 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0014 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0014 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0014 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0014 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0014 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0014 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0014 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0014 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0014 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0014 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0014 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0014 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0014 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0014 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0014 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0014 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0014 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0014 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0014 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0014 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0014 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0014 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0014 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0014 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0014 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0014 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0014 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0014 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0014 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0014 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0014 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0014 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0014 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0014 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0014 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0014 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0014 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0014 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0014 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0014 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0014 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0014 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0014 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0014 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0014 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0014 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0014 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0014 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0014 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0014 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0014 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0014 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0014 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0014 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0014 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0014 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0014 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0014 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0014 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0014 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0014 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0014 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0014 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0014 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0014 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0014 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0014 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0014 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0014 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0014 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0014 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0014 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0014 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0014 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0014 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0014 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0014 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0014 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0014 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0014 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0014 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0014 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0014 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0014 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0014 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0014 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0014 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0014 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0014 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0014 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0014 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0014 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0014 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0014 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0014 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0014 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0014 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0014 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0014 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0014 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0014 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0014 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0014 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0014 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0014 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0014 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0014 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0014 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0014 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0014 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0014 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0014 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0014 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0014 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0014 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0014 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0014 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0014 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0014 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0014 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0014 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0014 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0014 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0014 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0014 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0014 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0014 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0014 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0014 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0014 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0014 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0014 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0014 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0014 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0014 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0014 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0014 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0014 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0014 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0014 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0014 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0014 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0014 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0014 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0014 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0014 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0014 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0014 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0014 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0014 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0014 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0014 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0014 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0014 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0014 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0014 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0014 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0014 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0014 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0014 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0014 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0014 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0014 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0014 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0014 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0014 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0014 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0014 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0014 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0014 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0014 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0014 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0014 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0014 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0014 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0014 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0014 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0014 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0014 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0014 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0014 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0014 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0014 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0014 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0014 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0014 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0014 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0014 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0014 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0014 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0014 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0014 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0014 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0014 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0014 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0014 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0014 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0014 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0014 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0014 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0014 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0014 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0014 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0014 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0014 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0014 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0014 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0014 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0014 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0014 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0014 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0014 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0014 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0014 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0014 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0014 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0014 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0014 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0014 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0014 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0014 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0014 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0014 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0014 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0014 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0014 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0014 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0014 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0014 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0014 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0014 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0014 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0014 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0014 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0014 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0014 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0014 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0014 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0014 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0014 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0014 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0014 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0014 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0014 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0014 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0014 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0014 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0014 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0014 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0014 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0014 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0014 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0014 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0014 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0014 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0014 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0014 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0014 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0014 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0014 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0014 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0014 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0014 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0014 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0014 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0014 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0014 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0014 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0014 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0014 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0014 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0014 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0014 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0014 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0014 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0014 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0014 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0014 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0014 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0014 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0014 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0014 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0014 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0014 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0014 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0014 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0014 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0014 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0014 7.9613e-08 0)
IT11|T 0 T11  PWL(0 0 7e-12 0 1e-11 0.0014 1.3e-11 0 2.07e-10 0 2.1e-10 0.0014 2.13e-10 0 4.07e-10 0 4.1e-10 0.0014 4.13e-10 0 6.07e-10 0 6.1e-10 0.0014 6.13e-10 0 8.07e-10 0 8.1e-10 0.0014 8.13e-10 0 1.007e-09 0 1.01e-09 0.0014 1.013e-09 0 1.207e-09 0 1.21e-09 0.0014 1.213e-09 0 1.407e-09 0 1.41e-09 0.0014 1.413e-09 0 1.607e-09 0 1.61e-09 0.0014 1.613e-09 0 1.807e-09 0 1.81e-09 0.0014 1.813e-09 0 2.007e-09 0 2.01e-09 0.0014 2.013e-09 0 2.207e-09 0 2.21e-09 0.0014 2.213e-09 0 2.407e-09 0 2.41e-09 0.0014 2.413e-09 0 2.607e-09 0 2.61e-09 0.0014 2.613e-09 0 2.807e-09 0 2.81e-09 0.0014 2.813e-09 0 3.007e-09 0 3.01e-09 0.0014 3.013e-09 0 3.207e-09 0 3.21e-09 0.0014 3.213e-09 0 3.407e-09 0 3.41e-09 0.0014 3.413e-09 0 3.607e-09 0 3.61e-09 0.0014 3.613e-09 0 3.807e-09 0 3.81e-09 0.0014 3.813e-09 0 4.007e-09 0 4.01e-09 0.0014 4.013e-09 0 4.207e-09 0 4.21e-09 0.0014 4.213e-09 0 4.407e-09 0 4.41e-09 0.0014 4.413e-09 0 4.607e-09 0 4.61e-09 0.0014 4.613e-09 0 4.807e-09 0 4.81e-09 0.0014 4.813e-09 0 5.007e-09 0 5.01e-09 0.0014 5.013e-09 0 5.207e-09 0 5.21e-09 0.0014 5.213e-09 0 5.407e-09 0 5.41e-09 0.0014 5.413e-09 0 5.607e-09 0 5.61e-09 0.0014 5.613e-09 0 5.807e-09 0 5.81e-09 0.0014 5.813e-09 0 6.007e-09 0 6.01e-09 0.0014 6.013e-09 0 6.207e-09 0 6.21e-09 0.0014 6.213e-09 0 6.407e-09 0 6.41e-09 0.0014 6.413e-09 0 6.607e-09 0 6.61e-09 0.0014 6.613e-09 0 6.807e-09 0 6.81e-09 0.0014 6.813e-09 0 7.007e-09 0 7.01e-09 0.0014 7.013e-09 0 7.207e-09 0 7.21e-09 0.0014 7.213e-09 0 7.407e-09 0 7.41e-09 0.0014 7.413e-09 0 7.607e-09 0 7.61e-09 0.0014 7.613e-09 0 7.807e-09 0 7.81e-09 0.0014 7.813e-09 0 8.007e-09 0 8.01e-09 0.0014 8.013e-09 0 8.207e-09 0 8.21e-09 0.0014 8.213e-09 0 8.407e-09 0 8.41e-09 0.0014 8.413e-09 0 8.607e-09 0 8.61e-09 0.0014 8.613e-09 0 8.807e-09 0 8.81e-09 0.0014 8.813e-09 0 9.007e-09 0 9.01e-09 0.0014 9.013e-09 0 9.207e-09 0 9.21e-09 0.0014 9.213e-09 0 9.407e-09 0 9.41e-09 0.0014 9.413e-09 0 9.607e-09 0 9.61e-09 0.0014 9.613e-09 0 9.807e-09 0 9.81e-09 0.0014 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0014 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0014 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0014 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0014 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0014 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0014 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0014 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0014 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0014 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0014 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0014 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0014 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0014 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0014 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0014 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0014 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0014 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0014 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0014 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0014 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0014 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0014 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0014 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0014 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0014 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0014 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0014 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0014 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0014 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0014 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0014 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0014 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0014 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0014 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0014 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0014 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0014 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0014 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0014 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0014 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0014 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0014 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0014 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0014 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0014 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0014 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0014 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0014 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0014 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0014 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0014 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0014 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0014 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0014 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0014 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0014 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0014 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0014 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0014 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0014 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0014 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0014 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0014 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0014 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0014 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0014 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0014 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0014 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0014 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0014 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0014 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0014 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0014 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0014 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0014 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0014 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0014 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0014 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0014 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0014 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0014 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0014 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0014 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0014 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0014 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0014 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0014 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0014 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0014 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0014 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0014 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0014 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0014 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0014 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0014 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0014 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0014 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0014 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0014 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0014 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0014 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0014 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0014 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0014 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0014 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0014 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0014 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0014 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0014 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0014 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0014 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0014 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0014 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0014 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0014 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0014 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0014 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0014 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0014 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0014 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0014 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0014 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0014 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0014 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0014 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0014 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0014 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0014 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0014 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0014 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0014 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0014 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0014 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0014 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0014 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0014 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0014 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0014 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0014 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0014 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0014 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0014 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0014 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0014 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0014 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0014 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0014 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0014 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0014 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0014 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0014 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0014 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0014 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0014 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0014 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0014 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0014 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0014 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0014 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0014 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0014 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0014 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0014 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0014 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0014 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0014 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0014 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0014 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0014 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0014 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0014 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0014 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0014 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0014 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0014 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0014 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0014 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0014 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0014 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0014 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0014 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0014 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0014 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0014 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0014 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0014 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0014 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0014 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0014 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0014 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0014 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0014 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0014 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0014 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0014 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0014 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0014 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0014 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0014 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0014 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0014 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0014 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0014 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0014 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0014 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0014 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0014 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0014 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0014 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0014 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0014 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0014 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0014 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0014 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0014 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0014 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0014 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0014 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0014 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0014 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0014 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0014 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0014 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0014 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0014 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0014 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0014 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0014 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0014 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0014 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0014 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0014 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0014 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0014 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0014 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0014 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0014 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0014 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0014 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0014 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0014 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0014 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0014 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0014 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0014 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0014 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0014 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0014 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0014 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0014 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0014 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0014 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0014 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0014 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0014 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0014 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0014 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0014 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0014 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0014 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0014 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0014 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0014 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0014 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0014 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0014 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0014 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0014 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0014 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0014 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0014 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0014 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0014 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0014 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0014 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0014 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0014 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0014 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0014 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0014 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0014 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0014 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0014 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0014 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0014 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0014 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0014 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0014 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0014 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0014 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0014 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0014 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0014 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0014 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0014 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0014 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0014 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0014 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0014 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0014 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0014 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0014 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0014 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0014 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0014 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0014 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0014 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0014 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0014 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0014 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0014 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0014 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0014 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0014 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0014 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0014 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0014 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0014 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0014 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0014 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0014 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0014 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0014 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0014 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0014 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0014 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0014 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0014 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0014 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0014 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0014 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0014 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0014 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0014 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0014 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0014 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0014 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0014 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0014 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0014 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0014 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0014 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0014 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0014 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0014 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0014 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0014 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0014 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0014 7.9613e-08 0)
ID11|T 0 D11  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_DFF_IP1_12|1 IP1_1_OUT _DFF_IP1_12|A1  2.067833848e-12
L_DFF_IP1_12|2 _DFF_IP1_12|A1 _DFF_IP1_12|A2  4.135667696e-12
L_DFF_IP1_12|3 _DFF_IP1_12|A3 _DFF_IP1_12|A4  8.271335392e-12
L_DFF_IP1_12|T D11 _DFF_IP1_12|T1  2.067833848e-12
L_DFF_IP1_12|4 _DFF_IP1_12|T1 _DFF_IP1_12|T2  4.135667696e-12
L_DFF_IP1_12|5 _DFF_IP1_12|A4 _DFF_IP1_12|Q1  4.135667696e-12
L_DFF_IP1_12|6 _DFF_IP1_12|Q1 IP1_2_OUT  2.067833848e-12
ID12|T 0 D12  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_DFF_IP2_12|1 IP2_1_OUT _DFF_IP2_12|A1  2.067833848e-12
L_DFF_IP2_12|2 _DFF_IP2_12|A1 _DFF_IP2_12|A2  4.135667696e-12
L_DFF_IP2_12|3 _DFF_IP2_12|A3 _DFF_IP2_12|A4  8.271335392e-12
L_DFF_IP2_12|T D12 _DFF_IP2_12|T1  2.067833848e-12
L_DFF_IP2_12|4 _DFF_IP2_12|T1 _DFF_IP2_12|T2  4.135667696e-12
L_DFF_IP2_12|5 _DFF_IP2_12|A4 _DFF_IP2_12|Q1  4.135667696e-12
L_DFF_IP2_12|6 _DFF_IP2_12|Q1 IP2_2_OUT  2.067833848e-12
ID13|T 0 D13  PWL(0 0 7e-12 0 1e-11 0.0007 1.3e-11 0 2.07e-10 0 2.1e-10 0.0007 2.13e-10 0 4.07e-10 0 4.1e-10 0.0007 4.13e-10 0 6.07e-10 0 6.1e-10 0.0007 6.13e-10 0 8.07e-10 0 8.1e-10 0.0007 8.13e-10 0 1.007e-09 0 1.01e-09 0.0007 1.013e-09 0 1.207e-09 0 1.21e-09 0.0007 1.213e-09 0 1.407e-09 0 1.41e-09 0.0007 1.413e-09 0 1.607e-09 0 1.61e-09 0.0007 1.613e-09 0 1.807e-09 0 1.81e-09 0.0007 1.813e-09 0 2.007e-09 0 2.01e-09 0.0007 2.013e-09 0 2.207e-09 0 2.21e-09 0.0007 2.213e-09 0 2.407e-09 0 2.41e-09 0.0007 2.413e-09 0 2.607e-09 0 2.61e-09 0.0007 2.613e-09 0 2.807e-09 0 2.81e-09 0.0007 2.813e-09 0 3.007e-09 0 3.01e-09 0.0007 3.013e-09 0 3.207e-09 0 3.21e-09 0.0007 3.213e-09 0 3.407e-09 0 3.41e-09 0.0007 3.413e-09 0 3.607e-09 0 3.61e-09 0.0007 3.613e-09 0 3.807e-09 0 3.81e-09 0.0007 3.813e-09 0 4.007e-09 0 4.01e-09 0.0007 4.013e-09 0 4.207e-09 0 4.21e-09 0.0007 4.213e-09 0 4.407e-09 0 4.41e-09 0.0007 4.413e-09 0 4.607e-09 0 4.61e-09 0.0007 4.613e-09 0 4.807e-09 0 4.81e-09 0.0007 4.813e-09 0 5.007e-09 0 5.01e-09 0.0007 5.013e-09 0 5.207e-09 0 5.21e-09 0.0007 5.213e-09 0 5.407e-09 0 5.41e-09 0.0007 5.413e-09 0 5.607e-09 0 5.61e-09 0.0007 5.613e-09 0 5.807e-09 0 5.81e-09 0.0007 5.813e-09 0 6.007e-09 0 6.01e-09 0.0007 6.013e-09 0 6.207e-09 0 6.21e-09 0.0007 6.213e-09 0 6.407e-09 0 6.41e-09 0.0007 6.413e-09 0 6.607e-09 0 6.61e-09 0.0007 6.613e-09 0 6.807e-09 0 6.81e-09 0.0007 6.813e-09 0 7.007e-09 0 7.01e-09 0.0007 7.013e-09 0 7.207e-09 0 7.21e-09 0.0007 7.213e-09 0 7.407e-09 0 7.41e-09 0.0007 7.413e-09 0 7.607e-09 0 7.61e-09 0.0007 7.613e-09 0 7.807e-09 0 7.81e-09 0.0007 7.813e-09 0 8.007e-09 0 8.01e-09 0.0007 8.013e-09 0 8.207e-09 0 8.21e-09 0.0007 8.213e-09 0 8.407e-09 0 8.41e-09 0.0007 8.413e-09 0 8.607e-09 0 8.61e-09 0.0007 8.613e-09 0 8.807e-09 0 8.81e-09 0.0007 8.813e-09 0 9.007e-09 0 9.01e-09 0.0007 9.013e-09 0 9.207e-09 0 9.21e-09 0.0007 9.213e-09 0 9.407e-09 0 9.41e-09 0.0007 9.413e-09 0 9.607e-09 0 9.61e-09 0.0007 9.613e-09 0 9.807e-09 0 9.81e-09 0.0007 9.813e-09 0 1.0007e-08 0 1.001e-08 0.0007 1.0013e-08 0 1.0207e-08 0 1.021e-08 0.0007 1.0213e-08 0 1.0407e-08 0 1.041e-08 0.0007 1.0413e-08 0 1.0607e-08 0 1.061e-08 0.0007 1.0613e-08 0 1.0807e-08 0 1.081e-08 0.0007 1.0813e-08 0 1.1007e-08 0 1.101e-08 0.0007 1.1013e-08 0 1.1207e-08 0 1.121e-08 0.0007 1.1213e-08 0 1.1407e-08 0 1.141e-08 0.0007 1.1413e-08 0 1.1607e-08 0 1.161e-08 0.0007 1.1613e-08 0 1.1807e-08 0 1.181e-08 0.0007 1.1813e-08 0 1.2007e-08 0 1.201e-08 0.0007 1.2013e-08 0 1.2207e-08 0 1.221e-08 0.0007 1.2213e-08 0 1.2407e-08 0 1.241e-08 0.0007 1.2413e-08 0 1.2607e-08 0 1.261e-08 0.0007 1.2613e-08 0 1.2807e-08 0 1.281e-08 0.0007 1.2813e-08 0 1.3007e-08 0 1.301e-08 0.0007 1.3013e-08 0 1.3207e-08 0 1.321e-08 0.0007 1.3213e-08 0 1.3407e-08 0 1.341e-08 0.0007 1.3413e-08 0 1.3607e-08 0 1.361e-08 0.0007 1.3613e-08 0 1.3807e-08 0 1.381e-08 0.0007 1.3813e-08 0 1.4007e-08 0 1.401e-08 0.0007 1.4013e-08 0 1.4207e-08 0 1.421e-08 0.0007 1.4213e-08 0 1.4407e-08 0 1.441e-08 0.0007 1.4413e-08 0 1.4607e-08 0 1.461e-08 0.0007 1.4613e-08 0 1.4807e-08 0 1.481e-08 0.0007 1.4813e-08 0 1.5007e-08 0 1.501e-08 0.0007 1.5013e-08 0 1.5207e-08 0 1.521e-08 0.0007 1.5213e-08 0 1.5407e-08 0 1.541e-08 0.0007 1.5413e-08 0 1.5607e-08 0 1.561e-08 0.0007 1.5613e-08 0 1.5807e-08 0 1.581e-08 0.0007 1.5813e-08 0 1.6007e-08 0 1.601e-08 0.0007 1.6013e-08 0 1.6207e-08 0 1.621e-08 0.0007 1.6213e-08 0 1.6407e-08 0 1.641e-08 0.0007 1.6413e-08 0 1.6607e-08 0 1.661e-08 0.0007 1.6613e-08 0 1.6807e-08 0 1.681e-08 0.0007 1.6813e-08 0 1.7007e-08 0 1.701e-08 0.0007 1.7013e-08 0 1.7207e-08 0 1.721e-08 0.0007 1.7213e-08 0 1.7407e-08 0 1.741e-08 0.0007 1.7413e-08 0 1.7607e-08 0 1.761e-08 0.0007 1.7613e-08 0 1.7807e-08 0 1.781e-08 0.0007 1.7813e-08 0 1.8007e-08 0 1.801e-08 0.0007 1.8013e-08 0 1.8207e-08 0 1.821e-08 0.0007 1.8213e-08 0 1.8407e-08 0 1.841e-08 0.0007 1.8413e-08 0 1.8607e-08 0 1.861e-08 0.0007 1.8613e-08 0 1.8807e-08 0 1.881e-08 0.0007 1.8813e-08 0 1.9007e-08 0 1.901e-08 0.0007 1.9013e-08 0 1.9207e-08 0 1.921e-08 0.0007 1.9213e-08 0 1.9407e-08 0 1.941e-08 0.0007 1.9413e-08 0 1.9607e-08 0 1.961e-08 0.0007 1.9613e-08 0 1.9807e-08 0 1.981e-08 0.0007 1.9813e-08 0 2.0007e-08 0 2.001e-08 0.0007 2.0013e-08 0 2.0207e-08 0 2.021e-08 0.0007 2.0213e-08 0 2.0407e-08 0 2.041e-08 0.0007 2.0413e-08 0 2.0607e-08 0 2.061e-08 0.0007 2.0613e-08 0 2.0807e-08 0 2.081e-08 0.0007 2.0813e-08 0 2.1007e-08 0 2.101e-08 0.0007 2.1013e-08 0 2.1207e-08 0 2.121e-08 0.0007 2.1213e-08 0 2.1407e-08 0 2.141e-08 0.0007 2.1413e-08 0 2.1607e-08 0 2.161e-08 0.0007 2.1613e-08 0 2.1807e-08 0 2.181e-08 0.0007 2.1813e-08 0 2.2007e-08 0 2.201e-08 0.0007 2.2013e-08 0 2.2207e-08 0 2.221e-08 0.0007 2.2213e-08 0 2.2407e-08 0 2.241e-08 0.0007 2.2413e-08 0 2.2607e-08 0 2.261e-08 0.0007 2.2613e-08 0 2.2807e-08 0 2.281e-08 0.0007 2.2813e-08 0 2.3007e-08 0 2.301e-08 0.0007 2.3013e-08 0 2.3207e-08 0 2.321e-08 0.0007 2.3213e-08 0 2.3407e-08 0 2.341e-08 0.0007 2.3413e-08 0 2.3607e-08 0 2.361e-08 0.0007 2.3613e-08 0 2.3807e-08 0 2.381e-08 0.0007 2.3813e-08 0 2.4007e-08 0 2.401e-08 0.0007 2.4013e-08 0 2.4207e-08 0 2.421e-08 0.0007 2.4213e-08 0 2.4407e-08 0 2.441e-08 0.0007 2.4413e-08 0 2.4607e-08 0 2.461e-08 0.0007 2.4613e-08 0 2.4807e-08 0 2.481e-08 0.0007 2.4813e-08 0 2.5007e-08 0 2.501e-08 0.0007 2.5013e-08 0 2.5207e-08 0 2.521e-08 0.0007 2.5213e-08 0 2.5407e-08 0 2.541e-08 0.0007 2.5413e-08 0 2.5607e-08 0 2.561e-08 0.0007 2.5613e-08 0 2.5807e-08 0 2.581e-08 0.0007 2.5813e-08 0 2.6007e-08 0 2.601e-08 0.0007 2.6013e-08 0 2.6207e-08 0 2.621e-08 0.0007 2.6213e-08 0 2.6407e-08 0 2.641e-08 0.0007 2.6413e-08 0 2.6607e-08 0 2.661e-08 0.0007 2.6613e-08 0 2.6807e-08 0 2.681e-08 0.0007 2.6813e-08 0 2.7007e-08 0 2.701e-08 0.0007 2.7013e-08 0 2.7207e-08 0 2.721e-08 0.0007 2.7213e-08 0 2.7407e-08 0 2.741e-08 0.0007 2.7413e-08 0 2.7607e-08 0 2.761e-08 0.0007 2.7613e-08 0 2.7807e-08 0 2.781e-08 0.0007 2.7813e-08 0 2.8007e-08 0 2.801e-08 0.0007 2.8013e-08 0 2.8207e-08 0 2.821e-08 0.0007 2.8213e-08 0 2.8407e-08 0 2.841e-08 0.0007 2.8413e-08 0 2.8607e-08 0 2.861e-08 0.0007 2.8613e-08 0 2.8807e-08 0 2.881e-08 0.0007 2.8813e-08 0 2.9007e-08 0 2.901e-08 0.0007 2.9013e-08 0 2.9207e-08 0 2.921e-08 0.0007 2.9213e-08 0 2.9407e-08 0 2.941e-08 0.0007 2.9413e-08 0 2.9607e-08 0 2.961e-08 0.0007 2.9613e-08 0 2.9807e-08 0 2.981e-08 0.0007 2.9813e-08 0 3.0007e-08 0 3.001e-08 0.0007 3.0013e-08 0 3.0207e-08 0 3.021e-08 0.0007 3.0213e-08 0 3.0407e-08 0 3.041e-08 0.0007 3.0413e-08 0 3.0607e-08 0 3.061e-08 0.0007 3.0613e-08 0 3.0807e-08 0 3.081e-08 0.0007 3.0813e-08 0 3.1007e-08 0 3.101e-08 0.0007 3.1013e-08 0 3.1207e-08 0 3.121e-08 0.0007 3.1213e-08 0 3.1407e-08 0 3.141e-08 0.0007 3.1413e-08 0 3.1607e-08 0 3.161e-08 0.0007 3.1613e-08 0 3.1807e-08 0 3.181e-08 0.0007 3.1813e-08 0 3.2007e-08 0 3.201e-08 0.0007 3.2013e-08 0 3.2207e-08 0 3.221e-08 0.0007 3.2213e-08 0 3.2407e-08 0 3.241e-08 0.0007 3.2413e-08 0 3.2607e-08 0 3.261e-08 0.0007 3.2613e-08 0 3.2807e-08 0 3.281e-08 0.0007 3.2813e-08 0 3.3007e-08 0 3.301e-08 0.0007 3.3013e-08 0 3.3207e-08 0 3.321e-08 0.0007 3.3213e-08 0 3.3407e-08 0 3.341e-08 0.0007 3.3413e-08 0 3.3607e-08 0 3.361e-08 0.0007 3.3613e-08 0 3.3807e-08 0 3.381e-08 0.0007 3.3813e-08 0 3.4007e-08 0 3.401e-08 0.0007 3.4013e-08 0 3.4207e-08 0 3.421e-08 0.0007 3.4213e-08 0 3.4407e-08 0 3.441e-08 0.0007 3.4413e-08 0 3.4607e-08 0 3.461e-08 0.0007 3.4613e-08 0 3.4807e-08 0 3.481e-08 0.0007 3.4813e-08 0 3.5007e-08 0 3.501e-08 0.0007 3.5013e-08 0 3.5207e-08 0 3.521e-08 0.0007 3.5213e-08 0 3.5407e-08 0 3.541e-08 0.0007 3.5413e-08 0 3.5607e-08 0 3.561e-08 0.0007 3.5613e-08 0 3.5807e-08 0 3.581e-08 0.0007 3.5813e-08 0 3.6007e-08 0 3.601e-08 0.0007 3.6013e-08 0 3.6207e-08 0 3.621e-08 0.0007 3.6213e-08 0 3.6407e-08 0 3.641e-08 0.0007 3.6413e-08 0 3.6607e-08 0 3.661e-08 0.0007 3.6613e-08 0 3.6807e-08 0 3.681e-08 0.0007 3.6813e-08 0 3.7007e-08 0 3.701e-08 0.0007 3.7013e-08 0 3.7207e-08 0 3.721e-08 0.0007 3.7213e-08 0 3.7407e-08 0 3.741e-08 0.0007 3.7413e-08 0 3.7607e-08 0 3.761e-08 0.0007 3.7613e-08 0 3.7807e-08 0 3.781e-08 0.0007 3.7813e-08 0 3.8007e-08 0 3.801e-08 0.0007 3.8013e-08 0 3.8207e-08 0 3.821e-08 0.0007 3.8213e-08 0 3.8407e-08 0 3.841e-08 0.0007 3.8413e-08 0 3.8607e-08 0 3.861e-08 0.0007 3.8613e-08 0 3.8807e-08 0 3.881e-08 0.0007 3.8813e-08 0 3.9007e-08 0 3.901e-08 0.0007 3.9013e-08 0 3.9207e-08 0 3.921e-08 0.0007 3.9213e-08 0 3.9407e-08 0 3.941e-08 0.0007 3.9413e-08 0 3.9607e-08 0 3.961e-08 0.0007 3.9613e-08 0 3.9807e-08 0 3.981e-08 0.0007 3.9813e-08 0 4.0007e-08 0 4.001e-08 0.0007 4.0013e-08 0 4.0207e-08 0 4.021e-08 0.0007 4.0213e-08 0 4.0407e-08 0 4.041e-08 0.0007 4.0413e-08 0 4.0607e-08 0 4.061e-08 0.0007 4.0613e-08 0 4.0807e-08 0 4.081e-08 0.0007 4.0813e-08 0 4.1007e-08 0 4.101e-08 0.0007 4.1013e-08 0 4.1207e-08 0 4.121e-08 0.0007 4.1213e-08 0 4.1407e-08 0 4.141e-08 0.0007 4.1413e-08 0 4.1607e-08 0 4.161e-08 0.0007 4.1613e-08 0 4.1807e-08 0 4.181e-08 0.0007 4.1813e-08 0 4.2007e-08 0 4.201e-08 0.0007 4.2013e-08 0 4.2207e-08 0 4.221e-08 0.0007 4.2213e-08 0 4.2407e-08 0 4.241e-08 0.0007 4.2413e-08 0 4.2607e-08 0 4.261e-08 0.0007 4.2613e-08 0 4.2807e-08 0 4.281e-08 0.0007 4.2813e-08 0 4.3007e-08 0 4.301e-08 0.0007 4.3013e-08 0 4.3207e-08 0 4.321e-08 0.0007 4.3213e-08 0 4.3407e-08 0 4.341e-08 0.0007 4.3413e-08 0 4.3607e-08 0 4.361e-08 0.0007 4.3613e-08 0 4.3807e-08 0 4.381e-08 0.0007 4.3813e-08 0 4.4007e-08 0 4.401e-08 0.0007 4.4013e-08 0 4.4207e-08 0 4.421e-08 0.0007 4.4213e-08 0 4.4407e-08 0 4.441e-08 0.0007 4.4413e-08 0 4.4607e-08 0 4.461e-08 0.0007 4.4613e-08 0 4.4807e-08 0 4.481e-08 0.0007 4.4813e-08 0 4.5007e-08 0 4.501e-08 0.0007 4.5013e-08 0 4.5207e-08 0 4.521e-08 0.0007 4.5213e-08 0 4.5407e-08 0 4.541e-08 0.0007 4.5413e-08 0 4.5607e-08 0 4.561e-08 0.0007 4.5613e-08 0 4.5807e-08 0 4.581e-08 0.0007 4.5813e-08 0 4.6007e-08 0 4.601e-08 0.0007 4.6013e-08 0 4.6207e-08 0 4.621e-08 0.0007 4.6213e-08 0 4.6407e-08 0 4.641e-08 0.0007 4.6413e-08 0 4.6607e-08 0 4.661e-08 0.0007 4.6613e-08 0 4.6807e-08 0 4.681e-08 0.0007 4.6813e-08 0 4.7007e-08 0 4.701e-08 0.0007 4.7013e-08 0 4.7207e-08 0 4.721e-08 0.0007 4.7213e-08 0 4.7407e-08 0 4.741e-08 0.0007 4.7413e-08 0 4.7607e-08 0 4.761e-08 0.0007 4.7613e-08 0 4.7807e-08 0 4.781e-08 0.0007 4.7813e-08 0 4.8007e-08 0 4.801e-08 0.0007 4.8013e-08 0 4.8207e-08 0 4.821e-08 0.0007 4.8213e-08 0 4.8407e-08 0 4.841e-08 0.0007 4.8413e-08 0 4.8607e-08 0 4.861e-08 0.0007 4.8613e-08 0 4.8807e-08 0 4.881e-08 0.0007 4.8813e-08 0 4.9007e-08 0 4.901e-08 0.0007 4.9013e-08 0 4.9207e-08 0 4.921e-08 0.0007 4.9213e-08 0 4.9407e-08 0 4.941e-08 0.0007 4.9413e-08 0 4.9607e-08 0 4.961e-08 0.0007 4.9613e-08 0 4.9807e-08 0 4.981e-08 0.0007 4.9813e-08 0 5.0007e-08 0 5.001e-08 0.0007 5.0013e-08 0 5.0207e-08 0 5.021e-08 0.0007 5.0213e-08 0 5.0407e-08 0 5.041e-08 0.0007 5.0413e-08 0 5.0607e-08 0 5.061e-08 0.0007 5.0613e-08 0 5.0807e-08 0 5.081e-08 0.0007 5.0813e-08 0 5.1007e-08 0 5.101e-08 0.0007 5.1013e-08 0 5.1207e-08 0 5.121e-08 0.0007 5.1213e-08 0 5.1407e-08 0 5.141e-08 0.0007 5.1413e-08 0 5.1607e-08 0 5.161e-08 0.0007 5.1613e-08 0 5.1807e-08 0 5.181e-08 0.0007 5.1813e-08 0 5.2007e-08 0 5.201e-08 0.0007 5.2013e-08 0 5.2207e-08 0 5.221e-08 0.0007 5.2213e-08 0 5.2407e-08 0 5.241e-08 0.0007 5.2413e-08 0 5.2607e-08 0 5.261e-08 0.0007 5.2613e-08 0 5.2807e-08 0 5.281e-08 0.0007 5.2813e-08 0 5.3007e-08 0 5.301e-08 0.0007 5.3013e-08 0 5.3207e-08 0 5.321e-08 0.0007 5.3213e-08 0 5.3407e-08 0 5.341e-08 0.0007 5.3413e-08 0 5.3607e-08 0 5.361e-08 0.0007 5.3613e-08 0 5.3807e-08 0 5.381e-08 0.0007 5.3813e-08 0 5.4007e-08 0 5.401e-08 0.0007 5.4013e-08 0 5.4207e-08 0 5.421e-08 0.0007 5.4213e-08 0 5.4407e-08 0 5.441e-08 0.0007 5.4413e-08 0 5.4607e-08 0 5.461e-08 0.0007 5.4613e-08 0 5.4807e-08 0 5.481e-08 0.0007 5.4813e-08 0 5.5007e-08 0 5.501e-08 0.0007 5.5013e-08 0 5.5207e-08 0 5.521e-08 0.0007 5.5213e-08 0 5.5407e-08 0 5.541e-08 0.0007 5.5413e-08 0 5.5607e-08 0 5.561e-08 0.0007 5.5613e-08 0 5.5807e-08 0 5.581e-08 0.0007 5.5813e-08 0 5.6007e-08 0 5.601e-08 0.0007 5.6013e-08 0 5.6207e-08 0 5.621e-08 0.0007 5.6213e-08 0 5.6407e-08 0 5.641e-08 0.0007 5.6413e-08 0 5.6607e-08 0 5.661e-08 0.0007 5.6613e-08 0 5.6807e-08 0 5.681e-08 0.0007 5.6813e-08 0 5.7007e-08 0 5.701e-08 0.0007 5.7013e-08 0 5.7207e-08 0 5.721e-08 0.0007 5.7213e-08 0 5.7407e-08 0 5.741e-08 0.0007 5.7413e-08 0 5.7607e-08 0 5.761e-08 0.0007 5.7613e-08 0 5.7807e-08 0 5.781e-08 0.0007 5.7813e-08 0 5.8007e-08 0 5.801e-08 0.0007 5.8013e-08 0 5.8207e-08 0 5.821e-08 0.0007 5.8213e-08 0 5.8407e-08 0 5.841e-08 0.0007 5.8413e-08 0 5.8607e-08 0 5.861e-08 0.0007 5.8613e-08 0 5.8807e-08 0 5.881e-08 0.0007 5.8813e-08 0 5.9007e-08 0 5.901e-08 0.0007 5.9013e-08 0 5.9207e-08 0 5.921e-08 0.0007 5.9213e-08 0 5.9407e-08 0 5.941e-08 0.0007 5.9413e-08 0 5.9607e-08 0 5.961e-08 0.0007 5.9613e-08 0 5.9807e-08 0 5.981e-08 0.0007 5.9813e-08 0 6.0007e-08 0 6.001e-08 0.0007 6.0013e-08 0 6.0207e-08 0 6.021e-08 0.0007 6.0213e-08 0 6.0407e-08 0 6.041e-08 0.0007 6.0413e-08 0 6.0607e-08 0 6.061e-08 0.0007 6.0613e-08 0 6.0807e-08 0 6.081e-08 0.0007 6.0813e-08 0 6.1007e-08 0 6.101e-08 0.0007 6.1013e-08 0 6.1207e-08 0 6.121e-08 0.0007 6.1213e-08 0 6.1407e-08 0 6.141e-08 0.0007 6.1413e-08 0 6.1607e-08 0 6.161e-08 0.0007 6.1613e-08 0 6.1807e-08 0 6.181e-08 0.0007 6.1813e-08 0 6.2007e-08 0 6.201e-08 0.0007 6.2013e-08 0 6.2207e-08 0 6.221e-08 0.0007 6.2213e-08 0 6.2407e-08 0 6.241e-08 0.0007 6.2413e-08 0 6.2607e-08 0 6.261e-08 0.0007 6.2613e-08 0 6.2807e-08 0 6.281e-08 0.0007 6.2813e-08 0 6.3007e-08 0 6.301e-08 0.0007 6.3013e-08 0 6.3207e-08 0 6.321e-08 0.0007 6.3213e-08 0 6.3407e-08 0 6.341e-08 0.0007 6.3413e-08 0 6.3607e-08 0 6.361e-08 0.0007 6.3613e-08 0 6.3807e-08 0 6.381e-08 0.0007 6.3813e-08 0 6.4007e-08 0 6.401e-08 0.0007 6.4013e-08 0 6.4207e-08 0 6.421e-08 0.0007 6.4213e-08 0 6.4407e-08 0 6.441e-08 0.0007 6.4413e-08 0 6.4607e-08 0 6.461e-08 0.0007 6.4613e-08 0 6.4807e-08 0 6.481e-08 0.0007 6.4813e-08 0 6.5007e-08 0 6.501e-08 0.0007 6.5013e-08 0 6.5207e-08 0 6.521e-08 0.0007 6.5213e-08 0 6.5407e-08 0 6.541e-08 0.0007 6.5413e-08 0 6.5607e-08 0 6.561e-08 0.0007 6.5613e-08 0 6.5807e-08 0 6.581e-08 0.0007 6.5813e-08 0 6.6007e-08 0 6.601e-08 0.0007 6.6013e-08 0 6.6207e-08 0 6.621e-08 0.0007 6.6213e-08 0 6.6407e-08 0 6.641e-08 0.0007 6.6413e-08 0 6.6607e-08 0 6.661e-08 0.0007 6.6613e-08 0 6.6807e-08 0 6.681e-08 0.0007 6.6813e-08 0 6.7007e-08 0 6.701e-08 0.0007 6.7013e-08 0 6.7207e-08 0 6.721e-08 0.0007 6.7213e-08 0 6.7407e-08 0 6.741e-08 0.0007 6.7413e-08 0 6.7607e-08 0 6.761e-08 0.0007 6.7613e-08 0 6.7807e-08 0 6.781e-08 0.0007 6.7813e-08 0 6.8007e-08 0 6.801e-08 0.0007 6.8013e-08 0 6.8207e-08 0 6.821e-08 0.0007 6.8213e-08 0 6.8407e-08 0 6.841e-08 0.0007 6.8413e-08 0 6.8607e-08 0 6.861e-08 0.0007 6.8613e-08 0 6.8807e-08 0 6.881e-08 0.0007 6.8813e-08 0 6.9007e-08 0 6.901e-08 0.0007 6.9013e-08 0 6.9207e-08 0 6.921e-08 0.0007 6.9213e-08 0 6.9407e-08 0 6.941e-08 0.0007 6.9413e-08 0 6.9607e-08 0 6.961e-08 0.0007 6.9613e-08 0 6.9807e-08 0 6.981e-08 0.0007 6.9813e-08 0 7.0007e-08 0 7.001e-08 0.0007 7.0013e-08 0 7.0207e-08 0 7.021e-08 0.0007 7.0213e-08 0 7.0407e-08 0 7.041e-08 0.0007 7.0413e-08 0 7.0607e-08 0 7.061e-08 0.0007 7.0613e-08 0 7.0807e-08 0 7.081e-08 0.0007 7.0813e-08 0 7.1007e-08 0 7.101e-08 0.0007 7.1013e-08 0 7.1207e-08 0 7.121e-08 0.0007 7.1213e-08 0 7.1407e-08 0 7.141e-08 0.0007 7.1413e-08 0 7.1607e-08 0 7.161e-08 0.0007 7.1613e-08 0 7.1807e-08 0 7.181e-08 0.0007 7.1813e-08 0 7.2007e-08 0 7.201e-08 0.0007 7.2013e-08 0 7.2207e-08 0 7.221e-08 0.0007 7.2213e-08 0 7.2407e-08 0 7.241e-08 0.0007 7.2413e-08 0 7.2607e-08 0 7.261e-08 0.0007 7.2613e-08 0 7.2807e-08 0 7.281e-08 0.0007 7.2813e-08 0 7.3007e-08 0 7.301e-08 0.0007 7.3013e-08 0 7.3207e-08 0 7.321e-08 0.0007 7.3213e-08 0 7.3407e-08 0 7.341e-08 0.0007 7.3413e-08 0 7.3607e-08 0 7.361e-08 0.0007 7.3613e-08 0 7.3807e-08 0 7.381e-08 0.0007 7.3813e-08 0 7.4007e-08 0 7.401e-08 0.0007 7.4013e-08 0 7.4207e-08 0 7.421e-08 0.0007 7.4213e-08 0 7.4407e-08 0 7.441e-08 0.0007 7.4413e-08 0 7.4607e-08 0 7.461e-08 0.0007 7.4613e-08 0 7.4807e-08 0 7.481e-08 0.0007 7.4813e-08 0 7.5007e-08 0 7.501e-08 0.0007 7.5013e-08 0 7.5207e-08 0 7.521e-08 0.0007 7.5213e-08 0 7.5407e-08 0 7.541e-08 0.0007 7.5413e-08 0 7.5607e-08 0 7.561e-08 0.0007 7.5613e-08 0 7.5807e-08 0 7.581e-08 0.0007 7.5813e-08 0 7.6007e-08 0 7.601e-08 0.0007 7.6013e-08 0 7.6207e-08 0 7.621e-08 0.0007 7.6213e-08 0 7.6407e-08 0 7.641e-08 0.0007 7.6413e-08 0 7.6607e-08 0 7.661e-08 0.0007 7.6613e-08 0 7.6807e-08 0 7.681e-08 0.0007 7.6813e-08 0 7.7007e-08 0 7.701e-08 0.0007 7.7013e-08 0 7.7207e-08 0 7.721e-08 0.0007 7.7213e-08 0 7.7407e-08 0 7.741e-08 0.0007 7.7413e-08 0 7.7607e-08 0 7.761e-08 0.0007 7.7613e-08 0 7.7807e-08 0 7.781e-08 0.0007 7.7813e-08 0 7.8007e-08 0 7.801e-08 0.0007 7.8013e-08 0 7.8207e-08 0 7.821e-08 0.0007 7.8213e-08 0 7.8407e-08 0 7.841e-08 0.0007 7.8413e-08 0 7.8607e-08 0 7.861e-08 0.0007 7.8613e-08 0 7.8807e-08 0 7.881e-08 0.0007 7.8813e-08 0 7.9007e-08 0 7.901e-08 0.0007 7.9013e-08 0 7.9207e-08 0 7.921e-08 0.0007 7.9213e-08 0 7.9407e-08 0 7.941e-08 0.0007 7.9413e-08 0 7.9607e-08 0 7.961e-08 0.0007 7.9613e-08 0)
L_DFF_IP3_12|1 IP3_1_OUT _DFF_IP3_12|A1  2.067833848e-12
L_DFF_IP3_12|2 _DFF_IP3_12|A1 _DFF_IP3_12|A2  4.135667696e-12
L_DFF_IP3_12|3 _DFF_IP3_12|A3 _DFF_IP3_12|A4  8.271335392e-12
L_DFF_IP3_12|T D13 _DFF_IP3_12|T1  2.067833848e-12
L_DFF_IP3_12|4 _DFF_IP3_12|T1 _DFF_IP3_12|T2  4.135667696e-12
L_DFF_IP3_12|5 _DFF_IP3_12|A4 _DFF_IP3_12|Q1  4.135667696e-12
L_DFF_IP3_12|6 _DFF_IP3_12|Q1 IP3_2_OUT  2.067833848e-12
IT12|T 0 T12  PWL(0 0 2e-12 0 5e-12 0.0007 8e-12 0 2.02e-10 0 2.05e-10 0.0007 2.08e-10 0 4.02e-10 0 4.05e-10 0.0007 4.08e-10 0 6.02e-10 0 6.05e-10 0.0007 6.08e-10 0 8.02e-10 0 8.05e-10 0.0007 8.08e-10 0 1.002e-09 0 1.005e-09 0.0007 1.008e-09 0 1.202e-09 0 1.205e-09 0.0007 1.208e-09 0 1.402e-09 0 1.405e-09 0.0007 1.408e-09 0 1.602e-09 0 1.605e-09 0.0007 1.608e-09 0 1.802e-09 0 1.805e-09 0.0007 1.808e-09 0 2.002e-09 0 2.005e-09 0.0007 2.008e-09 0 2.202e-09 0 2.205e-09 0.0007 2.208e-09 0 2.402e-09 0 2.405e-09 0.0007 2.408e-09 0 2.602e-09 0 2.605e-09 0.0007 2.608e-09 0 2.802e-09 0 2.805e-09 0.0007 2.808e-09 0 3.002e-09 0 3.005e-09 0.0007 3.008e-09 0 3.202e-09 0 3.205e-09 0.0007 3.208e-09 0 3.402e-09 0 3.405e-09 0.0007 3.408e-09 0 3.602e-09 0 3.605e-09 0.0007 3.608e-09 0 3.802e-09 0 3.805e-09 0.0007 3.808e-09 0 4.002e-09 0 4.005e-09 0.0007 4.008e-09 0 4.202e-09 0 4.205e-09 0.0007 4.208e-09 0 4.402e-09 0 4.405e-09 0.0007 4.408e-09 0 4.602e-09 0 4.605e-09 0.0007 4.608e-09 0 4.802e-09 0 4.805e-09 0.0007 4.808e-09 0 5.002e-09 0 5.005e-09 0.0007 5.008e-09 0 5.202e-09 0 5.205e-09 0.0007 5.208e-09 0 5.402e-09 0 5.405e-09 0.0007 5.408e-09 0 5.602e-09 0 5.605e-09 0.0007 5.608e-09 0 5.802e-09 0 5.805e-09 0.0007 5.808e-09 0 6.002e-09 0 6.005e-09 0.0007 6.008e-09 0 6.202e-09 0 6.205e-09 0.0007 6.208e-09 0 6.402e-09 0 6.405e-09 0.0007 6.408e-09 0 6.602e-09 0 6.605e-09 0.0007 6.608e-09 0 6.802e-09 0 6.805e-09 0.0007 6.808e-09 0 7.002e-09 0 7.005e-09 0.0007 7.008e-09 0 7.202e-09 0 7.205e-09 0.0007 7.208e-09 0 7.402e-09 0 7.405e-09 0.0007 7.408e-09 0 7.602e-09 0 7.605e-09 0.0007 7.608e-09 0 7.802e-09 0 7.805e-09 0.0007 7.808e-09 0 8.002e-09 0 8.005e-09 0.0007 8.008e-09 0 8.202e-09 0 8.205e-09 0.0007 8.208e-09 0 8.402e-09 0 8.405e-09 0.0007 8.408e-09 0 8.602e-09 0 8.605e-09 0.0007 8.608e-09 0 8.802e-09 0 8.805e-09 0.0007 8.808e-09 0 9.002e-09 0 9.005e-09 0.0007 9.008e-09 0 9.202e-09 0 9.205e-09 0.0007 9.208e-09 0 9.402e-09 0 9.405e-09 0.0007 9.408e-09 0 9.602e-09 0 9.605e-09 0.0007 9.608e-09 0 9.802e-09 0 9.805e-09 0.0007 9.808e-09 0 1.0002e-08 0 1.0005e-08 0.0007 1.0008e-08 0 1.0202e-08 0 1.0205e-08 0.0007 1.0208e-08 0 1.0402e-08 0 1.0405e-08 0.0007 1.0408e-08 0 1.0602e-08 0 1.0605e-08 0.0007 1.0608e-08 0 1.0802e-08 0 1.0805e-08 0.0007 1.0808e-08 0 1.1002e-08 0 1.1005e-08 0.0007 1.1008e-08 0 1.1202e-08 0 1.1205e-08 0.0007 1.1208e-08 0 1.1402e-08 0 1.1405e-08 0.0007 1.1408e-08 0 1.1602e-08 0 1.1605e-08 0.0007 1.1608e-08 0 1.1802e-08 0 1.1805e-08 0.0007 1.1808e-08 0 1.2002e-08 0 1.2005e-08 0.0007 1.2008e-08 0 1.2202e-08 0 1.2205e-08 0.0007 1.2208e-08 0 1.2402e-08 0 1.2405e-08 0.0007 1.2408e-08 0 1.2602e-08 0 1.2605e-08 0.0007 1.2608e-08 0 1.2802e-08 0 1.2805e-08 0.0007 1.2808e-08 0 1.3002e-08 0 1.3005e-08 0.0007 1.3008e-08 0 1.3202e-08 0 1.3205e-08 0.0007 1.3208e-08 0 1.3402e-08 0 1.3405e-08 0.0007 1.3408e-08 0 1.3602e-08 0 1.3605e-08 0.0007 1.3608e-08 0 1.3802e-08 0 1.3805e-08 0.0007 1.3808e-08 0 1.4002e-08 0 1.4005e-08 0.0007 1.4008e-08 0 1.4202e-08 0 1.4205e-08 0.0007 1.4208e-08 0 1.4402e-08 0 1.4405e-08 0.0007 1.4408e-08 0 1.4602e-08 0 1.4605e-08 0.0007 1.4608e-08 0 1.4802e-08 0 1.4805e-08 0.0007 1.4808e-08 0 1.5002e-08 0 1.5005e-08 0.0007 1.5008e-08 0 1.5202e-08 0 1.5205e-08 0.0007 1.5208e-08 0 1.5402e-08 0 1.5405e-08 0.0007 1.5408e-08 0 1.5602e-08 0 1.5605e-08 0.0007 1.5608e-08 0 1.5802e-08 0 1.5805e-08 0.0007 1.5808e-08 0 1.6002e-08 0 1.6005e-08 0.0007 1.6008e-08 0 1.6202e-08 0 1.6205e-08 0.0007 1.6208e-08 0 1.6402e-08 0 1.6405e-08 0.0007 1.6408e-08 0 1.6602e-08 0 1.6605e-08 0.0007 1.6608e-08 0 1.6802e-08 0 1.6805e-08 0.0007 1.6808e-08 0 1.7002e-08 0 1.7005e-08 0.0007 1.7008e-08 0 1.7202e-08 0 1.7205e-08 0.0007 1.7208e-08 0 1.7402e-08 0 1.7405e-08 0.0007 1.7408e-08 0 1.7602e-08 0 1.7605e-08 0.0007 1.7608e-08 0 1.7802e-08 0 1.7805e-08 0.0007 1.7808e-08 0 1.8002e-08 0 1.8005e-08 0.0007 1.8008e-08 0 1.8202e-08 0 1.8205e-08 0.0007 1.8208e-08 0 1.8402e-08 0 1.8405e-08 0.0007 1.8408e-08 0 1.8602e-08 0 1.8605e-08 0.0007 1.8608e-08 0 1.8802e-08 0 1.8805e-08 0.0007 1.8808e-08 0 1.9002e-08 0 1.9005e-08 0.0007 1.9008e-08 0 1.9202e-08 0 1.9205e-08 0.0007 1.9208e-08 0 1.9402e-08 0 1.9405e-08 0.0007 1.9408e-08 0 1.9602e-08 0 1.9605e-08 0.0007 1.9608e-08 0 1.9802e-08 0 1.9805e-08 0.0007 1.9808e-08 0 2.0002e-08 0 2.0005e-08 0.0007 2.0008e-08 0 2.0202e-08 0 2.0205e-08 0.0007 2.0208e-08 0 2.0402e-08 0 2.0405e-08 0.0007 2.0408e-08 0 2.0602e-08 0 2.0605e-08 0.0007 2.0608e-08 0 2.0802e-08 0 2.0805e-08 0.0007 2.0808e-08 0 2.1002e-08 0 2.1005e-08 0.0007 2.1008e-08 0 2.1202e-08 0 2.1205e-08 0.0007 2.1208e-08 0 2.1402e-08 0 2.1405e-08 0.0007 2.1408e-08 0 2.1602e-08 0 2.1605e-08 0.0007 2.1608e-08 0 2.1802e-08 0 2.1805e-08 0.0007 2.1808e-08 0 2.2002e-08 0 2.2005e-08 0.0007 2.2008e-08 0 2.2202e-08 0 2.2205e-08 0.0007 2.2208e-08 0 2.2402e-08 0 2.2405e-08 0.0007 2.2408e-08 0 2.2602e-08 0 2.2605e-08 0.0007 2.2608e-08 0 2.2802e-08 0 2.2805e-08 0.0007 2.2808e-08 0 2.3002e-08 0 2.3005e-08 0.0007 2.3008e-08 0 2.3202e-08 0 2.3205e-08 0.0007 2.3208e-08 0 2.3402e-08 0 2.3405e-08 0.0007 2.3408e-08 0 2.3602e-08 0 2.3605e-08 0.0007 2.3608e-08 0 2.3802e-08 0 2.3805e-08 0.0007 2.3808e-08 0 2.4002e-08 0 2.4005e-08 0.0007 2.4008e-08 0 2.4202e-08 0 2.4205e-08 0.0007 2.4208e-08 0 2.4402e-08 0 2.4405e-08 0.0007 2.4408e-08 0 2.4602e-08 0 2.4605e-08 0.0007 2.4608e-08 0 2.4802e-08 0 2.4805e-08 0.0007 2.4808e-08 0 2.5002e-08 0 2.5005e-08 0.0007 2.5008e-08 0 2.5202e-08 0 2.5205e-08 0.0007 2.5208e-08 0 2.5402e-08 0 2.5405e-08 0.0007 2.5408e-08 0 2.5602e-08 0 2.5605e-08 0.0007 2.5608e-08 0 2.5802e-08 0 2.5805e-08 0.0007 2.5808e-08 0 2.6002e-08 0 2.6005e-08 0.0007 2.6008e-08 0 2.6202e-08 0 2.6205e-08 0.0007 2.6208e-08 0 2.6402e-08 0 2.6405e-08 0.0007 2.6408e-08 0 2.6602e-08 0 2.6605e-08 0.0007 2.6608e-08 0 2.6802e-08 0 2.6805e-08 0.0007 2.6808e-08 0 2.7002e-08 0 2.7005e-08 0.0007 2.7008e-08 0 2.7202e-08 0 2.7205e-08 0.0007 2.7208e-08 0 2.7402e-08 0 2.7405e-08 0.0007 2.7408e-08 0 2.7602e-08 0 2.7605e-08 0.0007 2.7608e-08 0 2.7802e-08 0 2.7805e-08 0.0007 2.7808e-08 0 2.8002e-08 0 2.8005e-08 0.0007 2.8008e-08 0 2.8202e-08 0 2.8205e-08 0.0007 2.8208e-08 0 2.8402e-08 0 2.8405e-08 0.0007 2.8408e-08 0 2.8602e-08 0 2.8605e-08 0.0007 2.8608e-08 0 2.8802e-08 0 2.8805e-08 0.0007 2.8808e-08 0 2.9002e-08 0 2.9005e-08 0.0007 2.9008e-08 0 2.9202e-08 0 2.9205e-08 0.0007 2.9208e-08 0 2.9402e-08 0 2.9405e-08 0.0007 2.9408e-08 0 2.9602e-08 0 2.9605e-08 0.0007 2.9608e-08 0 2.9802e-08 0 2.9805e-08 0.0007 2.9808e-08 0 3.0002e-08 0 3.0005e-08 0.0007 3.0008e-08 0 3.0202e-08 0 3.0205e-08 0.0007 3.0208e-08 0 3.0402e-08 0 3.0405e-08 0.0007 3.0408e-08 0 3.0602e-08 0 3.0605e-08 0.0007 3.0608e-08 0 3.0802e-08 0 3.0805e-08 0.0007 3.0808e-08 0 3.1002e-08 0 3.1005e-08 0.0007 3.1008e-08 0 3.1202e-08 0 3.1205e-08 0.0007 3.1208e-08 0 3.1402e-08 0 3.1405e-08 0.0007 3.1408e-08 0 3.1602e-08 0 3.1605e-08 0.0007 3.1608e-08 0 3.1802e-08 0 3.1805e-08 0.0007 3.1808e-08 0 3.2002e-08 0 3.2005e-08 0.0007 3.2008e-08 0 3.2202e-08 0 3.2205e-08 0.0007 3.2208e-08 0 3.2402e-08 0 3.2405e-08 0.0007 3.2408e-08 0 3.2602e-08 0 3.2605e-08 0.0007 3.2608e-08 0 3.2802e-08 0 3.2805e-08 0.0007 3.2808e-08 0 3.3002e-08 0 3.3005e-08 0.0007 3.3008e-08 0 3.3202e-08 0 3.3205e-08 0.0007 3.3208e-08 0 3.3402e-08 0 3.3405e-08 0.0007 3.3408e-08 0 3.3602e-08 0 3.3605e-08 0.0007 3.3608e-08 0 3.3802e-08 0 3.3805e-08 0.0007 3.3808e-08 0 3.4002e-08 0 3.4005e-08 0.0007 3.4008e-08 0 3.4202e-08 0 3.4205e-08 0.0007 3.4208e-08 0 3.4402e-08 0 3.4405e-08 0.0007 3.4408e-08 0 3.4602e-08 0 3.4605e-08 0.0007 3.4608e-08 0 3.4802e-08 0 3.4805e-08 0.0007 3.4808e-08 0 3.5002e-08 0 3.5005e-08 0.0007 3.5008e-08 0 3.5202e-08 0 3.5205e-08 0.0007 3.5208e-08 0 3.5402e-08 0 3.5405e-08 0.0007 3.5408e-08 0 3.5602e-08 0 3.5605e-08 0.0007 3.5608e-08 0 3.5802e-08 0 3.5805e-08 0.0007 3.5808e-08 0 3.6002e-08 0 3.6005e-08 0.0007 3.6008e-08 0 3.6202e-08 0 3.6205e-08 0.0007 3.6208e-08 0 3.6402e-08 0 3.6405e-08 0.0007 3.6408e-08 0 3.6602e-08 0 3.6605e-08 0.0007 3.6608e-08 0 3.6802e-08 0 3.6805e-08 0.0007 3.6808e-08 0 3.7002e-08 0 3.7005e-08 0.0007 3.7008e-08 0 3.7202e-08 0 3.7205e-08 0.0007 3.7208e-08 0 3.7402e-08 0 3.7405e-08 0.0007 3.7408e-08 0 3.7602e-08 0 3.7605e-08 0.0007 3.7608e-08 0 3.7802e-08 0 3.7805e-08 0.0007 3.7808e-08 0 3.8002e-08 0 3.8005e-08 0.0007 3.8008e-08 0 3.8202e-08 0 3.8205e-08 0.0007 3.8208e-08 0 3.8402e-08 0 3.8405e-08 0.0007 3.8408e-08 0 3.8602e-08 0 3.8605e-08 0.0007 3.8608e-08 0 3.8802e-08 0 3.8805e-08 0.0007 3.8808e-08 0 3.9002e-08 0 3.9005e-08 0.0007 3.9008e-08 0 3.9202e-08 0 3.9205e-08 0.0007 3.9208e-08 0 3.9402e-08 0 3.9405e-08 0.0007 3.9408e-08 0 3.9602e-08 0 3.9605e-08 0.0007 3.9608e-08 0 3.9802e-08 0 3.9805e-08 0.0007 3.9808e-08 0 4.0002e-08 0 4.0005e-08 0.0007 4.0008e-08 0 4.0202e-08 0 4.0205e-08 0.0007 4.0208e-08 0 4.0402e-08 0 4.0405e-08 0.0007 4.0408e-08 0 4.0602e-08 0 4.0605e-08 0.0007 4.0608e-08 0 4.0802e-08 0 4.0805e-08 0.0007 4.0808e-08 0 4.1002e-08 0 4.1005e-08 0.0007 4.1008e-08 0 4.1202e-08 0 4.1205e-08 0.0007 4.1208e-08 0 4.1402e-08 0 4.1405e-08 0.0007 4.1408e-08 0 4.1602e-08 0 4.1605e-08 0.0007 4.1608e-08 0 4.1802e-08 0 4.1805e-08 0.0007 4.1808e-08 0 4.2002e-08 0 4.2005e-08 0.0007 4.2008e-08 0 4.2202e-08 0 4.2205e-08 0.0007 4.2208e-08 0 4.2402e-08 0 4.2405e-08 0.0007 4.2408e-08 0 4.2602e-08 0 4.2605e-08 0.0007 4.2608e-08 0 4.2802e-08 0 4.2805e-08 0.0007 4.2808e-08 0 4.3002e-08 0 4.3005e-08 0.0007 4.3008e-08 0 4.3202e-08 0 4.3205e-08 0.0007 4.3208e-08 0 4.3402e-08 0 4.3405e-08 0.0007 4.3408e-08 0 4.3602e-08 0 4.3605e-08 0.0007 4.3608e-08 0 4.3802e-08 0 4.3805e-08 0.0007 4.3808e-08 0 4.4002e-08 0 4.4005e-08 0.0007 4.4008e-08 0 4.4202e-08 0 4.4205e-08 0.0007 4.4208e-08 0 4.4402e-08 0 4.4405e-08 0.0007 4.4408e-08 0 4.4602e-08 0 4.4605e-08 0.0007 4.4608e-08 0 4.4802e-08 0 4.4805e-08 0.0007 4.4808e-08 0 4.5002e-08 0 4.5005e-08 0.0007 4.5008e-08 0 4.5202e-08 0 4.5205e-08 0.0007 4.5208e-08 0 4.5402e-08 0 4.5405e-08 0.0007 4.5408e-08 0 4.5602e-08 0 4.5605e-08 0.0007 4.5608e-08 0 4.5802e-08 0 4.5805e-08 0.0007 4.5808e-08 0 4.6002e-08 0 4.6005e-08 0.0007 4.6008e-08 0 4.6202e-08 0 4.6205e-08 0.0007 4.6208e-08 0 4.6402e-08 0 4.6405e-08 0.0007 4.6408e-08 0 4.6602e-08 0 4.6605e-08 0.0007 4.6608e-08 0 4.6802e-08 0 4.6805e-08 0.0007 4.6808e-08 0 4.7002e-08 0 4.7005e-08 0.0007 4.7008e-08 0 4.7202e-08 0 4.7205e-08 0.0007 4.7208e-08 0 4.7402e-08 0 4.7405e-08 0.0007 4.7408e-08 0 4.7602e-08 0 4.7605e-08 0.0007 4.7608e-08 0 4.7802e-08 0 4.7805e-08 0.0007 4.7808e-08 0 4.8002e-08 0 4.8005e-08 0.0007 4.8008e-08 0 4.8202e-08 0 4.8205e-08 0.0007 4.8208e-08 0 4.8402e-08 0 4.8405e-08 0.0007 4.8408e-08 0 4.8602e-08 0 4.8605e-08 0.0007 4.8608e-08 0 4.8802e-08 0 4.8805e-08 0.0007 4.8808e-08 0 4.9002e-08 0 4.9005e-08 0.0007 4.9008e-08 0 4.9202e-08 0 4.9205e-08 0.0007 4.9208e-08 0 4.9402e-08 0 4.9405e-08 0.0007 4.9408e-08 0 4.9602e-08 0 4.9605e-08 0.0007 4.9608e-08 0 4.9802e-08 0 4.9805e-08 0.0007 4.9808e-08 0 5.0002e-08 0 5.0005e-08 0.0007 5.0008e-08 0 5.0202e-08 0 5.0205e-08 0.0007 5.0208e-08 0 5.0402e-08 0 5.0405e-08 0.0007 5.0408e-08 0 5.0602e-08 0 5.0605e-08 0.0007 5.0608e-08 0 5.0802e-08 0 5.0805e-08 0.0007 5.0808e-08 0 5.1002e-08 0 5.1005e-08 0.0007 5.1008e-08 0 5.1202e-08 0 5.1205e-08 0.0007 5.1208e-08 0 5.1402e-08 0 5.1405e-08 0.0007 5.1408e-08 0 5.1602e-08 0 5.1605e-08 0.0007 5.1608e-08 0 5.1802e-08 0 5.1805e-08 0.0007 5.1808e-08 0 5.2002e-08 0 5.2005e-08 0.0007 5.2008e-08 0 5.2202e-08 0 5.2205e-08 0.0007 5.2208e-08 0 5.2402e-08 0 5.2405e-08 0.0007 5.2408e-08 0 5.2602e-08 0 5.2605e-08 0.0007 5.2608e-08 0 5.2802e-08 0 5.2805e-08 0.0007 5.2808e-08 0 5.3002e-08 0 5.3005e-08 0.0007 5.3008e-08 0 5.3202e-08 0 5.3205e-08 0.0007 5.3208e-08 0 5.3402e-08 0 5.3405e-08 0.0007 5.3408e-08 0 5.3602e-08 0 5.3605e-08 0.0007 5.3608e-08 0 5.3802e-08 0 5.3805e-08 0.0007 5.3808e-08 0 5.4002e-08 0 5.4005e-08 0.0007 5.4008e-08 0 5.4202e-08 0 5.4205e-08 0.0007 5.4208e-08 0 5.4402e-08 0 5.4405e-08 0.0007 5.4408e-08 0 5.4602e-08 0 5.4605e-08 0.0007 5.4608e-08 0 5.4802e-08 0 5.4805e-08 0.0007 5.4808e-08 0 5.5002e-08 0 5.5005e-08 0.0007 5.5008e-08 0 5.5202e-08 0 5.5205e-08 0.0007 5.5208e-08 0 5.5402e-08 0 5.5405e-08 0.0007 5.5408e-08 0 5.5602e-08 0 5.5605e-08 0.0007 5.5608e-08 0 5.5802e-08 0 5.5805e-08 0.0007 5.5808e-08 0 5.6002e-08 0 5.6005e-08 0.0007 5.6008e-08 0 5.6202e-08 0 5.6205e-08 0.0007 5.6208e-08 0 5.6402e-08 0 5.6405e-08 0.0007 5.6408e-08 0 5.6602e-08 0 5.6605e-08 0.0007 5.6608e-08 0 5.6802e-08 0 5.6805e-08 0.0007 5.6808e-08 0 5.7002e-08 0 5.7005e-08 0.0007 5.7008e-08 0 5.7202e-08 0 5.7205e-08 0.0007 5.7208e-08 0 5.7402e-08 0 5.7405e-08 0.0007 5.7408e-08 0 5.7602e-08 0 5.7605e-08 0.0007 5.7608e-08 0 5.7802e-08 0 5.7805e-08 0.0007 5.7808e-08 0 5.8002e-08 0 5.8005e-08 0.0007 5.8008e-08 0 5.8202e-08 0 5.8205e-08 0.0007 5.8208e-08 0 5.8402e-08 0 5.8405e-08 0.0007 5.8408e-08 0 5.8602e-08 0 5.8605e-08 0.0007 5.8608e-08 0 5.8802e-08 0 5.8805e-08 0.0007 5.8808e-08 0 5.9002e-08 0 5.9005e-08 0.0007 5.9008e-08 0 5.9202e-08 0 5.9205e-08 0.0007 5.9208e-08 0 5.9402e-08 0 5.9405e-08 0.0007 5.9408e-08 0 5.9602e-08 0 5.9605e-08 0.0007 5.9608e-08 0 5.9802e-08 0 5.9805e-08 0.0007 5.9808e-08 0 6.0002e-08 0 6.0005e-08 0.0007 6.0008e-08 0 6.0202e-08 0 6.0205e-08 0.0007 6.0208e-08 0 6.0402e-08 0 6.0405e-08 0.0007 6.0408e-08 0 6.0602e-08 0 6.0605e-08 0.0007 6.0608e-08 0 6.0802e-08 0 6.0805e-08 0.0007 6.0808e-08 0 6.1002e-08 0 6.1005e-08 0.0007 6.1008e-08 0 6.1202e-08 0 6.1205e-08 0.0007 6.1208e-08 0 6.1402e-08 0 6.1405e-08 0.0007 6.1408e-08 0 6.1602e-08 0 6.1605e-08 0.0007 6.1608e-08 0 6.1802e-08 0 6.1805e-08 0.0007 6.1808e-08 0 6.2002e-08 0 6.2005e-08 0.0007 6.2008e-08 0 6.2202e-08 0 6.2205e-08 0.0007 6.2208e-08 0 6.2402e-08 0 6.2405e-08 0.0007 6.2408e-08 0 6.2602e-08 0 6.2605e-08 0.0007 6.2608e-08 0 6.2802e-08 0 6.2805e-08 0.0007 6.2808e-08 0 6.3002e-08 0 6.3005e-08 0.0007 6.3008e-08 0 6.3202e-08 0 6.3205e-08 0.0007 6.3208e-08 0 6.3402e-08 0 6.3405e-08 0.0007 6.3408e-08 0 6.3602e-08 0 6.3605e-08 0.0007 6.3608e-08 0 6.3802e-08 0 6.3805e-08 0.0007 6.3808e-08 0 6.4002e-08 0 6.4005e-08 0.0007 6.4008e-08 0 6.4202e-08 0 6.4205e-08 0.0007 6.4208e-08 0 6.4402e-08 0 6.4405e-08 0.0007 6.4408e-08 0 6.4602e-08 0 6.4605e-08 0.0007 6.4608e-08 0 6.4802e-08 0 6.4805e-08 0.0007 6.4808e-08 0 6.5002e-08 0 6.5005e-08 0.0007 6.5008e-08 0 6.5202e-08 0 6.5205e-08 0.0007 6.5208e-08 0 6.5402e-08 0 6.5405e-08 0.0007 6.5408e-08 0 6.5602e-08 0 6.5605e-08 0.0007 6.5608e-08 0 6.5802e-08 0 6.5805e-08 0.0007 6.5808e-08 0 6.6002e-08 0 6.6005e-08 0.0007 6.6008e-08 0 6.6202e-08 0 6.6205e-08 0.0007 6.6208e-08 0 6.6402e-08 0 6.6405e-08 0.0007 6.6408e-08 0 6.6602e-08 0 6.6605e-08 0.0007 6.6608e-08 0 6.6802e-08 0 6.6805e-08 0.0007 6.6808e-08 0 6.7002e-08 0 6.7005e-08 0.0007 6.7008e-08 0 6.7202e-08 0 6.7205e-08 0.0007 6.7208e-08 0 6.7402e-08 0 6.7405e-08 0.0007 6.7408e-08 0 6.7602e-08 0 6.7605e-08 0.0007 6.7608e-08 0 6.7802e-08 0 6.7805e-08 0.0007 6.7808e-08 0 6.8002e-08 0 6.8005e-08 0.0007 6.8008e-08 0 6.8202e-08 0 6.8205e-08 0.0007 6.8208e-08 0 6.8402e-08 0 6.8405e-08 0.0007 6.8408e-08 0 6.8602e-08 0 6.8605e-08 0.0007 6.8608e-08 0 6.8802e-08 0 6.8805e-08 0.0007 6.8808e-08 0 6.9002e-08 0 6.9005e-08 0.0007 6.9008e-08 0 6.9202e-08 0 6.9205e-08 0.0007 6.9208e-08 0 6.9402e-08 0 6.9405e-08 0.0007 6.9408e-08 0 6.9602e-08 0 6.9605e-08 0.0007 6.9608e-08 0 6.9802e-08 0 6.9805e-08 0.0007 6.9808e-08 0 7.0002e-08 0 7.0005e-08 0.0007 7.0008e-08 0 7.0202e-08 0 7.0205e-08 0.0007 7.0208e-08 0 7.0402e-08 0 7.0405e-08 0.0007 7.0408e-08 0 7.0602e-08 0 7.0605e-08 0.0007 7.0608e-08 0 7.0802e-08 0 7.0805e-08 0.0007 7.0808e-08 0 7.1002e-08 0 7.1005e-08 0.0007 7.1008e-08 0 7.1202e-08 0 7.1205e-08 0.0007 7.1208e-08 0 7.1402e-08 0 7.1405e-08 0.0007 7.1408e-08 0 7.1602e-08 0 7.1605e-08 0.0007 7.1608e-08 0 7.1802e-08 0 7.1805e-08 0.0007 7.1808e-08 0 7.2002e-08 0 7.2005e-08 0.0007 7.2008e-08 0 7.2202e-08 0 7.2205e-08 0.0007 7.2208e-08 0 7.2402e-08 0 7.2405e-08 0.0007 7.2408e-08 0 7.2602e-08 0 7.2605e-08 0.0007 7.2608e-08 0 7.2802e-08 0 7.2805e-08 0.0007 7.2808e-08 0 7.3002e-08 0 7.3005e-08 0.0007 7.3008e-08 0 7.3202e-08 0 7.3205e-08 0.0007 7.3208e-08 0 7.3402e-08 0 7.3405e-08 0.0007 7.3408e-08 0 7.3602e-08 0 7.3605e-08 0.0007 7.3608e-08 0 7.3802e-08 0 7.3805e-08 0.0007 7.3808e-08 0 7.4002e-08 0 7.4005e-08 0.0007 7.4008e-08 0 7.4202e-08 0 7.4205e-08 0.0007 7.4208e-08 0 7.4402e-08 0 7.4405e-08 0.0007 7.4408e-08 0 7.4602e-08 0 7.4605e-08 0.0007 7.4608e-08 0 7.4802e-08 0 7.4805e-08 0.0007 7.4808e-08 0 7.5002e-08 0 7.5005e-08 0.0007 7.5008e-08 0 7.5202e-08 0 7.5205e-08 0.0007 7.5208e-08 0 7.5402e-08 0 7.5405e-08 0.0007 7.5408e-08 0 7.5602e-08 0 7.5605e-08 0.0007 7.5608e-08 0 7.5802e-08 0 7.5805e-08 0.0007 7.5808e-08 0 7.6002e-08 0 7.6005e-08 0.0007 7.6008e-08 0 7.6202e-08 0 7.6205e-08 0.0007 7.6208e-08 0 7.6402e-08 0 7.6405e-08 0.0007 7.6408e-08 0 7.6602e-08 0 7.6605e-08 0.0007 7.6608e-08 0 7.6802e-08 0 7.6805e-08 0.0007 7.6808e-08 0 7.7002e-08 0 7.7005e-08 0.0007 7.7008e-08 0 7.7202e-08 0 7.7205e-08 0.0007 7.7208e-08 0 7.7402e-08 0 7.7405e-08 0.0007 7.7408e-08 0 7.7602e-08 0 7.7605e-08 0.0007 7.7608e-08 0 7.7802e-08 0 7.7805e-08 0.0007 7.7808e-08 0 7.8002e-08 0 7.8005e-08 0.0007 7.8008e-08 0 7.8202e-08 0 7.8205e-08 0.0007 7.8208e-08 0 7.8402e-08 0 7.8405e-08 0.0007 7.8408e-08 0 7.8602e-08 0 7.8605e-08 0.0007 7.8608e-08 0 7.8802e-08 0 7.8805e-08 0.0007 7.8808e-08 0 7.9002e-08 0 7.9005e-08 0.0007 7.9008e-08 0 7.9202e-08 0 7.9205e-08 0.0007 7.9208e-08 0 7.9402e-08 0 7.9405e-08 0.0007 7.9408e-08 0 7.9602e-08 0 7.9605e-08 0.0007 7.9608e-08 0)
L_S0|1 P0_2 _S0|A1  2.067833848e-12
L_S0|2 _S0|A1 _S0|A2  4.135667696e-12
L_S0|3 _S0|A3 _S0|A4  8.271335392e-12
L_S0|T T12 _S0|T1  2.067833848e-12
L_S0|4 _S0|T1 _S0|T2  4.135667696e-12
L_S0|5 _S0|A4 _S0|Q1  4.135667696e-12
L_S0|6 _S0|Q1 S0  2.067833848e-12
IT13|T 0 T13  PWL(0 0 2e-12 0 5e-12 0.0007 8e-12 0 2.02e-10 0 2.05e-10 0.0007 2.08e-10 0 4.02e-10 0 4.05e-10 0.0007 4.08e-10 0 6.02e-10 0 6.05e-10 0.0007 6.08e-10 0 8.02e-10 0 8.05e-10 0.0007 8.08e-10 0 1.002e-09 0 1.005e-09 0.0007 1.008e-09 0 1.202e-09 0 1.205e-09 0.0007 1.208e-09 0 1.402e-09 0 1.405e-09 0.0007 1.408e-09 0 1.602e-09 0 1.605e-09 0.0007 1.608e-09 0 1.802e-09 0 1.805e-09 0.0007 1.808e-09 0 2.002e-09 0 2.005e-09 0.0007 2.008e-09 0 2.202e-09 0 2.205e-09 0.0007 2.208e-09 0 2.402e-09 0 2.405e-09 0.0007 2.408e-09 0 2.602e-09 0 2.605e-09 0.0007 2.608e-09 0 2.802e-09 0 2.805e-09 0.0007 2.808e-09 0 3.002e-09 0 3.005e-09 0.0007 3.008e-09 0 3.202e-09 0 3.205e-09 0.0007 3.208e-09 0 3.402e-09 0 3.405e-09 0.0007 3.408e-09 0 3.602e-09 0 3.605e-09 0.0007 3.608e-09 0 3.802e-09 0 3.805e-09 0.0007 3.808e-09 0 4.002e-09 0 4.005e-09 0.0007 4.008e-09 0 4.202e-09 0 4.205e-09 0.0007 4.208e-09 0 4.402e-09 0 4.405e-09 0.0007 4.408e-09 0 4.602e-09 0 4.605e-09 0.0007 4.608e-09 0 4.802e-09 0 4.805e-09 0.0007 4.808e-09 0 5.002e-09 0 5.005e-09 0.0007 5.008e-09 0 5.202e-09 0 5.205e-09 0.0007 5.208e-09 0 5.402e-09 0 5.405e-09 0.0007 5.408e-09 0 5.602e-09 0 5.605e-09 0.0007 5.608e-09 0 5.802e-09 0 5.805e-09 0.0007 5.808e-09 0 6.002e-09 0 6.005e-09 0.0007 6.008e-09 0 6.202e-09 0 6.205e-09 0.0007 6.208e-09 0 6.402e-09 0 6.405e-09 0.0007 6.408e-09 0 6.602e-09 0 6.605e-09 0.0007 6.608e-09 0 6.802e-09 0 6.805e-09 0.0007 6.808e-09 0 7.002e-09 0 7.005e-09 0.0007 7.008e-09 0 7.202e-09 0 7.205e-09 0.0007 7.208e-09 0 7.402e-09 0 7.405e-09 0.0007 7.408e-09 0 7.602e-09 0 7.605e-09 0.0007 7.608e-09 0 7.802e-09 0 7.805e-09 0.0007 7.808e-09 0 8.002e-09 0 8.005e-09 0.0007 8.008e-09 0 8.202e-09 0 8.205e-09 0.0007 8.208e-09 0 8.402e-09 0 8.405e-09 0.0007 8.408e-09 0 8.602e-09 0 8.605e-09 0.0007 8.608e-09 0 8.802e-09 0 8.805e-09 0.0007 8.808e-09 0 9.002e-09 0 9.005e-09 0.0007 9.008e-09 0 9.202e-09 0 9.205e-09 0.0007 9.208e-09 0 9.402e-09 0 9.405e-09 0.0007 9.408e-09 0 9.602e-09 0 9.605e-09 0.0007 9.608e-09 0 9.802e-09 0 9.805e-09 0.0007 9.808e-09 0 1.0002e-08 0 1.0005e-08 0.0007 1.0008e-08 0 1.0202e-08 0 1.0205e-08 0.0007 1.0208e-08 0 1.0402e-08 0 1.0405e-08 0.0007 1.0408e-08 0 1.0602e-08 0 1.0605e-08 0.0007 1.0608e-08 0 1.0802e-08 0 1.0805e-08 0.0007 1.0808e-08 0 1.1002e-08 0 1.1005e-08 0.0007 1.1008e-08 0 1.1202e-08 0 1.1205e-08 0.0007 1.1208e-08 0 1.1402e-08 0 1.1405e-08 0.0007 1.1408e-08 0 1.1602e-08 0 1.1605e-08 0.0007 1.1608e-08 0 1.1802e-08 0 1.1805e-08 0.0007 1.1808e-08 0 1.2002e-08 0 1.2005e-08 0.0007 1.2008e-08 0 1.2202e-08 0 1.2205e-08 0.0007 1.2208e-08 0 1.2402e-08 0 1.2405e-08 0.0007 1.2408e-08 0 1.2602e-08 0 1.2605e-08 0.0007 1.2608e-08 0 1.2802e-08 0 1.2805e-08 0.0007 1.2808e-08 0 1.3002e-08 0 1.3005e-08 0.0007 1.3008e-08 0 1.3202e-08 0 1.3205e-08 0.0007 1.3208e-08 0 1.3402e-08 0 1.3405e-08 0.0007 1.3408e-08 0 1.3602e-08 0 1.3605e-08 0.0007 1.3608e-08 0 1.3802e-08 0 1.3805e-08 0.0007 1.3808e-08 0 1.4002e-08 0 1.4005e-08 0.0007 1.4008e-08 0 1.4202e-08 0 1.4205e-08 0.0007 1.4208e-08 0 1.4402e-08 0 1.4405e-08 0.0007 1.4408e-08 0 1.4602e-08 0 1.4605e-08 0.0007 1.4608e-08 0 1.4802e-08 0 1.4805e-08 0.0007 1.4808e-08 0 1.5002e-08 0 1.5005e-08 0.0007 1.5008e-08 0 1.5202e-08 0 1.5205e-08 0.0007 1.5208e-08 0 1.5402e-08 0 1.5405e-08 0.0007 1.5408e-08 0 1.5602e-08 0 1.5605e-08 0.0007 1.5608e-08 0 1.5802e-08 0 1.5805e-08 0.0007 1.5808e-08 0 1.6002e-08 0 1.6005e-08 0.0007 1.6008e-08 0 1.6202e-08 0 1.6205e-08 0.0007 1.6208e-08 0 1.6402e-08 0 1.6405e-08 0.0007 1.6408e-08 0 1.6602e-08 0 1.6605e-08 0.0007 1.6608e-08 0 1.6802e-08 0 1.6805e-08 0.0007 1.6808e-08 0 1.7002e-08 0 1.7005e-08 0.0007 1.7008e-08 0 1.7202e-08 0 1.7205e-08 0.0007 1.7208e-08 0 1.7402e-08 0 1.7405e-08 0.0007 1.7408e-08 0 1.7602e-08 0 1.7605e-08 0.0007 1.7608e-08 0 1.7802e-08 0 1.7805e-08 0.0007 1.7808e-08 0 1.8002e-08 0 1.8005e-08 0.0007 1.8008e-08 0 1.8202e-08 0 1.8205e-08 0.0007 1.8208e-08 0 1.8402e-08 0 1.8405e-08 0.0007 1.8408e-08 0 1.8602e-08 0 1.8605e-08 0.0007 1.8608e-08 0 1.8802e-08 0 1.8805e-08 0.0007 1.8808e-08 0 1.9002e-08 0 1.9005e-08 0.0007 1.9008e-08 0 1.9202e-08 0 1.9205e-08 0.0007 1.9208e-08 0 1.9402e-08 0 1.9405e-08 0.0007 1.9408e-08 0 1.9602e-08 0 1.9605e-08 0.0007 1.9608e-08 0 1.9802e-08 0 1.9805e-08 0.0007 1.9808e-08 0 2.0002e-08 0 2.0005e-08 0.0007 2.0008e-08 0 2.0202e-08 0 2.0205e-08 0.0007 2.0208e-08 0 2.0402e-08 0 2.0405e-08 0.0007 2.0408e-08 0 2.0602e-08 0 2.0605e-08 0.0007 2.0608e-08 0 2.0802e-08 0 2.0805e-08 0.0007 2.0808e-08 0 2.1002e-08 0 2.1005e-08 0.0007 2.1008e-08 0 2.1202e-08 0 2.1205e-08 0.0007 2.1208e-08 0 2.1402e-08 0 2.1405e-08 0.0007 2.1408e-08 0 2.1602e-08 0 2.1605e-08 0.0007 2.1608e-08 0 2.1802e-08 0 2.1805e-08 0.0007 2.1808e-08 0 2.2002e-08 0 2.2005e-08 0.0007 2.2008e-08 0 2.2202e-08 0 2.2205e-08 0.0007 2.2208e-08 0 2.2402e-08 0 2.2405e-08 0.0007 2.2408e-08 0 2.2602e-08 0 2.2605e-08 0.0007 2.2608e-08 0 2.2802e-08 0 2.2805e-08 0.0007 2.2808e-08 0 2.3002e-08 0 2.3005e-08 0.0007 2.3008e-08 0 2.3202e-08 0 2.3205e-08 0.0007 2.3208e-08 0 2.3402e-08 0 2.3405e-08 0.0007 2.3408e-08 0 2.3602e-08 0 2.3605e-08 0.0007 2.3608e-08 0 2.3802e-08 0 2.3805e-08 0.0007 2.3808e-08 0 2.4002e-08 0 2.4005e-08 0.0007 2.4008e-08 0 2.4202e-08 0 2.4205e-08 0.0007 2.4208e-08 0 2.4402e-08 0 2.4405e-08 0.0007 2.4408e-08 0 2.4602e-08 0 2.4605e-08 0.0007 2.4608e-08 0 2.4802e-08 0 2.4805e-08 0.0007 2.4808e-08 0 2.5002e-08 0 2.5005e-08 0.0007 2.5008e-08 0 2.5202e-08 0 2.5205e-08 0.0007 2.5208e-08 0 2.5402e-08 0 2.5405e-08 0.0007 2.5408e-08 0 2.5602e-08 0 2.5605e-08 0.0007 2.5608e-08 0 2.5802e-08 0 2.5805e-08 0.0007 2.5808e-08 0 2.6002e-08 0 2.6005e-08 0.0007 2.6008e-08 0 2.6202e-08 0 2.6205e-08 0.0007 2.6208e-08 0 2.6402e-08 0 2.6405e-08 0.0007 2.6408e-08 0 2.6602e-08 0 2.6605e-08 0.0007 2.6608e-08 0 2.6802e-08 0 2.6805e-08 0.0007 2.6808e-08 0 2.7002e-08 0 2.7005e-08 0.0007 2.7008e-08 0 2.7202e-08 0 2.7205e-08 0.0007 2.7208e-08 0 2.7402e-08 0 2.7405e-08 0.0007 2.7408e-08 0 2.7602e-08 0 2.7605e-08 0.0007 2.7608e-08 0 2.7802e-08 0 2.7805e-08 0.0007 2.7808e-08 0 2.8002e-08 0 2.8005e-08 0.0007 2.8008e-08 0 2.8202e-08 0 2.8205e-08 0.0007 2.8208e-08 0 2.8402e-08 0 2.8405e-08 0.0007 2.8408e-08 0 2.8602e-08 0 2.8605e-08 0.0007 2.8608e-08 0 2.8802e-08 0 2.8805e-08 0.0007 2.8808e-08 0 2.9002e-08 0 2.9005e-08 0.0007 2.9008e-08 0 2.9202e-08 0 2.9205e-08 0.0007 2.9208e-08 0 2.9402e-08 0 2.9405e-08 0.0007 2.9408e-08 0 2.9602e-08 0 2.9605e-08 0.0007 2.9608e-08 0 2.9802e-08 0 2.9805e-08 0.0007 2.9808e-08 0 3.0002e-08 0 3.0005e-08 0.0007 3.0008e-08 0 3.0202e-08 0 3.0205e-08 0.0007 3.0208e-08 0 3.0402e-08 0 3.0405e-08 0.0007 3.0408e-08 0 3.0602e-08 0 3.0605e-08 0.0007 3.0608e-08 0 3.0802e-08 0 3.0805e-08 0.0007 3.0808e-08 0 3.1002e-08 0 3.1005e-08 0.0007 3.1008e-08 0 3.1202e-08 0 3.1205e-08 0.0007 3.1208e-08 0 3.1402e-08 0 3.1405e-08 0.0007 3.1408e-08 0 3.1602e-08 0 3.1605e-08 0.0007 3.1608e-08 0 3.1802e-08 0 3.1805e-08 0.0007 3.1808e-08 0 3.2002e-08 0 3.2005e-08 0.0007 3.2008e-08 0 3.2202e-08 0 3.2205e-08 0.0007 3.2208e-08 0 3.2402e-08 0 3.2405e-08 0.0007 3.2408e-08 0 3.2602e-08 0 3.2605e-08 0.0007 3.2608e-08 0 3.2802e-08 0 3.2805e-08 0.0007 3.2808e-08 0 3.3002e-08 0 3.3005e-08 0.0007 3.3008e-08 0 3.3202e-08 0 3.3205e-08 0.0007 3.3208e-08 0 3.3402e-08 0 3.3405e-08 0.0007 3.3408e-08 0 3.3602e-08 0 3.3605e-08 0.0007 3.3608e-08 0 3.3802e-08 0 3.3805e-08 0.0007 3.3808e-08 0 3.4002e-08 0 3.4005e-08 0.0007 3.4008e-08 0 3.4202e-08 0 3.4205e-08 0.0007 3.4208e-08 0 3.4402e-08 0 3.4405e-08 0.0007 3.4408e-08 0 3.4602e-08 0 3.4605e-08 0.0007 3.4608e-08 0 3.4802e-08 0 3.4805e-08 0.0007 3.4808e-08 0 3.5002e-08 0 3.5005e-08 0.0007 3.5008e-08 0 3.5202e-08 0 3.5205e-08 0.0007 3.5208e-08 0 3.5402e-08 0 3.5405e-08 0.0007 3.5408e-08 0 3.5602e-08 0 3.5605e-08 0.0007 3.5608e-08 0 3.5802e-08 0 3.5805e-08 0.0007 3.5808e-08 0 3.6002e-08 0 3.6005e-08 0.0007 3.6008e-08 0 3.6202e-08 0 3.6205e-08 0.0007 3.6208e-08 0 3.6402e-08 0 3.6405e-08 0.0007 3.6408e-08 0 3.6602e-08 0 3.6605e-08 0.0007 3.6608e-08 0 3.6802e-08 0 3.6805e-08 0.0007 3.6808e-08 0 3.7002e-08 0 3.7005e-08 0.0007 3.7008e-08 0 3.7202e-08 0 3.7205e-08 0.0007 3.7208e-08 0 3.7402e-08 0 3.7405e-08 0.0007 3.7408e-08 0 3.7602e-08 0 3.7605e-08 0.0007 3.7608e-08 0 3.7802e-08 0 3.7805e-08 0.0007 3.7808e-08 0 3.8002e-08 0 3.8005e-08 0.0007 3.8008e-08 0 3.8202e-08 0 3.8205e-08 0.0007 3.8208e-08 0 3.8402e-08 0 3.8405e-08 0.0007 3.8408e-08 0 3.8602e-08 0 3.8605e-08 0.0007 3.8608e-08 0 3.8802e-08 0 3.8805e-08 0.0007 3.8808e-08 0 3.9002e-08 0 3.9005e-08 0.0007 3.9008e-08 0 3.9202e-08 0 3.9205e-08 0.0007 3.9208e-08 0 3.9402e-08 0 3.9405e-08 0.0007 3.9408e-08 0 3.9602e-08 0 3.9605e-08 0.0007 3.9608e-08 0 3.9802e-08 0 3.9805e-08 0.0007 3.9808e-08 0 4.0002e-08 0 4.0005e-08 0.0007 4.0008e-08 0 4.0202e-08 0 4.0205e-08 0.0007 4.0208e-08 0 4.0402e-08 0 4.0405e-08 0.0007 4.0408e-08 0 4.0602e-08 0 4.0605e-08 0.0007 4.0608e-08 0 4.0802e-08 0 4.0805e-08 0.0007 4.0808e-08 0 4.1002e-08 0 4.1005e-08 0.0007 4.1008e-08 0 4.1202e-08 0 4.1205e-08 0.0007 4.1208e-08 0 4.1402e-08 0 4.1405e-08 0.0007 4.1408e-08 0 4.1602e-08 0 4.1605e-08 0.0007 4.1608e-08 0 4.1802e-08 0 4.1805e-08 0.0007 4.1808e-08 0 4.2002e-08 0 4.2005e-08 0.0007 4.2008e-08 0 4.2202e-08 0 4.2205e-08 0.0007 4.2208e-08 0 4.2402e-08 0 4.2405e-08 0.0007 4.2408e-08 0 4.2602e-08 0 4.2605e-08 0.0007 4.2608e-08 0 4.2802e-08 0 4.2805e-08 0.0007 4.2808e-08 0 4.3002e-08 0 4.3005e-08 0.0007 4.3008e-08 0 4.3202e-08 0 4.3205e-08 0.0007 4.3208e-08 0 4.3402e-08 0 4.3405e-08 0.0007 4.3408e-08 0 4.3602e-08 0 4.3605e-08 0.0007 4.3608e-08 0 4.3802e-08 0 4.3805e-08 0.0007 4.3808e-08 0 4.4002e-08 0 4.4005e-08 0.0007 4.4008e-08 0 4.4202e-08 0 4.4205e-08 0.0007 4.4208e-08 0 4.4402e-08 0 4.4405e-08 0.0007 4.4408e-08 0 4.4602e-08 0 4.4605e-08 0.0007 4.4608e-08 0 4.4802e-08 0 4.4805e-08 0.0007 4.4808e-08 0 4.5002e-08 0 4.5005e-08 0.0007 4.5008e-08 0 4.5202e-08 0 4.5205e-08 0.0007 4.5208e-08 0 4.5402e-08 0 4.5405e-08 0.0007 4.5408e-08 0 4.5602e-08 0 4.5605e-08 0.0007 4.5608e-08 0 4.5802e-08 0 4.5805e-08 0.0007 4.5808e-08 0 4.6002e-08 0 4.6005e-08 0.0007 4.6008e-08 0 4.6202e-08 0 4.6205e-08 0.0007 4.6208e-08 0 4.6402e-08 0 4.6405e-08 0.0007 4.6408e-08 0 4.6602e-08 0 4.6605e-08 0.0007 4.6608e-08 0 4.6802e-08 0 4.6805e-08 0.0007 4.6808e-08 0 4.7002e-08 0 4.7005e-08 0.0007 4.7008e-08 0 4.7202e-08 0 4.7205e-08 0.0007 4.7208e-08 0 4.7402e-08 0 4.7405e-08 0.0007 4.7408e-08 0 4.7602e-08 0 4.7605e-08 0.0007 4.7608e-08 0 4.7802e-08 0 4.7805e-08 0.0007 4.7808e-08 0 4.8002e-08 0 4.8005e-08 0.0007 4.8008e-08 0 4.8202e-08 0 4.8205e-08 0.0007 4.8208e-08 0 4.8402e-08 0 4.8405e-08 0.0007 4.8408e-08 0 4.8602e-08 0 4.8605e-08 0.0007 4.8608e-08 0 4.8802e-08 0 4.8805e-08 0.0007 4.8808e-08 0 4.9002e-08 0 4.9005e-08 0.0007 4.9008e-08 0 4.9202e-08 0 4.9205e-08 0.0007 4.9208e-08 0 4.9402e-08 0 4.9405e-08 0.0007 4.9408e-08 0 4.9602e-08 0 4.9605e-08 0.0007 4.9608e-08 0 4.9802e-08 0 4.9805e-08 0.0007 4.9808e-08 0 5.0002e-08 0 5.0005e-08 0.0007 5.0008e-08 0 5.0202e-08 0 5.0205e-08 0.0007 5.0208e-08 0 5.0402e-08 0 5.0405e-08 0.0007 5.0408e-08 0 5.0602e-08 0 5.0605e-08 0.0007 5.0608e-08 0 5.0802e-08 0 5.0805e-08 0.0007 5.0808e-08 0 5.1002e-08 0 5.1005e-08 0.0007 5.1008e-08 0 5.1202e-08 0 5.1205e-08 0.0007 5.1208e-08 0 5.1402e-08 0 5.1405e-08 0.0007 5.1408e-08 0 5.1602e-08 0 5.1605e-08 0.0007 5.1608e-08 0 5.1802e-08 0 5.1805e-08 0.0007 5.1808e-08 0 5.2002e-08 0 5.2005e-08 0.0007 5.2008e-08 0 5.2202e-08 0 5.2205e-08 0.0007 5.2208e-08 0 5.2402e-08 0 5.2405e-08 0.0007 5.2408e-08 0 5.2602e-08 0 5.2605e-08 0.0007 5.2608e-08 0 5.2802e-08 0 5.2805e-08 0.0007 5.2808e-08 0 5.3002e-08 0 5.3005e-08 0.0007 5.3008e-08 0 5.3202e-08 0 5.3205e-08 0.0007 5.3208e-08 0 5.3402e-08 0 5.3405e-08 0.0007 5.3408e-08 0 5.3602e-08 0 5.3605e-08 0.0007 5.3608e-08 0 5.3802e-08 0 5.3805e-08 0.0007 5.3808e-08 0 5.4002e-08 0 5.4005e-08 0.0007 5.4008e-08 0 5.4202e-08 0 5.4205e-08 0.0007 5.4208e-08 0 5.4402e-08 0 5.4405e-08 0.0007 5.4408e-08 0 5.4602e-08 0 5.4605e-08 0.0007 5.4608e-08 0 5.4802e-08 0 5.4805e-08 0.0007 5.4808e-08 0 5.5002e-08 0 5.5005e-08 0.0007 5.5008e-08 0 5.5202e-08 0 5.5205e-08 0.0007 5.5208e-08 0 5.5402e-08 0 5.5405e-08 0.0007 5.5408e-08 0 5.5602e-08 0 5.5605e-08 0.0007 5.5608e-08 0 5.5802e-08 0 5.5805e-08 0.0007 5.5808e-08 0 5.6002e-08 0 5.6005e-08 0.0007 5.6008e-08 0 5.6202e-08 0 5.6205e-08 0.0007 5.6208e-08 0 5.6402e-08 0 5.6405e-08 0.0007 5.6408e-08 0 5.6602e-08 0 5.6605e-08 0.0007 5.6608e-08 0 5.6802e-08 0 5.6805e-08 0.0007 5.6808e-08 0 5.7002e-08 0 5.7005e-08 0.0007 5.7008e-08 0 5.7202e-08 0 5.7205e-08 0.0007 5.7208e-08 0 5.7402e-08 0 5.7405e-08 0.0007 5.7408e-08 0 5.7602e-08 0 5.7605e-08 0.0007 5.7608e-08 0 5.7802e-08 0 5.7805e-08 0.0007 5.7808e-08 0 5.8002e-08 0 5.8005e-08 0.0007 5.8008e-08 0 5.8202e-08 0 5.8205e-08 0.0007 5.8208e-08 0 5.8402e-08 0 5.8405e-08 0.0007 5.8408e-08 0 5.8602e-08 0 5.8605e-08 0.0007 5.8608e-08 0 5.8802e-08 0 5.8805e-08 0.0007 5.8808e-08 0 5.9002e-08 0 5.9005e-08 0.0007 5.9008e-08 0 5.9202e-08 0 5.9205e-08 0.0007 5.9208e-08 0 5.9402e-08 0 5.9405e-08 0.0007 5.9408e-08 0 5.9602e-08 0 5.9605e-08 0.0007 5.9608e-08 0 5.9802e-08 0 5.9805e-08 0.0007 5.9808e-08 0 6.0002e-08 0 6.0005e-08 0.0007 6.0008e-08 0 6.0202e-08 0 6.0205e-08 0.0007 6.0208e-08 0 6.0402e-08 0 6.0405e-08 0.0007 6.0408e-08 0 6.0602e-08 0 6.0605e-08 0.0007 6.0608e-08 0 6.0802e-08 0 6.0805e-08 0.0007 6.0808e-08 0 6.1002e-08 0 6.1005e-08 0.0007 6.1008e-08 0 6.1202e-08 0 6.1205e-08 0.0007 6.1208e-08 0 6.1402e-08 0 6.1405e-08 0.0007 6.1408e-08 0 6.1602e-08 0 6.1605e-08 0.0007 6.1608e-08 0 6.1802e-08 0 6.1805e-08 0.0007 6.1808e-08 0 6.2002e-08 0 6.2005e-08 0.0007 6.2008e-08 0 6.2202e-08 0 6.2205e-08 0.0007 6.2208e-08 0 6.2402e-08 0 6.2405e-08 0.0007 6.2408e-08 0 6.2602e-08 0 6.2605e-08 0.0007 6.2608e-08 0 6.2802e-08 0 6.2805e-08 0.0007 6.2808e-08 0 6.3002e-08 0 6.3005e-08 0.0007 6.3008e-08 0 6.3202e-08 0 6.3205e-08 0.0007 6.3208e-08 0 6.3402e-08 0 6.3405e-08 0.0007 6.3408e-08 0 6.3602e-08 0 6.3605e-08 0.0007 6.3608e-08 0 6.3802e-08 0 6.3805e-08 0.0007 6.3808e-08 0 6.4002e-08 0 6.4005e-08 0.0007 6.4008e-08 0 6.4202e-08 0 6.4205e-08 0.0007 6.4208e-08 0 6.4402e-08 0 6.4405e-08 0.0007 6.4408e-08 0 6.4602e-08 0 6.4605e-08 0.0007 6.4608e-08 0 6.4802e-08 0 6.4805e-08 0.0007 6.4808e-08 0 6.5002e-08 0 6.5005e-08 0.0007 6.5008e-08 0 6.5202e-08 0 6.5205e-08 0.0007 6.5208e-08 0 6.5402e-08 0 6.5405e-08 0.0007 6.5408e-08 0 6.5602e-08 0 6.5605e-08 0.0007 6.5608e-08 0 6.5802e-08 0 6.5805e-08 0.0007 6.5808e-08 0 6.6002e-08 0 6.6005e-08 0.0007 6.6008e-08 0 6.6202e-08 0 6.6205e-08 0.0007 6.6208e-08 0 6.6402e-08 0 6.6405e-08 0.0007 6.6408e-08 0 6.6602e-08 0 6.6605e-08 0.0007 6.6608e-08 0 6.6802e-08 0 6.6805e-08 0.0007 6.6808e-08 0 6.7002e-08 0 6.7005e-08 0.0007 6.7008e-08 0 6.7202e-08 0 6.7205e-08 0.0007 6.7208e-08 0 6.7402e-08 0 6.7405e-08 0.0007 6.7408e-08 0 6.7602e-08 0 6.7605e-08 0.0007 6.7608e-08 0 6.7802e-08 0 6.7805e-08 0.0007 6.7808e-08 0 6.8002e-08 0 6.8005e-08 0.0007 6.8008e-08 0 6.8202e-08 0 6.8205e-08 0.0007 6.8208e-08 0 6.8402e-08 0 6.8405e-08 0.0007 6.8408e-08 0 6.8602e-08 0 6.8605e-08 0.0007 6.8608e-08 0 6.8802e-08 0 6.8805e-08 0.0007 6.8808e-08 0 6.9002e-08 0 6.9005e-08 0.0007 6.9008e-08 0 6.9202e-08 0 6.9205e-08 0.0007 6.9208e-08 0 6.9402e-08 0 6.9405e-08 0.0007 6.9408e-08 0 6.9602e-08 0 6.9605e-08 0.0007 6.9608e-08 0 6.9802e-08 0 6.9805e-08 0.0007 6.9808e-08 0 7.0002e-08 0 7.0005e-08 0.0007 7.0008e-08 0 7.0202e-08 0 7.0205e-08 0.0007 7.0208e-08 0 7.0402e-08 0 7.0405e-08 0.0007 7.0408e-08 0 7.0602e-08 0 7.0605e-08 0.0007 7.0608e-08 0 7.0802e-08 0 7.0805e-08 0.0007 7.0808e-08 0 7.1002e-08 0 7.1005e-08 0.0007 7.1008e-08 0 7.1202e-08 0 7.1205e-08 0.0007 7.1208e-08 0 7.1402e-08 0 7.1405e-08 0.0007 7.1408e-08 0 7.1602e-08 0 7.1605e-08 0.0007 7.1608e-08 0 7.1802e-08 0 7.1805e-08 0.0007 7.1808e-08 0 7.2002e-08 0 7.2005e-08 0.0007 7.2008e-08 0 7.2202e-08 0 7.2205e-08 0.0007 7.2208e-08 0 7.2402e-08 0 7.2405e-08 0.0007 7.2408e-08 0 7.2602e-08 0 7.2605e-08 0.0007 7.2608e-08 0 7.2802e-08 0 7.2805e-08 0.0007 7.2808e-08 0 7.3002e-08 0 7.3005e-08 0.0007 7.3008e-08 0 7.3202e-08 0 7.3205e-08 0.0007 7.3208e-08 0 7.3402e-08 0 7.3405e-08 0.0007 7.3408e-08 0 7.3602e-08 0 7.3605e-08 0.0007 7.3608e-08 0 7.3802e-08 0 7.3805e-08 0.0007 7.3808e-08 0 7.4002e-08 0 7.4005e-08 0.0007 7.4008e-08 0 7.4202e-08 0 7.4205e-08 0.0007 7.4208e-08 0 7.4402e-08 0 7.4405e-08 0.0007 7.4408e-08 0 7.4602e-08 0 7.4605e-08 0.0007 7.4608e-08 0 7.4802e-08 0 7.4805e-08 0.0007 7.4808e-08 0 7.5002e-08 0 7.5005e-08 0.0007 7.5008e-08 0 7.5202e-08 0 7.5205e-08 0.0007 7.5208e-08 0 7.5402e-08 0 7.5405e-08 0.0007 7.5408e-08 0 7.5602e-08 0 7.5605e-08 0.0007 7.5608e-08 0 7.5802e-08 0 7.5805e-08 0.0007 7.5808e-08 0 7.6002e-08 0 7.6005e-08 0.0007 7.6008e-08 0 7.6202e-08 0 7.6205e-08 0.0007 7.6208e-08 0 7.6402e-08 0 7.6405e-08 0.0007 7.6408e-08 0 7.6602e-08 0 7.6605e-08 0.0007 7.6608e-08 0 7.6802e-08 0 7.6805e-08 0.0007 7.6808e-08 0 7.7002e-08 0 7.7005e-08 0.0007 7.7008e-08 0 7.7202e-08 0 7.7205e-08 0.0007 7.7208e-08 0 7.7402e-08 0 7.7405e-08 0.0007 7.7408e-08 0 7.7602e-08 0 7.7605e-08 0.0007 7.7608e-08 0 7.7802e-08 0 7.7805e-08 0.0007 7.7808e-08 0 7.8002e-08 0 7.8005e-08 0.0007 7.8008e-08 0 7.8202e-08 0 7.8205e-08 0.0007 7.8208e-08 0 7.8402e-08 0 7.8405e-08 0.0007 7.8408e-08 0 7.8602e-08 0 7.8605e-08 0.0007 7.8608e-08 0 7.8802e-08 0 7.8805e-08 0.0007 7.8808e-08 0 7.9002e-08 0 7.9005e-08 0.0007 7.9008e-08 0 7.9202e-08 0 7.9205e-08 0.0007 7.9208e-08 0 7.9402e-08 0 7.9405e-08 0.0007 7.9408e-08 0 7.9602e-08 0 7.9605e-08 0.0007 7.9608e-08 0)
BBUF_G0_2_TMP|1 BUF_G0_2_TMP|1 BUF_G0_2_TMP|2 JJMIT AREA=2.5
BBUF_G0_2_TMP|2 BUF_G0_2_TMP|4 BUF_G0_2_TMP|5 JJMIT AREA=2.5
BBUF_G0_2_TMP|3 BUF_G0_2_TMP|7 BUF_G0_2_TMP|8 JJMIT AREA=2.5
BBUF_G0_2_TMP|4 BUF_G0_2_TMP|10 BUF_G0_2_TMP|11 JJMIT AREA=2.5
IBUF_G0_2_TMP|B1 0 BUF_G0_2_TMP|3  PWL(0 0 5e-12 0.000175)
IBUF_G0_2_TMP|B2 0 BUF_G0_2_TMP|6  PWL(0 0 5e-12 0.0002375)
IBUF_G0_2_TMP|B3 0 BUF_G0_2_TMP|9  PWL(0 0 5e-12 0.0002375)
IBUF_G0_2_TMP|B4 0 BUF_G0_2_TMP|12  PWL(0 0 5e-12 0.000175)
LBUF_G0_2_TMP|1 G0_2 BUF_G0_2_TMP|1  2.067833848e-12
LBUF_G0_2_TMP|2 BUF_G0_2_TMP|1 BUF_G0_2_TMP|4  4.135667696e-12
LBUF_G0_2_TMP|3 BUF_G0_2_TMP|4 BUF_G0_2_TMP|7  4.135667696e-12
LBUF_G0_2_TMP|4 BUF_G0_2_TMP|7 BUF_G0_2_TMP|10  4.135667696e-12
LBUF_G0_2_TMP|5 BUF_G0_2_TMP|10 G0_2_TMP  2.067833848e-12
LBUF_G0_2_TMP|P1 BUF_G0_2_TMP|2 0  5e-13
LBUF_G0_2_TMP|P2 BUF_G0_2_TMP|5 0  5e-13
LBUF_G0_2_TMP|P3 BUF_G0_2_TMP|8 0  5e-13
LBUF_G0_2_TMP|P4 BUF_G0_2_TMP|11 0  5e-13
LBUF_G0_2_TMP|B1 BUF_G0_2_TMP|1 BUF_G0_2_TMP|3  2e-12
LBUF_G0_2_TMP|B2 BUF_G0_2_TMP|4 BUF_G0_2_TMP|6  2e-12
LBUF_G0_2_TMP|B3 BUF_G0_2_TMP|7 BUF_G0_2_TMP|9  2e-12
LBUF_G0_2_TMP|B4 BUF_G0_2_TMP|10 BUF_G0_2_TMP|12  2e-12
RBUF_G0_2_TMP|B1 BUF_G0_2_TMP|1 BUF_G0_2_TMP|101  2.7439617672
RBUF_G0_2_TMP|B2 BUF_G0_2_TMP|4 BUF_G0_2_TMP|104  2.7439617672
RBUF_G0_2_TMP|B3 BUF_G0_2_TMP|7 BUF_G0_2_TMP|107  2.7439617672
RBUF_G0_2_TMP|B4 BUF_G0_2_TMP|10 BUF_G0_2_TMP|110  2.7439617672
LBUF_G0_2_TMP|RB1 BUF_G0_2_TMP|101 0  2.050338398468e-12
LBUF_G0_2_TMP|RB2 BUF_G0_2_TMP|104 0  2.050338398468e-12
LBUF_G0_2_TMP|RB3 BUF_G0_2_TMP|107 0  2.050338398468e-12
LBUF_G0_2_TMP|RB4 BUF_G0_2_TMP|110 0  2.050338398468e-12
LBUF_G0_2|1 G0_2_TMP BUF_G0_2|1  2.067833848e-12
LBUF_G0_2|2 BUF_G0_2|1 BUF_G0_2|4  2.067833848e-12
LBUF_G0_2|3 BUF_G0_2|4 BUF_G0_2|6  2.067833848e-12
LBUF_G0_2|4 BUF_G0_2|6 G0_2_BUF  2.067833848e-12
BBUF_IP1_2_TMP|1 BUF_IP1_2_TMP|1 BUF_IP1_2_TMP|2 JJMIT AREA=2.5
BBUF_IP1_2_TMP|2 BUF_IP1_2_TMP|4 BUF_IP1_2_TMP|5 JJMIT AREA=2.5
BBUF_IP1_2_TMP|3 BUF_IP1_2_TMP|7 BUF_IP1_2_TMP|8 JJMIT AREA=2.5
BBUF_IP1_2_TMP|4 BUF_IP1_2_TMP|10 BUF_IP1_2_TMP|11 JJMIT AREA=2.5
IBUF_IP1_2_TMP|B1 0 BUF_IP1_2_TMP|3  PWL(0 0 5e-12 0.000175)
IBUF_IP1_2_TMP|B2 0 BUF_IP1_2_TMP|6  PWL(0 0 5e-12 0.0002375)
IBUF_IP1_2_TMP|B3 0 BUF_IP1_2_TMP|9  PWL(0 0 5e-12 0.0002375)
IBUF_IP1_2_TMP|B4 0 BUF_IP1_2_TMP|12  PWL(0 0 5e-12 0.000175)
LBUF_IP1_2_TMP|1 IP1_2_OUT BUF_IP1_2_TMP|1  2.067833848e-12
LBUF_IP1_2_TMP|2 BUF_IP1_2_TMP|1 BUF_IP1_2_TMP|4  4.135667696e-12
LBUF_IP1_2_TMP|3 BUF_IP1_2_TMP|4 BUF_IP1_2_TMP|7  4.135667696e-12
LBUF_IP1_2_TMP|4 BUF_IP1_2_TMP|7 BUF_IP1_2_TMP|10  4.135667696e-12
LBUF_IP1_2_TMP|5 BUF_IP1_2_TMP|10 IP1_2_TMP  2.067833848e-12
LBUF_IP1_2_TMP|P1 BUF_IP1_2_TMP|2 0  5e-13
LBUF_IP1_2_TMP|P2 BUF_IP1_2_TMP|5 0  5e-13
LBUF_IP1_2_TMP|P3 BUF_IP1_2_TMP|8 0  5e-13
LBUF_IP1_2_TMP|P4 BUF_IP1_2_TMP|11 0  5e-13
LBUF_IP1_2_TMP|B1 BUF_IP1_2_TMP|1 BUF_IP1_2_TMP|3  2e-12
LBUF_IP1_2_TMP|B2 BUF_IP1_2_TMP|4 BUF_IP1_2_TMP|6  2e-12
LBUF_IP1_2_TMP|B3 BUF_IP1_2_TMP|7 BUF_IP1_2_TMP|9  2e-12
LBUF_IP1_2_TMP|B4 BUF_IP1_2_TMP|10 BUF_IP1_2_TMP|12  2e-12
RBUF_IP1_2_TMP|B1 BUF_IP1_2_TMP|1 BUF_IP1_2_TMP|101  2.7439617672
RBUF_IP1_2_TMP|B2 BUF_IP1_2_TMP|4 BUF_IP1_2_TMP|104  2.7439617672
RBUF_IP1_2_TMP|B3 BUF_IP1_2_TMP|7 BUF_IP1_2_TMP|107  2.7439617672
RBUF_IP1_2_TMP|B4 BUF_IP1_2_TMP|10 BUF_IP1_2_TMP|110  2.7439617672
LBUF_IP1_2_TMP|RB1 BUF_IP1_2_TMP|101 0  2.050338398468e-12
LBUF_IP1_2_TMP|RB2 BUF_IP1_2_TMP|104 0  2.050338398468e-12
LBUF_IP1_2_TMP|RB3 BUF_IP1_2_TMP|107 0  2.050338398468e-12
LBUF_IP1_2_TMP|RB4 BUF_IP1_2_TMP|110 0  2.050338398468e-12
LBUF_IP1_2|1 IP1_2_TMP BUF_IP1_2|1  2.067833848e-12
LBUF_IP1_2|2 BUF_IP1_2|1 BUF_IP1_2|4  2.067833848e-12
LBUF_IP1_2|3 BUF_IP1_2|4 BUF_IP1_2|6  2.067833848e-12
LBUF_IP1_2|4 BUF_IP1_2|6 IP1_2_OUT_BUF  2.067833848e-12
L_S1|A1 G0_2_BUF _S1|A1  2.067833848e-12
L_S1|A2 _S1|A1 _S1|A2  4.135667696e-12
L_S1|A3 _S1|A3 _S1|AB  8.271335392e-12
L_S1|B1 IP1_2_OUT_BUF _S1|B1  2.067833848e-12
L_S1|B2 _S1|B1 _S1|B2  4.135667696e-12
L_S1|B3 _S1|B3 _S1|AB  8.271335392e-12
L_S1|T1 T13 _S1|T1  2.067833848e-12
L_S1|T2 _S1|T1 _S1|T2  4.135667696e-12
L_S1|Q2 _S1|ABTQ _S1|Q1  4.135667696e-12
L_S1|Q1 _S1|Q1 S1  2.067833848e-12
IT14|T 0 T14  PWL(0 0 2e-12 0 5e-12 0.0007 8e-12 0 2.02e-10 0 2.05e-10 0.0007 2.08e-10 0 4.02e-10 0 4.05e-10 0.0007 4.08e-10 0 6.02e-10 0 6.05e-10 0.0007 6.08e-10 0 8.02e-10 0 8.05e-10 0.0007 8.08e-10 0 1.002e-09 0 1.005e-09 0.0007 1.008e-09 0 1.202e-09 0 1.205e-09 0.0007 1.208e-09 0 1.402e-09 0 1.405e-09 0.0007 1.408e-09 0 1.602e-09 0 1.605e-09 0.0007 1.608e-09 0 1.802e-09 0 1.805e-09 0.0007 1.808e-09 0 2.002e-09 0 2.005e-09 0.0007 2.008e-09 0 2.202e-09 0 2.205e-09 0.0007 2.208e-09 0 2.402e-09 0 2.405e-09 0.0007 2.408e-09 0 2.602e-09 0 2.605e-09 0.0007 2.608e-09 0 2.802e-09 0 2.805e-09 0.0007 2.808e-09 0 3.002e-09 0 3.005e-09 0.0007 3.008e-09 0 3.202e-09 0 3.205e-09 0.0007 3.208e-09 0 3.402e-09 0 3.405e-09 0.0007 3.408e-09 0 3.602e-09 0 3.605e-09 0.0007 3.608e-09 0 3.802e-09 0 3.805e-09 0.0007 3.808e-09 0 4.002e-09 0 4.005e-09 0.0007 4.008e-09 0 4.202e-09 0 4.205e-09 0.0007 4.208e-09 0 4.402e-09 0 4.405e-09 0.0007 4.408e-09 0 4.602e-09 0 4.605e-09 0.0007 4.608e-09 0 4.802e-09 0 4.805e-09 0.0007 4.808e-09 0 5.002e-09 0 5.005e-09 0.0007 5.008e-09 0 5.202e-09 0 5.205e-09 0.0007 5.208e-09 0 5.402e-09 0 5.405e-09 0.0007 5.408e-09 0 5.602e-09 0 5.605e-09 0.0007 5.608e-09 0 5.802e-09 0 5.805e-09 0.0007 5.808e-09 0 6.002e-09 0 6.005e-09 0.0007 6.008e-09 0 6.202e-09 0 6.205e-09 0.0007 6.208e-09 0 6.402e-09 0 6.405e-09 0.0007 6.408e-09 0 6.602e-09 0 6.605e-09 0.0007 6.608e-09 0 6.802e-09 0 6.805e-09 0.0007 6.808e-09 0 7.002e-09 0 7.005e-09 0.0007 7.008e-09 0 7.202e-09 0 7.205e-09 0.0007 7.208e-09 0 7.402e-09 0 7.405e-09 0.0007 7.408e-09 0 7.602e-09 0 7.605e-09 0.0007 7.608e-09 0 7.802e-09 0 7.805e-09 0.0007 7.808e-09 0 8.002e-09 0 8.005e-09 0.0007 8.008e-09 0 8.202e-09 0 8.205e-09 0.0007 8.208e-09 0 8.402e-09 0 8.405e-09 0.0007 8.408e-09 0 8.602e-09 0 8.605e-09 0.0007 8.608e-09 0 8.802e-09 0 8.805e-09 0.0007 8.808e-09 0 9.002e-09 0 9.005e-09 0.0007 9.008e-09 0 9.202e-09 0 9.205e-09 0.0007 9.208e-09 0 9.402e-09 0 9.405e-09 0.0007 9.408e-09 0 9.602e-09 0 9.605e-09 0.0007 9.608e-09 0 9.802e-09 0 9.805e-09 0.0007 9.808e-09 0 1.0002e-08 0 1.0005e-08 0.0007 1.0008e-08 0 1.0202e-08 0 1.0205e-08 0.0007 1.0208e-08 0 1.0402e-08 0 1.0405e-08 0.0007 1.0408e-08 0 1.0602e-08 0 1.0605e-08 0.0007 1.0608e-08 0 1.0802e-08 0 1.0805e-08 0.0007 1.0808e-08 0 1.1002e-08 0 1.1005e-08 0.0007 1.1008e-08 0 1.1202e-08 0 1.1205e-08 0.0007 1.1208e-08 0 1.1402e-08 0 1.1405e-08 0.0007 1.1408e-08 0 1.1602e-08 0 1.1605e-08 0.0007 1.1608e-08 0 1.1802e-08 0 1.1805e-08 0.0007 1.1808e-08 0 1.2002e-08 0 1.2005e-08 0.0007 1.2008e-08 0 1.2202e-08 0 1.2205e-08 0.0007 1.2208e-08 0 1.2402e-08 0 1.2405e-08 0.0007 1.2408e-08 0 1.2602e-08 0 1.2605e-08 0.0007 1.2608e-08 0 1.2802e-08 0 1.2805e-08 0.0007 1.2808e-08 0 1.3002e-08 0 1.3005e-08 0.0007 1.3008e-08 0 1.3202e-08 0 1.3205e-08 0.0007 1.3208e-08 0 1.3402e-08 0 1.3405e-08 0.0007 1.3408e-08 0 1.3602e-08 0 1.3605e-08 0.0007 1.3608e-08 0 1.3802e-08 0 1.3805e-08 0.0007 1.3808e-08 0 1.4002e-08 0 1.4005e-08 0.0007 1.4008e-08 0 1.4202e-08 0 1.4205e-08 0.0007 1.4208e-08 0 1.4402e-08 0 1.4405e-08 0.0007 1.4408e-08 0 1.4602e-08 0 1.4605e-08 0.0007 1.4608e-08 0 1.4802e-08 0 1.4805e-08 0.0007 1.4808e-08 0 1.5002e-08 0 1.5005e-08 0.0007 1.5008e-08 0 1.5202e-08 0 1.5205e-08 0.0007 1.5208e-08 0 1.5402e-08 0 1.5405e-08 0.0007 1.5408e-08 0 1.5602e-08 0 1.5605e-08 0.0007 1.5608e-08 0 1.5802e-08 0 1.5805e-08 0.0007 1.5808e-08 0 1.6002e-08 0 1.6005e-08 0.0007 1.6008e-08 0 1.6202e-08 0 1.6205e-08 0.0007 1.6208e-08 0 1.6402e-08 0 1.6405e-08 0.0007 1.6408e-08 0 1.6602e-08 0 1.6605e-08 0.0007 1.6608e-08 0 1.6802e-08 0 1.6805e-08 0.0007 1.6808e-08 0 1.7002e-08 0 1.7005e-08 0.0007 1.7008e-08 0 1.7202e-08 0 1.7205e-08 0.0007 1.7208e-08 0 1.7402e-08 0 1.7405e-08 0.0007 1.7408e-08 0 1.7602e-08 0 1.7605e-08 0.0007 1.7608e-08 0 1.7802e-08 0 1.7805e-08 0.0007 1.7808e-08 0 1.8002e-08 0 1.8005e-08 0.0007 1.8008e-08 0 1.8202e-08 0 1.8205e-08 0.0007 1.8208e-08 0 1.8402e-08 0 1.8405e-08 0.0007 1.8408e-08 0 1.8602e-08 0 1.8605e-08 0.0007 1.8608e-08 0 1.8802e-08 0 1.8805e-08 0.0007 1.8808e-08 0 1.9002e-08 0 1.9005e-08 0.0007 1.9008e-08 0 1.9202e-08 0 1.9205e-08 0.0007 1.9208e-08 0 1.9402e-08 0 1.9405e-08 0.0007 1.9408e-08 0 1.9602e-08 0 1.9605e-08 0.0007 1.9608e-08 0 1.9802e-08 0 1.9805e-08 0.0007 1.9808e-08 0 2.0002e-08 0 2.0005e-08 0.0007 2.0008e-08 0 2.0202e-08 0 2.0205e-08 0.0007 2.0208e-08 0 2.0402e-08 0 2.0405e-08 0.0007 2.0408e-08 0 2.0602e-08 0 2.0605e-08 0.0007 2.0608e-08 0 2.0802e-08 0 2.0805e-08 0.0007 2.0808e-08 0 2.1002e-08 0 2.1005e-08 0.0007 2.1008e-08 0 2.1202e-08 0 2.1205e-08 0.0007 2.1208e-08 0 2.1402e-08 0 2.1405e-08 0.0007 2.1408e-08 0 2.1602e-08 0 2.1605e-08 0.0007 2.1608e-08 0 2.1802e-08 0 2.1805e-08 0.0007 2.1808e-08 0 2.2002e-08 0 2.2005e-08 0.0007 2.2008e-08 0 2.2202e-08 0 2.2205e-08 0.0007 2.2208e-08 0 2.2402e-08 0 2.2405e-08 0.0007 2.2408e-08 0 2.2602e-08 0 2.2605e-08 0.0007 2.2608e-08 0 2.2802e-08 0 2.2805e-08 0.0007 2.2808e-08 0 2.3002e-08 0 2.3005e-08 0.0007 2.3008e-08 0 2.3202e-08 0 2.3205e-08 0.0007 2.3208e-08 0 2.3402e-08 0 2.3405e-08 0.0007 2.3408e-08 0 2.3602e-08 0 2.3605e-08 0.0007 2.3608e-08 0 2.3802e-08 0 2.3805e-08 0.0007 2.3808e-08 0 2.4002e-08 0 2.4005e-08 0.0007 2.4008e-08 0 2.4202e-08 0 2.4205e-08 0.0007 2.4208e-08 0 2.4402e-08 0 2.4405e-08 0.0007 2.4408e-08 0 2.4602e-08 0 2.4605e-08 0.0007 2.4608e-08 0 2.4802e-08 0 2.4805e-08 0.0007 2.4808e-08 0 2.5002e-08 0 2.5005e-08 0.0007 2.5008e-08 0 2.5202e-08 0 2.5205e-08 0.0007 2.5208e-08 0 2.5402e-08 0 2.5405e-08 0.0007 2.5408e-08 0 2.5602e-08 0 2.5605e-08 0.0007 2.5608e-08 0 2.5802e-08 0 2.5805e-08 0.0007 2.5808e-08 0 2.6002e-08 0 2.6005e-08 0.0007 2.6008e-08 0 2.6202e-08 0 2.6205e-08 0.0007 2.6208e-08 0 2.6402e-08 0 2.6405e-08 0.0007 2.6408e-08 0 2.6602e-08 0 2.6605e-08 0.0007 2.6608e-08 0 2.6802e-08 0 2.6805e-08 0.0007 2.6808e-08 0 2.7002e-08 0 2.7005e-08 0.0007 2.7008e-08 0 2.7202e-08 0 2.7205e-08 0.0007 2.7208e-08 0 2.7402e-08 0 2.7405e-08 0.0007 2.7408e-08 0 2.7602e-08 0 2.7605e-08 0.0007 2.7608e-08 0 2.7802e-08 0 2.7805e-08 0.0007 2.7808e-08 0 2.8002e-08 0 2.8005e-08 0.0007 2.8008e-08 0 2.8202e-08 0 2.8205e-08 0.0007 2.8208e-08 0 2.8402e-08 0 2.8405e-08 0.0007 2.8408e-08 0 2.8602e-08 0 2.8605e-08 0.0007 2.8608e-08 0 2.8802e-08 0 2.8805e-08 0.0007 2.8808e-08 0 2.9002e-08 0 2.9005e-08 0.0007 2.9008e-08 0 2.9202e-08 0 2.9205e-08 0.0007 2.9208e-08 0 2.9402e-08 0 2.9405e-08 0.0007 2.9408e-08 0 2.9602e-08 0 2.9605e-08 0.0007 2.9608e-08 0 2.9802e-08 0 2.9805e-08 0.0007 2.9808e-08 0 3.0002e-08 0 3.0005e-08 0.0007 3.0008e-08 0 3.0202e-08 0 3.0205e-08 0.0007 3.0208e-08 0 3.0402e-08 0 3.0405e-08 0.0007 3.0408e-08 0 3.0602e-08 0 3.0605e-08 0.0007 3.0608e-08 0 3.0802e-08 0 3.0805e-08 0.0007 3.0808e-08 0 3.1002e-08 0 3.1005e-08 0.0007 3.1008e-08 0 3.1202e-08 0 3.1205e-08 0.0007 3.1208e-08 0 3.1402e-08 0 3.1405e-08 0.0007 3.1408e-08 0 3.1602e-08 0 3.1605e-08 0.0007 3.1608e-08 0 3.1802e-08 0 3.1805e-08 0.0007 3.1808e-08 0 3.2002e-08 0 3.2005e-08 0.0007 3.2008e-08 0 3.2202e-08 0 3.2205e-08 0.0007 3.2208e-08 0 3.2402e-08 0 3.2405e-08 0.0007 3.2408e-08 0 3.2602e-08 0 3.2605e-08 0.0007 3.2608e-08 0 3.2802e-08 0 3.2805e-08 0.0007 3.2808e-08 0 3.3002e-08 0 3.3005e-08 0.0007 3.3008e-08 0 3.3202e-08 0 3.3205e-08 0.0007 3.3208e-08 0 3.3402e-08 0 3.3405e-08 0.0007 3.3408e-08 0 3.3602e-08 0 3.3605e-08 0.0007 3.3608e-08 0 3.3802e-08 0 3.3805e-08 0.0007 3.3808e-08 0 3.4002e-08 0 3.4005e-08 0.0007 3.4008e-08 0 3.4202e-08 0 3.4205e-08 0.0007 3.4208e-08 0 3.4402e-08 0 3.4405e-08 0.0007 3.4408e-08 0 3.4602e-08 0 3.4605e-08 0.0007 3.4608e-08 0 3.4802e-08 0 3.4805e-08 0.0007 3.4808e-08 0 3.5002e-08 0 3.5005e-08 0.0007 3.5008e-08 0 3.5202e-08 0 3.5205e-08 0.0007 3.5208e-08 0 3.5402e-08 0 3.5405e-08 0.0007 3.5408e-08 0 3.5602e-08 0 3.5605e-08 0.0007 3.5608e-08 0 3.5802e-08 0 3.5805e-08 0.0007 3.5808e-08 0 3.6002e-08 0 3.6005e-08 0.0007 3.6008e-08 0 3.6202e-08 0 3.6205e-08 0.0007 3.6208e-08 0 3.6402e-08 0 3.6405e-08 0.0007 3.6408e-08 0 3.6602e-08 0 3.6605e-08 0.0007 3.6608e-08 0 3.6802e-08 0 3.6805e-08 0.0007 3.6808e-08 0 3.7002e-08 0 3.7005e-08 0.0007 3.7008e-08 0 3.7202e-08 0 3.7205e-08 0.0007 3.7208e-08 0 3.7402e-08 0 3.7405e-08 0.0007 3.7408e-08 0 3.7602e-08 0 3.7605e-08 0.0007 3.7608e-08 0 3.7802e-08 0 3.7805e-08 0.0007 3.7808e-08 0 3.8002e-08 0 3.8005e-08 0.0007 3.8008e-08 0 3.8202e-08 0 3.8205e-08 0.0007 3.8208e-08 0 3.8402e-08 0 3.8405e-08 0.0007 3.8408e-08 0 3.8602e-08 0 3.8605e-08 0.0007 3.8608e-08 0 3.8802e-08 0 3.8805e-08 0.0007 3.8808e-08 0 3.9002e-08 0 3.9005e-08 0.0007 3.9008e-08 0 3.9202e-08 0 3.9205e-08 0.0007 3.9208e-08 0 3.9402e-08 0 3.9405e-08 0.0007 3.9408e-08 0 3.9602e-08 0 3.9605e-08 0.0007 3.9608e-08 0 3.9802e-08 0 3.9805e-08 0.0007 3.9808e-08 0 4.0002e-08 0 4.0005e-08 0.0007 4.0008e-08 0 4.0202e-08 0 4.0205e-08 0.0007 4.0208e-08 0 4.0402e-08 0 4.0405e-08 0.0007 4.0408e-08 0 4.0602e-08 0 4.0605e-08 0.0007 4.0608e-08 0 4.0802e-08 0 4.0805e-08 0.0007 4.0808e-08 0 4.1002e-08 0 4.1005e-08 0.0007 4.1008e-08 0 4.1202e-08 0 4.1205e-08 0.0007 4.1208e-08 0 4.1402e-08 0 4.1405e-08 0.0007 4.1408e-08 0 4.1602e-08 0 4.1605e-08 0.0007 4.1608e-08 0 4.1802e-08 0 4.1805e-08 0.0007 4.1808e-08 0 4.2002e-08 0 4.2005e-08 0.0007 4.2008e-08 0 4.2202e-08 0 4.2205e-08 0.0007 4.2208e-08 0 4.2402e-08 0 4.2405e-08 0.0007 4.2408e-08 0 4.2602e-08 0 4.2605e-08 0.0007 4.2608e-08 0 4.2802e-08 0 4.2805e-08 0.0007 4.2808e-08 0 4.3002e-08 0 4.3005e-08 0.0007 4.3008e-08 0 4.3202e-08 0 4.3205e-08 0.0007 4.3208e-08 0 4.3402e-08 0 4.3405e-08 0.0007 4.3408e-08 0 4.3602e-08 0 4.3605e-08 0.0007 4.3608e-08 0 4.3802e-08 0 4.3805e-08 0.0007 4.3808e-08 0 4.4002e-08 0 4.4005e-08 0.0007 4.4008e-08 0 4.4202e-08 0 4.4205e-08 0.0007 4.4208e-08 0 4.4402e-08 0 4.4405e-08 0.0007 4.4408e-08 0 4.4602e-08 0 4.4605e-08 0.0007 4.4608e-08 0 4.4802e-08 0 4.4805e-08 0.0007 4.4808e-08 0 4.5002e-08 0 4.5005e-08 0.0007 4.5008e-08 0 4.5202e-08 0 4.5205e-08 0.0007 4.5208e-08 0 4.5402e-08 0 4.5405e-08 0.0007 4.5408e-08 0 4.5602e-08 0 4.5605e-08 0.0007 4.5608e-08 0 4.5802e-08 0 4.5805e-08 0.0007 4.5808e-08 0 4.6002e-08 0 4.6005e-08 0.0007 4.6008e-08 0 4.6202e-08 0 4.6205e-08 0.0007 4.6208e-08 0 4.6402e-08 0 4.6405e-08 0.0007 4.6408e-08 0 4.6602e-08 0 4.6605e-08 0.0007 4.6608e-08 0 4.6802e-08 0 4.6805e-08 0.0007 4.6808e-08 0 4.7002e-08 0 4.7005e-08 0.0007 4.7008e-08 0 4.7202e-08 0 4.7205e-08 0.0007 4.7208e-08 0 4.7402e-08 0 4.7405e-08 0.0007 4.7408e-08 0 4.7602e-08 0 4.7605e-08 0.0007 4.7608e-08 0 4.7802e-08 0 4.7805e-08 0.0007 4.7808e-08 0 4.8002e-08 0 4.8005e-08 0.0007 4.8008e-08 0 4.8202e-08 0 4.8205e-08 0.0007 4.8208e-08 0 4.8402e-08 0 4.8405e-08 0.0007 4.8408e-08 0 4.8602e-08 0 4.8605e-08 0.0007 4.8608e-08 0 4.8802e-08 0 4.8805e-08 0.0007 4.8808e-08 0 4.9002e-08 0 4.9005e-08 0.0007 4.9008e-08 0 4.9202e-08 0 4.9205e-08 0.0007 4.9208e-08 0 4.9402e-08 0 4.9405e-08 0.0007 4.9408e-08 0 4.9602e-08 0 4.9605e-08 0.0007 4.9608e-08 0 4.9802e-08 0 4.9805e-08 0.0007 4.9808e-08 0 5.0002e-08 0 5.0005e-08 0.0007 5.0008e-08 0 5.0202e-08 0 5.0205e-08 0.0007 5.0208e-08 0 5.0402e-08 0 5.0405e-08 0.0007 5.0408e-08 0 5.0602e-08 0 5.0605e-08 0.0007 5.0608e-08 0 5.0802e-08 0 5.0805e-08 0.0007 5.0808e-08 0 5.1002e-08 0 5.1005e-08 0.0007 5.1008e-08 0 5.1202e-08 0 5.1205e-08 0.0007 5.1208e-08 0 5.1402e-08 0 5.1405e-08 0.0007 5.1408e-08 0 5.1602e-08 0 5.1605e-08 0.0007 5.1608e-08 0 5.1802e-08 0 5.1805e-08 0.0007 5.1808e-08 0 5.2002e-08 0 5.2005e-08 0.0007 5.2008e-08 0 5.2202e-08 0 5.2205e-08 0.0007 5.2208e-08 0 5.2402e-08 0 5.2405e-08 0.0007 5.2408e-08 0 5.2602e-08 0 5.2605e-08 0.0007 5.2608e-08 0 5.2802e-08 0 5.2805e-08 0.0007 5.2808e-08 0 5.3002e-08 0 5.3005e-08 0.0007 5.3008e-08 0 5.3202e-08 0 5.3205e-08 0.0007 5.3208e-08 0 5.3402e-08 0 5.3405e-08 0.0007 5.3408e-08 0 5.3602e-08 0 5.3605e-08 0.0007 5.3608e-08 0 5.3802e-08 0 5.3805e-08 0.0007 5.3808e-08 0 5.4002e-08 0 5.4005e-08 0.0007 5.4008e-08 0 5.4202e-08 0 5.4205e-08 0.0007 5.4208e-08 0 5.4402e-08 0 5.4405e-08 0.0007 5.4408e-08 0 5.4602e-08 0 5.4605e-08 0.0007 5.4608e-08 0 5.4802e-08 0 5.4805e-08 0.0007 5.4808e-08 0 5.5002e-08 0 5.5005e-08 0.0007 5.5008e-08 0 5.5202e-08 0 5.5205e-08 0.0007 5.5208e-08 0 5.5402e-08 0 5.5405e-08 0.0007 5.5408e-08 0 5.5602e-08 0 5.5605e-08 0.0007 5.5608e-08 0 5.5802e-08 0 5.5805e-08 0.0007 5.5808e-08 0 5.6002e-08 0 5.6005e-08 0.0007 5.6008e-08 0 5.6202e-08 0 5.6205e-08 0.0007 5.6208e-08 0 5.6402e-08 0 5.6405e-08 0.0007 5.6408e-08 0 5.6602e-08 0 5.6605e-08 0.0007 5.6608e-08 0 5.6802e-08 0 5.6805e-08 0.0007 5.6808e-08 0 5.7002e-08 0 5.7005e-08 0.0007 5.7008e-08 0 5.7202e-08 0 5.7205e-08 0.0007 5.7208e-08 0 5.7402e-08 0 5.7405e-08 0.0007 5.7408e-08 0 5.7602e-08 0 5.7605e-08 0.0007 5.7608e-08 0 5.7802e-08 0 5.7805e-08 0.0007 5.7808e-08 0 5.8002e-08 0 5.8005e-08 0.0007 5.8008e-08 0 5.8202e-08 0 5.8205e-08 0.0007 5.8208e-08 0 5.8402e-08 0 5.8405e-08 0.0007 5.8408e-08 0 5.8602e-08 0 5.8605e-08 0.0007 5.8608e-08 0 5.8802e-08 0 5.8805e-08 0.0007 5.8808e-08 0 5.9002e-08 0 5.9005e-08 0.0007 5.9008e-08 0 5.9202e-08 0 5.9205e-08 0.0007 5.9208e-08 0 5.9402e-08 0 5.9405e-08 0.0007 5.9408e-08 0 5.9602e-08 0 5.9605e-08 0.0007 5.9608e-08 0 5.9802e-08 0 5.9805e-08 0.0007 5.9808e-08 0 6.0002e-08 0 6.0005e-08 0.0007 6.0008e-08 0 6.0202e-08 0 6.0205e-08 0.0007 6.0208e-08 0 6.0402e-08 0 6.0405e-08 0.0007 6.0408e-08 0 6.0602e-08 0 6.0605e-08 0.0007 6.0608e-08 0 6.0802e-08 0 6.0805e-08 0.0007 6.0808e-08 0 6.1002e-08 0 6.1005e-08 0.0007 6.1008e-08 0 6.1202e-08 0 6.1205e-08 0.0007 6.1208e-08 0 6.1402e-08 0 6.1405e-08 0.0007 6.1408e-08 0 6.1602e-08 0 6.1605e-08 0.0007 6.1608e-08 0 6.1802e-08 0 6.1805e-08 0.0007 6.1808e-08 0 6.2002e-08 0 6.2005e-08 0.0007 6.2008e-08 0 6.2202e-08 0 6.2205e-08 0.0007 6.2208e-08 0 6.2402e-08 0 6.2405e-08 0.0007 6.2408e-08 0 6.2602e-08 0 6.2605e-08 0.0007 6.2608e-08 0 6.2802e-08 0 6.2805e-08 0.0007 6.2808e-08 0 6.3002e-08 0 6.3005e-08 0.0007 6.3008e-08 0 6.3202e-08 0 6.3205e-08 0.0007 6.3208e-08 0 6.3402e-08 0 6.3405e-08 0.0007 6.3408e-08 0 6.3602e-08 0 6.3605e-08 0.0007 6.3608e-08 0 6.3802e-08 0 6.3805e-08 0.0007 6.3808e-08 0 6.4002e-08 0 6.4005e-08 0.0007 6.4008e-08 0 6.4202e-08 0 6.4205e-08 0.0007 6.4208e-08 0 6.4402e-08 0 6.4405e-08 0.0007 6.4408e-08 0 6.4602e-08 0 6.4605e-08 0.0007 6.4608e-08 0 6.4802e-08 0 6.4805e-08 0.0007 6.4808e-08 0 6.5002e-08 0 6.5005e-08 0.0007 6.5008e-08 0 6.5202e-08 0 6.5205e-08 0.0007 6.5208e-08 0 6.5402e-08 0 6.5405e-08 0.0007 6.5408e-08 0 6.5602e-08 0 6.5605e-08 0.0007 6.5608e-08 0 6.5802e-08 0 6.5805e-08 0.0007 6.5808e-08 0 6.6002e-08 0 6.6005e-08 0.0007 6.6008e-08 0 6.6202e-08 0 6.6205e-08 0.0007 6.6208e-08 0 6.6402e-08 0 6.6405e-08 0.0007 6.6408e-08 0 6.6602e-08 0 6.6605e-08 0.0007 6.6608e-08 0 6.6802e-08 0 6.6805e-08 0.0007 6.6808e-08 0 6.7002e-08 0 6.7005e-08 0.0007 6.7008e-08 0 6.7202e-08 0 6.7205e-08 0.0007 6.7208e-08 0 6.7402e-08 0 6.7405e-08 0.0007 6.7408e-08 0 6.7602e-08 0 6.7605e-08 0.0007 6.7608e-08 0 6.7802e-08 0 6.7805e-08 0.0007 6.7808e-08 0 6.8002e-08 0 6.8005e-08 0.0007 6.8008e-08 0 6.8202e-08 0 6.8205e-08 0.0007 6.8208e-08 0 6.8402e-08 0 6.8405e-08 0.0007 6.8408e-08 0 6.8602e-08 0 6.8605e-08 0.0007 6.8608e-08 0 6.8802e-08 0 6.8805e-08 0.0007 6.8808e-08 0 6.9002e-08 0 6.9005e-08 0.0007 6.9008e-08 0 6.9202e-08 0 6.9205e-08 0.0007 6.9208e-08 0 6.9402e-08 0 6.9405e-08 0.0007 6.9408e-08 0 6.9602e-08 0 6.9605e-08 0.0007 6.9608e-08 0 6.9802e-08 0 6.9805e-08 0.0007 6.9808e-08 0 7.0002e-08 0 7.0005e-08 0.0007 7.0008e-08 0 7.0202e-08 0 7.0205e-08 0.0007 7.0208e-08 0 7.0402e-08 0 7.0405e-08 0.0007 7.0408e-08 0 7.0602e-08 0 7.0605e-08 0.0007 7.0608e-08 0 7.0802e-08 0 7.0805e-08 0.0007 7.0808e-08 0 7.1002e-08 0 7.1005e-08 0.0007 7.1008e-08 0 7.1202e-08 0 7.1205e-08 0.0007 7.1208e-08 0 7.1402e-08 0 7.1405e-08 0.0007 7.1408e-08 0 7.1602e-08 0 7.1605e-08 0.0007 7.1608e-08 0 7.1802e-08 0 7.1805e-08 0.0007 7.1808e-08 0 7.2002e-08 0 7.2005e-08 0.0007 7.2008e-08 0 7.2202e-08 0 7.2205e-08 0.0007 7.2208e-08 0 7.2402e-08 0 7.2405e-08 0.0007 7.2408e-08 0 7.2602e-08 0 7.2605e-08 0.0007 7.2608e-08 0 7.2802e-08 0 7.2805e-08 0.0007 7.2808e-08 0 7.3002e-08 0 7.3005e-08 0.0007 7.3008e-08 0 7.3202e-08 0 7.3205e-08 0.0007 7.3208e-08 0 7.3402e-08 0 7.3405e-08 0.0007 7.3408e-08 0 7.3602e-08 0 7.3605e-08 0.0007 7.3608e-08 0 7.3802e-08 0 7.3805e-08 0.0007 7.3808e-08 0 7.4002e-08 0 7.4005e-08 0.0007 7.4008e-08 0 7.4202e-08 0 7.4205e-08 0.0007 7.4208e-08 0 7.4402e-08 0 7.4405e-08 0.0007 7.4408e-08 0 7.4602e-08 0 7.4605e-08 0.0007 7.4608e-08 0 7.4802e-08 0 7.4805e-08 0.0007 7.4808e-08 0 7.5002e-08 0 7.5005e-08 0.0007 7.5008e-08 0 7.5202e-08 0 7.5205e-08 0.0007 7.5208e-08 0 7.5402e-08 0 7.5405e-08 0.0007 7.5408e-08 0 7.5602e-08 0 7.5605e-08 0.0007 7.5608e-08 0 7.5802e-08 0 7.5805e-08 0.0007 7.5808e-08 0 7.6002e-08 0 7.6005e-08 0.0007 7.6008e-08 0 7.6202e-08 0 7.6205e-08 0.0007 7.6208e-08 0 7.6402e-08 0 7.6405e-08 0.0007 7.6408e-08 0 7.6602e-08 0 7.6605e-08 0.0007 7.6608e-08 0 7.6802e-08 0 7.6805e-08 0.0007 7.6808e-08 0 7.7002e-08 0 7.7005e-08 0.0007 7.7008e-08 0 7.7202e-08 0 7.7205e-08 0.0007 7.7208e-08 0 7.7402e-08 0 7.7405e-08 0.0007 7.7408e-08 0 7.7602e-08 0 7.7605e-08 0.0007 7.7608e-08 0 7.7802e-08 0 7.7805e-08 0.0007 7.7808e-08 0 7.8002e-08 0 7.8005e-08 0.0007 7.8008e-08 0 7.8202e-08 0 7.8205e-08 0.0007 7.8208e-08 0 7.8402e-08 0 7.8405e-08 0.0007 7.8408e-08 0 7.8602e-08 0 7.8605e-08 0.0007 7.8608e-08 0 7.8802e-08 0 7.8805e-08 0.0007 7.8808e-08 0 7.9002e-08 0 7.9005e-08 0.0007 7.9008e-08 0 7.9202e-08 0 7.9205e-08 0.0007 7.9208e-08 0 7.9402e-08 0 7.9405e-08 0.0007 7.9408e-08 0 7.9602e-08 0 7.9605e-08 0.0007 7.9608e-08 0)
BBUF_G1_2_TMP|1 BUF_G1_2_TMP|1 BUF_G1_2_TMP|2 JJMIT AREA=2.5
BBUF_G1_2_TMP|2 BUF_G1_2_TMP|4 BUF_G1_2_TMP|5 JJMIT AREA=2.5
BBUF_G1_2_TMP|3 BUF_G1_2_TMP|7 BUF_G1_2_TMP|8 JJMIT AREA=2.5
BBUF_G1_2_TMP|4 BUF_G1_2_TMP|10 BUF_G1_2_TMP|11 JJMIT AREA=2.5
IBUF_G1_2_TMP|B1 0 BUF_G1_2_TMP|3  PWL(0 0 5e-12 0.000175)
IBUF_G1_2_TMP|B2 0 BUF_G1_2_TMP|6  PWL(0 0 5e-12 0.0002375)
IBUF_G1_2_TMP|B3 0 BUF_G1_2_TMP|9  PWL(0 0 5e-12 0.0002375)
IBUF_G1_2_TMP|B4 0 BUF_G1_2_TMP|12  PWL(0 0 5e-12 0.000175)
LBUF_G1_2_TMP|1 G1_2 BUF_G1_2_TMP|1  2.067833848e-12
LBUF_G1_2_TMP|2 BUF_G1_2_TMP|1 BUF_G1_2_TMP|4  4.135667696e-12
LBUF_G1_2_TMP|3 BUF_G1_2_TMP|4 BUF_G1_2_TMP|7  4.135667696e-12
LBUF_G1_2_TMP|4 BUF_G1_2_TMP|7 BUF_G1_2_TMP|10  4.135667696e-12
LBUF_G1_2_TMP|5 BUF_G1_2_TMP|10 G1_2_TMP  2.067833848e-12
LBUF_G1_2_TMP|P1 BUF_G1_2_TMP|2 0  5e-13
LBUF_G1_2_TMP|P2 BUF_G1_2_TMP|5 0  5e-13
LBUF_G1_2_TMP|P3 BUF_G1_2_TMP|8 0  5e-13
LBUF_G1_2_TMP|P4 BUF_G1_2_TMP|11 0  5e-13
LBUF_G1_2_TMP|B1 BUF_G1_2_TMP|1 BUF_G1_2_TMP|3  2e-12
LBUF_G1_2_TMP|B2 BUF_G1_2_TMP|4 BUF_G1_2_TMP|6  2e-12
LBUF_G1_2_TMP|B3 BUF_G1_2_TMP|7 BUF_G1_2_TMP|9  2e-12
LBUF_G1_2_TMP|B4 BUF_G1_2_TMP|10 BUF_G1_2_TMP|12  2e-12
RBUF_G1_2_TMP|B1 BUF_G1_2_TMP|1 BUF_G1_2_TMP|101  2.7439617672
RBUF_G1_2_TMP|B2 BUF_G1_2_TMP|4 BUF_G1_2_TMP|104  2.7439617672
RBUF_G1_2_TMP|B3 BUF_G1_2_TMP|7 BUF_G1_2_TMP|107  2.7439617672
RBUF_G1_2_TMP|B4 BUF_G1_2_TMP|10 BUF_G1_2_TMP|110  2.7439617672
LBUF_G1_2_TMP|RB1 BUF_G1_2_TMP|101 0  2.050338398468e-12
LBUF_G1_2_TMP|RB2 BUF_G1_2_TMP|104 0  2.050338398468e-12
LBUF_G1_2_TMP|RB3 BUF_G1_2_TMP|107 0  2.050338398468e-12
LBUF_G1_2_TMP|RB4 BUF_G1_2_TMP|110 0  2.050338398468e-12
LBUF_G1_2|1 G1_2_TMP BUF_G1_2|1  2.067833848e-12
LBUF_G1_2|2 BUF_G1_2|1 BUF_G1_2|4  2.067833848e-12
LBUF_G1_2|3 BUF_G1_2|4 BUF_G1_2|6  2.067833848e-12
LBUF_G1_2|4 BUF_G1_2|6 G1_2_BUF  2.067833848e-12
BBUF_IP2_2_TMP|1 BUF_IP2_2_TMP|1 BUF_IP2_2_TMP|2 JJMIT AREA=2.5
BBUF_IP2_2_TMP|2 BUF_IP2_2_TMP|4 BUF_IP2_2_TMP|5 JJMIT AREA=2.5
BBUF_IP2_2_TMP|3 BUF_IP2_2_TMP|7 BUF_IP2_2_TMP|8 JJMIT AREA=2.5
BBUF_IP2_2_TMP|4 BUF_IP2_2_TMP|10 BUF_IP2_2_TMP|11 JJMIT AREA=2.5
IBUF_IP2_2_TMP|B1 0 BUF_IP2_2_TMP|3  PWL(0 0 5e-12 0.000175)
IBUF_IP2_2_TMP|B2 0 BUF_IP2_2_TMP|6  PWL(0 0 5e-12 0.0002375)
IBUF_IP2_2_TMP|B3 0 BUF_IP2_2_TMP|9  PWL(0 0 5e-12 0.0002375)
IBUF_IP2_2_TMP|B4 0 BUF_IP2_2_TMP|12  PWL(0 0 5e-12 0.000175)
LBUF_IP2_2_TMP|1 IP2_2_OUT BUF_IP2_2_TMP|1  2.067833848e-12
LBUF_IP2_2_TMP|2 BUF_IP2_2_TMP|1 BUF_IP2_2_TMP|4  4.135667696e-12
LBUF_IP2_2_TMP|3 BUF_IP2_2_TMP|4 BUF_IP2_2_TMP|7  4.135667696e-12
LBUF_IP2_2_TMP|4 BUF_IP2_2_TMP|7 BUF_IP2_2_TMP|10  4.135667696e-12
LBUF_IP2_2_TMP|5 BUF_IP2_2_TMP|10 IP2_2_TMP  2.067833848e-12
LBUF_IP2_2_TMP|P1 BUF_IP2_2_TMP|2 0  5e-13
LBUF_IP2_2_TMP|P2 BUF_IP2_2_TMP|5 0  5e-13
LBUF_IP2_2_TMP|P3 BUF_IP2_2_TMP|8 0  5e-13
LBUF_IP2_2_TMP|P4 BUF_IP2_2_TMP|11 0  5e-13
LBUF_IP2_2_TMP|B1 BUF_IP2_2_TMP|1 BUF_IP2_2_TMP|3  2e-12
LBUF_IP2_2_TMP|B2 BUF_IP2_2_TMP|4 BUF_IP2_2_TMP|6  2e-12
LBUF_IP2_2_TMP|B3 BUF_IP2_2_TMP|7 BUF_IP2_2_TMP|9  2e-12
LBUF_IP2_2_TMP|B4 BUF_IP2_2_TMP|10 BUF_IP2_2_TMP|12  2e-12
RBUF_IP2_2_TMP|B1 BUF_IP2_2_TMP|1 BUF_IP2_2_TMP|101  2.7439617672
RBUF_IP2_2_TMP|B2 BUF_IP2_2_TMP|4 BUF_IP2_2_TMP|104  2.7439617672
RBUF_IP2_2_TMP|B3 BUF_IP2_2_TMP|7 BUF_IP2_2_TMP|107  2.7439617672
RBUF_IP2_2_TMP|B4 BUF_IP2_2_TMP|10 BUF_IP2_2_TMP|110  2.7439617672
LBUF_IP2_2_TMP|RB1 BUF_IP2_2_TMP|101 0  2.050338398468e-12
LBUF_IP2_2_TMP|RB2 BUF_IP2_2_TMP|104 0  2.050338398468e-12
LBUF_IP2_2_TMP|RB3 BUF_IP2_2_TMP|107 0  2.050338398468e-12
LBUF_IP2_2_TMP|RB4 BUF_IP2_2_TMP|110 0  2.050338398468e-12
LBUF_IP2_2|1 IP2_2_TMP BUF_IP2_2|1  2.067833848e-12
LBUF_IP2_2|2 BUF_IP2_2|1 BUF_IP2_2|4  2.067833848e-12
LBUF_IP2_2|3 BUF_IP2_2|4 BUF_IP2_2|6  2.067833848e-12
LBUF_IP2_2|4 BUF_IP2_2|6 IP2_2_OUT_BUF  2.067833848e-12
L_S2|A1 G1_2_BUF _S2|A1  2.067833848e-12
L_S2|A2 _S2|A1 _S2|A2  4.135667696e-12
L_S2|A3 _S2|A3 _S2|AB  8.271335392e-12
L_S2|B1 IP2_2_OUT_BUF _S2|B1  2.067833848e-12
L_S2|B2 _S2|B1 _S2|B2  4.135667696e-12
L_S2|B3 _S2|B3 _S2|AB  8.271335392e-12
L_S2|T1 T14 _S2|T1  2.067833848e-12
L_S2|T2 _S2|T1 _S2|T2  4.135667696e-12
L_S2|Q2 _S2|ABTQ _S2|Q1  4.135667696e-12
L_S2|Q1 _S2|Q1 S2  2.067833848e-12
IT15|T 0 T15  PWL(0 0 2e-12 0 5e-12 0.0007 8e-12 0 2.02e-10 0 2.05e-10 0.0007 2.08e-10 0 4.02e-10 0 4.05e-10 0.0007 4.08e-10 0 6.02e-10 0 6.05e-10 0.0007 6.08e-10 0 8.02e-10 0 8.05e-10 0.0007 8.08e-10 0 1.002e-09 0 1.005e-09 0.0007 1.008e-09 0 1.202e-09 0 1.205e-09 0.0007 1.208e-09 0 1.402e-09 0 1.405e-09 0.0007 1.408e-09 0 1.602e-09 0 1.605e-09 0.0007 1.608e-09 0 1.802e-09 0 1.805e-09 0.0007 1.808e-09 0 2.002e-09 0 2.005e-09 0.0007 2.008e-09 0 2.202e-09 0 2.205e-09 0.0007 2.208e-09 0 2.402e-09 0 2.405e-09 0.0007 2.408e-09 0 2.602e-09 0 2.605e-09 0.0007 2.608e-09 0 2.802e-09 0 2.805e-09 0.0007 2.808e-09 0 3.002e-09 0 3.005e-09 0.0007 3.008e-09 0 3.202e-09 0 3.205e-09 0.0007 3.208e-09 0 3.402e-09 0 3.405e-09 0.0007 3.408e-09 0 3.602e-09 0 3.605e-09 0.0007 3.608e-09 0 3.802e-09 0 3.805e-09 0.0007 3.808e-09 0 4.002e-09 0 4.005e-09 0.0007 4.008e-09 0 4.202e-09 0 4.205e-09 0.0007 4.208e-09 0 4.402e-09 0 4.405e-09 0.0007 4.408e-09 0 4.602e-09 0 4.605e-09 0.0007 4.608e-09 0 4.802e-09 0 4.805e-09 0.0007 4.808e-09 0 5.002e-09 0 5.005e-09 0.0007 5.008e-09 0 5.202e-09 0 5.205e-09 0.0007 5.208e-09 0 5.402e-09 0 5.405e-09 0.0007 5.408e-09 0 5.602e-09 0 5.605e-09 0.0007 5.608e-09 0 5.802e-09 0 5.805e-09 0.0007 5.808e-09 0 6.002e-09 0 6.005e-09 0.0007 6.008e-09 0 6.202e-09 0 6.205e-09 0.0007 6.208e-09 0 6.402e-09 0 6.405e-09 0.0007 6.408e-09 0 6.602e-09 0 6.605e-09 0.0007 6.608e-09 0 6.802e-09 0 6.805e-09 0.0007 6.808e-09 0 7.002e-09 0 7.005e-09 0.0007 7.008e-09 0 7.202e-09 0 7.205e-09 0.0007 7.208e-09 0 7.402e-09 0 7.405e-09 0.0007 7.408e-09 0 7.602e-09 0 7.605e-09 0.0007 7.608e-09 0 7.802e-09 0 7.805e-09 0.0007 7.808e-09 0 8.002e-09 0 8.005e-09 0.0007 8.008e-09 0 8.202e-09 0 8.205e-09 0.0007 8.208e-09 0 8.402e-09 0 8.405e-09 0.0007 8.408e-09 0 8.602e-09 0 8.605e-09 0.0007 8.608e-09 0 8.802e-09 0 8.805e-09 0.0007 8.808e-09 0 9.002e-09 0 9.005e-09 0.0007 9.008e-09 0 9.202e-09 0 9.205e-09 0.0007 9.208e-09 0 9.402e-09 0 9.405e-09 0.0007 9.408e-09 0 9.602e-09 0 9.605e-09 0.0007 9.608e-09 0 9.802e-09 0 9.805e-09 0.0007 9.808e-09 0 1.0002e-08 0 1.0005e-08 0.0007 1.0008e-08 0 1.0202e-08 0 1.0205e-08 0.0007 1.0208e-08 0 1.0402e-08 0 1.0405e-08 0.0007 1.0408e-08 0 1.0602e-08 0 1.0605e-08 0.0007 1.0608e-08 0 1.0802e-08 0 1.0805e-08 0.0007 1.0808e-08 0 1.1002e-08 0 1.1005e-08 0.0007 1.1008e-08 0 1.1202e-08 0 1.1205e-08 0.0007 1.1208e-08 0 1.1402e-08 0 1.1405e-08 0.0007 1.1408e-08 0 1.1602e-08 0 1.1605e-08 0.0007 1.1608e-08 0 1.1802e-08 0 1.1805e-08 0.0007 1.1808e-08 0 1.2002e-08 0 1.2005e-08 0.0007 1.2008e-08 0 1.2202e-08 0 1.2205e-08 0.0007 1.2208e-08 0 1.2402e-08 0 1.2405e-08 0.0007 1.2408e-08 0 1.2602e-08 0 1.2605e-08 0.0007 1.2608e-08 0 1.2802e-08 0 1.2805e-08 0.0007 1.2808e-08 0 1.3002e-08 0 1.3005e-08 0.0007 1.3008e-08 0 1.3202e-08 0 1.3205e-08 0.0007 1.3208e-08 0 1.3402e-08 0 1.3405e-08 0.0007 1.3408e-08 0 1.3602e-08 0 1.3605e-08 0.0007 1.3608e-08 0 1.3802e-08 0 1.3805e-08 0.0007 1.3808e-08 0 1.4002e-08 0 1.4005e-08 0.0007 1.4008e-08 0 1.4202e-08 0 1.4205e-08 0.0007 1.4208e-08 0 1.4402e-08 0 1.4405e-08 0.0007 1.4408e-08 0 1.4602e-08 0 1.4605e-08 0.0007 1.4608e-08 0 1.4802e-08 0 1.4805e-08 0.0007 1.4808e-08 0 1.5002e-08 0 1.5005e-08 0.0007 1.5008e-08 0 1.5202e-08 0 1.5205e-08 0.0007 1.5208e-08 0 1.5402e-08 0 1.5405e-08 0.0007 1.5408e-08 0 1.5602e-08 0 1.5605e-08 0.0007 1.5608e-08 0 1.5802e-08 0 1.5805e-08 0.0007 1.5808e-08 0 1.6002e-08 0 1.6005e-08 0.0007 1.6008e-08 0 1.6202e-08 0 1.6205e-08 0.0007 1.6208e-08 0 1.6402e-08 0 1.6405e-08 0.0007 1.6408e-08 0 1.6602e-08 0 1.6605e-08 0.0007 1.6608e-08 0 1.6802e-08 0 1.6805e-08 0.0007 1.6808e-08 0 1.7002e-08 0 1.7005e-08 0.0007 1.7008e-08 0 1.7202e-08 0 1.7205e-08 0.0007 1.7208e-08 0 1.7402e-08 0 1.7405e-08 0.0007 1.7408e-08 0 1.7602e-08 0 1.7605e-08 0.0007 1.7608e-08 0 1.7802e-08 0 1.7805e-08 0.0007 1.7808e-08 0 1.8002e-08 0 1.8005e-08 0.0007 1.8008e-08 0 1.8202e-08 0 1.8205e-08 0.0007 1.8208e-08 0 1.8402e-08 0 1.8405e-08 0.0007 1.8408e-08 0 1.8602e-08 0 1.8605e-08 0.0007 1.8608e-08 0 1.8802e-08 0 1.8805e-08 0.0007 1.8808e-08 0 1.9002e-08 0 1.9005e-08 0.0007 1.9008e-08 0 1.9202e-08 0 1.9205e-08 0.0007 1.9208e-08 0 1.9402e-08 0 1.9405e-08 0.0007 1.9408e-08 0 1.9602e-08 0 1.9605e-08 0.0007 1.9608e-08 0 1.9802e-08 0 1.9805e-08 0.0007 1.9808e-08 0 2.0002e-08 0 2.0005e-08 0.0007 2.0008e-08 0 2.0202e-08 0 2.0205e-08 0.0007 2.0208e-08 0 2.0402e-08 0 2.0405e-08 0.0007 2.0408e-08 0 2.0602e-08 0 2.0605e-08 0.0007 2.0608e-08 0 2.0802e-08 0 2.0805e-08 0.0007 2.0808e-08 0 2.1002e-08 0 2.1005e-08 0.0007 2.1008e-08 0 2.1202e-08 0 2.1205e-08 0.0007 2.1208e-08 0 2.1402e-08 0 2.1405e-08 0.0007 2.1408e-08 0 2.1602e-08 0 2.1605e-08 0.0007 2.1608e-08 0 2.1802e-08 0 2.1805e-08 0.0007 2.1808e-08 0 2.2002e-08 0 2.2005e-08 0.0007 2.2008e-08 0 2.2202e-08 0 2.2205e-08 0.0007 2.2208e-08 0 2.2402e-08 0 2.2405e-08 0.0007 2.2408e-08 0 2.2602e-08 0 2.2605e-08 0.0007 2.2608e-08 0 2.2802e-08 0 2.2805e-08 0.0007 2.2808e-08 0 2.3002e-08 0 2.3005e-08 0.0007 2.3008e-08 0 2.3202e-08 0 2.3205e-08 0.0007 2.3208e-08 0 2.3402e-08 0 2.3405e-08 0.0007 2.3408e-08 0 2.3602e-08 0 2.3605e-08 0.0007 2.3608e-08 0 2.3802e-08 0 2.3805e-08 0.0007 2.3808e-08 0 2.4002e-08 0 2.4005e-08 0.0007 2.4008e-08 0 2.4202e-08 0 2.4205e-08 0.0007 2.4208e-08 0 2.4402e-08 0 2.4405e-08 0.0007 2.4408e-08 0 2.4602e-08 0 2.4605e-08 0.0007 2.4608e-08 0 2.4802e-08 0 2.4805e-08 0.0007 2.4808e-08 0 2.5002e-08 0 2.5005e-08 0.0007 2.5008e-08 0 2.5202e-08 0 2.5205e-08 0.0007 2.5208e-08 0 2.5402e-08 0 2.5405e-08 0.0007 2.5408e-08 0 2.5602e-08 0 2.5605e-08 0.0007 2.5608e-08 0 2.5802e-08 0 2.5805e-08 0.0007 2.5808e-08 0 2.6002e-08 0 2.6005e-08 0.0007 2.6008e-08 0 2.6202e-08 0 2.6205e-08 0.0007 2.6208e-08 0 2.6402e-08 0 2.6405e-08 0.0007 2.6408e-08 0 2.6602e-08 0 2.6605e-08 0.0007 2.6608e-08 0 2.6802e-08 0 2.6805e-08 0.0007 2.6808e-08 0 2.7002e-08 0 2.7005e-08 0.0007 2.7008e-08 0 2.7202e-08 0 2.7205e-08 0.0007 2.7208e-08 0 2.7402e-08 0 2.7405e-08 0.0007 2.7408e-08 0 2.7602e-08 0 2.7605e-08 0.0007 2.7608e-08 0 2.7802e-08 0 2.7805e-08 0.0007 2.7808e-08 0 2.8002e-08 0 2.8005e-08 0.0007 2.8008e-08 0 2.8202e-08 0 2.8205e-08 0.0007 2.8208e-08 0 2.8402e-08 0 2.8405e-08 0.0007 2.8408e-08 0 2.8602e-08 0 2.8605e-08 0.0007 2.8608e-08 0 2.8802e-08 0 2.8805e-08 0.0007 2.8808e-08 0 2.9002e-08 0 2.9005e-08 0.0007 2.9008e-08 0 2.9202e-08 0 2.9205e-08 0.0007 2.9208e-08 0 2.9402e-08 0 2.9405e-08 0.0007 2.9408e-08 0 2.9602e-08 0 2.9605e-08 0.0007 2.9608e-08 0 2.9802e-08 0 2.9805e-08 0.0007 2.9808e-08 0 3.0002e-08 0 3.0005e-08 0.0007 3.0008e-08 0 3.0202e-08 0 3.0205e-08 0.0007 3.0208e-08 0 3.0402e-08 0 3.0405e-08 0.0007 3.0408e-08 0 3.0602e-08 0 3.0605e-08 0.0007 3.0608e-08 0 3.0802e-08 0 3.0805e-08 0.0007 3.0808e-08 0 3.1002e-08 0 3.1005e-08 0.0007 3.1008e-08 0 3.1202e-08 0 3.1205e-08 0.0007 3.1208e-08 0 3.1402e-08 0 3.1405e-08 0.0007 3.1408e-08 0 3.1602e-08 0 3.1605e-08 0.0007 3.1608e-08 0 3.1802e-08 0 3.1805e-08 0.0007 3.1808e-08 0 3.2002e-08 0 3.2005e-08 0.0007 3.2008e-08 0 3.2202e-08 0 3.2205e-08 0.0007 3.2208e-08 0 3.2402e-08 0 3.2405e-08 0.0007 3.2408e-08 0 3.2602e-08 0 3.2605e-08 0.0007 3.2608e-08 0 3.2802e-08 0 3.2805e-08 0.0007 3.2808e-08 0 3.3002e-08 0 3.3005e-08 0.0007 3.3008e-08 0 3.3202e-08 0 3.3205e-08 0.0007 3.3208e-08 0 3.3402e-08 0 3.3405e-08 0.0007 3.3408e-08 0 3.3602e-08 0 3.3605e-08 0.0007 3.3608e-08 0 3.3802e-08 0 3.3805e-08 0.0007 3.3808e-08 0 3.4002e-08 0 3.4005e-08 0.0007 3.4008e-08 0 3.4202e-08 0 3.4205e-08 0.0007 3.4208e-08 0 3.4402e-08 0 3.4405e-08 0.0007 3.4408e-08 0 3.4602e-08 0 3.4605e-08 0.0007 3.4608e-08 0 3.4802e-08 0 3.4805e-08 0.0007 3.4808e-08 0 3.5002e-08 0 3.5005e-08 0.0007 3.5008e-08 0 3.5202e-08 0 3.5205e-08 0.0007 3.5208e-08 0 3.5402e-08 0 3.5405e-08 0.0007 3.5408e-08 0 3.5602e-08 0 3.5605e-08 0.0007 3.5608e-08 0 3.5802e-08 0 3.5805e-08 0.0007 3.5808e-08 0 3.6002e-08 0 3.6005e-08 0.0007 3.6008e-08 0 3.6202e-08 0 3.6205e-08 0.0007 3.6208e-08 0 3.6402e-08 0 3.6405e-08 0.0007 3.6408e-08 0 3.6602e-08 0 3.6605e-08 0.0007 3.6608e-08 0 3.6802e-08 0 3.6805e-08 0.0007 3.6808e-08 0 3.7002e-08 0 3.7005e-08 0.0007 3.7008e-08 0 3.7202e-08 0 3.7205e-08 0.0007 3.7208e-08 0 3.7402e-08 0 3.7405e-08 0.0007 3.7408e-08 0 3.7602e-08 0 3.7605e-08 0.0007 3.7608e-08 0 3.7802e-08 0 3.7805e-08 0.0007 3.7808e-08 0 3.8002e-08 0 3.8005e-08 0.0007 3.8008e-08 0 3.8202e-08 0 3.8205e-08 0.0007 3.8208e-08 0 3.8402e-08 0 3.8405e-08 0.0007 3.8408e-08 0 3.8602e-08 0 3.8605e-08 0.0007 3.8608e-08 0 3.8802e-08 0 3.8805e-08 0.0007 3.8808e-08 0 3.9002e-08 0 3.9005e-08 0.0007 3.9008e-08 0 3.9202e-08 0 3.9205e-08 0.0007 3.9208e-08 0 3.9402e-08 0 3.9405e-08 0.0007 3.9408e-08 0 3.9602e-08 0 3.9605e-08 0.0007 3.9608e-08 0 3.9802e-08 0 3.9805e-08 0.0007 3.9808e-08 0 4.0002e-08 0 4.0005e-08 0.0007 4.0008e-08 0 4.0202e-08 0 4.0205e-08 0.0007 4.0208e-08 0 4.0402e-08 0 4.0405e-08 0.0007 4.0408e-08 0 4.0602e-08 0 4.0605e-08 0.0007 4.0608e-08 0 4.0802e-08 0 4.0805e-08 0.0007 4.0808e-08 0 4.1002e-08 0 4.1005e-08 0.0007 4.1008e-08 0 4.1202e-08 0 4.1205e-08 0.0007 4.1208e-08 0 4.1402e-08 0 4.1405e-08 0.0007 4.1408e-08 0 4.1602e-08 0 4.1605e-08 0.0007 4.1608e-08 0 4.1802e-08 0 4.1805e-08 0.0007 4.1808e-08 0 4.2002e-08 0 4.2005e-08 0.0007 4.2008e-08 0 4.2202e-08 0 4.2205e-08 0.0007 4.2208e-08 0 4.2402e-08 0 4.2405e-08 0.0007 4.2408e-08 0 4.2602e-08 0 4.2605e-08 0.0007 4.2608e-08 0 4.2802e-08 0 4.2805e-08 0.0007 4.2808e-08 0 4.3002e-08 0 4.3005e-08 0.0007 4.3008e-08 0 4.3202e-08 0 4.3205e-08 0.0007 4.3208e-08 0 4.3402e-08 0 4.3405e-08 0.0007 4.3408e-08 0 4.3602e-08 0 4.3605e-08 0.0007 4.3608e-08 0 4.3802e-08 0 4.3805e-08 0.0007 4.3808e-08 0 4.4002e-08 0 4.4005e-08 0.0007 4.4008e-08 0 4.4202e-08 0 4.4205e-08 0.0007 4.4208e-08 0 4.4402e-08 0 4.4405e-08 0.0007 4.4408e-08 0 4.4602e-08 0 4.4605e-08 0.0007 4.4608e-08 0 4.4802e-08 0 4.4805e-08 0.0007 4.4808e-08 0 4.5002e-08 0 4.5005e-08 0.0007 4.5008e-08 0 4.5202e-08 0 4.5205e-08 0.0007 4.5208e-08 0 4.5402e-08 0 4.5405e-08 0.0007 4.5408e-08 0 4.5602e-08 0 4.5605e-08 0.0007 4.5608e-08 0 4.5802e-08 0 4.5805e-08 0.0007 4.5808e-08 0 4.6002e-08 0 4.6005e-08 0.0007 4.6008e-08 0 4.6202e-08 0 4.6205e-08 0.0007 4.6208e-08 0 4.6402e-08 0 4.6405e-08 0.0007 4.6408e-08 0 4.6602e-08 0 4.6605e-08 0.0007 4.6608e-08 0 4.6802e-08 0 4.6805e-08 0.0007 4.6808e-08 0 4.7002e-08 0 4.7005e-08 0.0007 4.7008e-08 0 4.7202e-08 0 4.7205e-08 0.0007 4.7208e-08 0 4.7402e-08 0 4.7405e-08 0.0007 4.7408e-08 0 4.7602e-08 0 4.7605e-08 0.0007 4.7608e-08 0 4.7802e-08 0 4.7805e-08 0.0007 4.7808e-08 0 4.8002e-08 0 4.8005e-08 0.0007 4.8008e-08 0 4.8202e-08 0 4.8205e-08 0.0007 4.8208e-08 0 4.8402e-08 0 4.8405e-08 0.0007 4.8408e-08 0 4.8602e-08 0 4.8605e-08 0.0007 4.8608e-08 0 4.8802e-08 0 4.8805e-08 0.0007 4.8808e-08 0 4.9002e-08 0 4.9005e-08 0.0007 4.9008e-08 0 4.9202e-08 0 4.9205e-08 0.0007 4.9208e-08 0 4.9402e-08 0 4.9405e-08 0.0007 4.9408e-08 0 4.9602e-08 0 4.9605e-08 0.0007 4.9608e-08 0 4.9802e-08 0 4.9805e-08 0.0007 4.9808e-08 0 5.0002e-08 0 5.0005e-08 0.0007 5.0008e-08 0 5.0202e-08 0 5.0205e-08 0.0007 5.0208e-08 0 5.0402e-08 0 5.0405e-08 0.0007 5.0408e-08 0 5.0602e-08 0 5.0605e-08 0.0007 5.0608e-08 0 5.0802e-08 0 5.0805e-08 0.0007 5.0808e-08 0 5.1002e-08 0 5.1005e-08 0.0007 5.1008e-08 0 5.1202e-08 0 5.1205e-08 0.0007 5.1208e-08 0 5.1402e-08 0 5.1405e-08 0.0007 5.1408e-08 0 5.1602e-08 0 5.1605e-08 0.0007 5.1608e-08 0 5.1802e-08 0 5.1805e-08 0.0007 5.1808e-08 0 5.2002e-08 0 5.2005e-08 0.0007 5.2008e-08 0 5.2202e-08 0 5.2205e-08 0.0007 5.2208e-08 0 5.2402e-08 0 5.2405e-08 0.0007 5.2408e-08 0 5.2602e-08 0 5.2605e-08 0.0007 5.2608e-08 0 5.2802e-08 0 5.2805e-08 0.0007 5.2808e-08 0 5.3002e-08 0 5.3005e-08 0.0007 5.3008e-08 0 5.3202e-08 0 5.3205e-08 0.0007 5.3208e-08 0 5.3402e-08 0 5.3405e-08 0.0007 5.3408e-08 0 5.3602e-08 0 5.3605e-08 0.0007 5.3608e-08 0 5.3802e-08 0 5.3805e-08 0.0007 5.3808e-08 0 5.4002e-08 0 5.4005e-08 0.0007 5.4008e-08 0 5.4202e-08 0 5.4205e-08 0.0007 5.4208e-08 0 5.4402e-08 0 5.4405e-08 0.0007 5.4408e-08 0 5.4602e-08 0 5.4605e-08 0.0007 5.4608e-08 0 5.4802e-08 0 5.4805e-08 0.0007 5.4808e-08 0 5.5002e-08 0 5.5005e-08 0.0007 5.5008e-08 0 5.5202e-08 0 5.5205e-08 0.0007 5.5208e-08 0 5.5402e-08 0 5.5405e-08 0.0007 5.5408e-08 0 5.5602e-08 0 5.5605e-08 0.0007 5.5608e-08 0 5.5802e-08 0 5.5805e-08 0.0007 5.5808e-08 0 5.6002e-08 0 5.6005e-08 0.0007 5.6008e-08 0 5.6202e-08 0 5.6205e-08 0.0007 5.6208e-08 0 5.6402e-08 0 5.6405e-08 0.0007 5.6408e-08 0 5.6602e-08 0 5.6605e-08 0.0007 5.6608e-08 0 5.6802e-08 0 5.6805e-08 0.0007 5.6808e-08 0 5.7002e-08 0 5.7005e-08 0.0007 5.7008e-08 0 5.7202e-08 0 5.7205e-08 0.0007 5.7208e-08 0 5.7402e-08 0 5.7405e-08 0.0007 5.7408e-08 0 5.7602e-08 0 5.7605e-08 0.0007 5.7608e-08 0 5.7802e-08 0 5.7805e-08 0.0007 5.7808e-08 0 5.8002e-08 0 5.8005e-08 0.0007 5.8008e-08 0 5.8202e-08 0 5.8205e-08 0.0007 5.8208e-08 0 5.8402e-08 0 5.8405e-08 0.0007 5.8408e-08 0 5.8602e-08 0 5.8605e-08 0.0007 5.8608e-08 0 5.8802e-08 0 5.8805e-08 0.0007 5.8808e-08 0 5.9002e-08 0 5.9005e-08 0.0007 5.9008e-08 0 5.9202e-08 0 5.9205e-08 0.0007 5.9208e-08 0 5.9402e-08 0 5.9405e-08 0.0007 5.9408e-08 0 5.9602e-08 0 5.9605e-08 0.0007 5.9608e-08 0 5.9802e-08 0 5.9805e-08 0.0007 5.9808e-08 0 6.0002e-08 0 6.0005e-08 0.0007 6.0008e-08 0 6.0202e-08 0 6.0205e-08 0.0007 6.0208e-08 0 6.0402e-08 0 6.0405e-08 0.0007 6.0408e-08 0 6.0602e-08 0 6.0605e-08 0.0007 6.0608e-08 0 6.0802e-08 0 6.0805e-08 0.0007 6.0808e-08 0 6.1002e-08 0 6.1005e-08 0.0007 6.1008e-08 0 6.1202e-08 0 6.1205e-08 0.0007 6.1208e-08 0 6.1402e-08 0 6.1405e-08 0.0007 6.1408e-08 0 6.1602e-08 0 6.1605e-08 0.0007 6.1608e-08 0 6.1802e-08 0 6.1805e-08 0.0007 6.1808e-08 0 6.2002e-08 0 6.2005e-08 0.0007 6.2008e-08 0 6.2202e-08 0 6.2205e-08 0.0007 6.2208e-08 0 6.2402e-08 0 6.2405e-08 0.0007 6.2408e-08 0 6.2602e-08 0 6.2605e-08 0.0007 6.2608e-08 0 6.2802e-08 0 6.2805e-08 0.0007 6.2808e-08 0 6.3002e-08 0 6.3005e-08 0.0007 6.3008e-08 0 6.3202e-08 0 6.3205e-08 0.0007 6.3208e-08 0 6.3402e-08 0 6.3405e-08 0.0007 6.3408e-08 0 6.3602e-08 0 6.3605e-08 0.0007 6.3608e-08 0 6.3802e-08 0 6.3805e-08 0.0007 6.3808e-08 0 6.4002e-08 0 6.4005e-08 0.0007 6.4008e-08 0 6.4202e-08 0 6.4205e-08 0.0007 6.4208e-08 0 6.4402e-08 0 6.4405e-08 0.0007 6.4408e-08 0 6.4602e-08 0 6.4605e-08 0.0007 6.4608e-08 0 6.4802e-08 0 6.4805e-08 0.0007 6.4808e-08 0 6.5002e-08 0 6.5005e-08 0.0007 6.5008e-08 0 6.5202e-08 0 6.5205e-08 0.0007 6.5208e-08 0 6.5402e-08 0 6.5405e-08 0.0007 6.5408e-08 0 6.5602e-08 0 6.5605e-08 0.0007 6.5608e-08 0 6.5802e-08 0 6.5805e-08 0.0007 6.5808e-08 0 6.6002e-08 0 6.6005e-08 0.0007 6.6008e-08 0 6.6202e-08 0 6.6205e-08 0.0007 6.6208e-08 0 6.6402e-08 0 6.6405e-08 0.0007 6.6408e-08 0 6.6602e-08 0 6.6605e-08 0.0007 6.6608e-08 0 6.6802e-08 0 6.6805e-08 0.0007 6.6808e-08 0 6.7002e-08 0 6.7005e-08 0.0007 6.7008e-08 0 6.7202e-08 0 6.7205e-08 0.0007 6.7208e-08 0 6.7402e-08 0 6.7405e-08 0.0007 6.7408e-08 0 6.7602e-08 0 6.7605e-08 0.0007 6.7608e-08 0 6.7802e-08 0 6.7805e-08 0.0007 6.7808e-08 0 6.8002e-08 0 6.8005e-08 0.0007 6.8008e-08 0 6.8202e-08 0 6.8205e-08 0.0007 6.8208e-08 0 6.8402e-08 0 6.8405e-08 0.0007 6.8408e-08 0 6.8602e-08 0 6.8605e-08 0.0007 6.8608e-08 0 6.8802e-08 0 6.8805e-08 0.0007 6.8808e-08 0 6.9002e-08 0 6.9005e-08 0.0007 6.9008e-08 0 6.9202e-08 0 6.9205e-08 0.0007 6.9208e-08 0 6.9402e-08 0 6.9405e-08 0.0007 6.9408e-08 0 6.9602e-08 0 6.9605e-08 0.0007 6.9608e-08 0 6.9802e-08 0 6.9805e-08 0.0007 6.9808e-08 0 7.0002e-08 0 7.0005e-08 0.0007 7.0008e-08 0 7.0202e-08 0 7.0205e-08 0.0007 7.0208e-08 0 7.0402e-08 0 7.0405e-08 0.0007 7.0408e-08 0 7.0602e-08 0 7.0605e-08 0.0007 7.0608e-08 0 7.0802e-08 0 7.0805e-08 0.0007 7.0808e-08 0 7.1002e-08 0 7.1005e-08 0.0007 7.1008e-08 0 7.1202e-08 0 7.1205e-08 0.0007 7.1208e-08 0 7.1402e-08 0 7.1405e-08 0.0007 7.1408e-08 0 7.1602e-08 0 7.1605e-08 0.0007 7.1608e-08 0 7.1802e-08 0 7.1805e-08 0.0007 7.1808e-08 0 7.2002e-08 0 7.2005e-08 0.0007 7.2008e-08 0 7.2202e-08 0 7.2205e-08 0.0007 7.2208e-08 0 7.2402e-08 0 7.2405e-08 0.0007 7.2408e-08 0 7.2602e-08 0 7.2605e-08 0.0007 7.2608e-08 0 7.2802e-08 0 7.2805e-08 0.0007 7.2808e-08 0 7.3002e-08 0 7.3005e-08 0.0007 7.3008e-08 0 7.3202e-08 0 7.3205e-08 0.0007 7.3208e-08 0 7.3402e-08 0 7.3405e-08 0.0007 7.3408e-08 0 7.3602e-08 0 7.3605e-08 0.0007 7.3608e-08 0 7.3802e-08 0 7.3805e-08 0.0007 7.3808e-08 0 7.4002e-08 0 7.4005e-08 0.0007 7.4008e-08 0 7.4202e-08 0 7.4205e-08 0.0007 7.4208e-08 0 7.4402e-08 0 7.4405e-08 0.0007 7.4408e-08 0 7.4602e-08 0 7.4605e-08 0.0007 7.4608e-08 0 7.4802e-08 0 7.4805e-08 0.0007 7.4808e-08 0 7.5002e-08 0 7.5005e-08 0.0007 7.5008e-08 0 7.5202e-08 0 7.5205e-08 0.0007 7.5208e-08 0 7.5402e-08 0 7.5405e-08 0.0007 7.5408e-08 0 7.5602e-08 0 7.5605e-08 0.0007 7.5608e-08 0 7.5802e-08 0 7.5805e-08 0.0007 7.5808e-08 0 7.6002e-08 0 7.6005e-08 0.0007 7.6008e-08 0 7.6202e-08 0 7.6205e-08 0.0007 7.6208e-08 0 7.6402e-08 0 7.6405e-08 0.0007 7.6408e-08 0 7.6602e-08 0 7.6605e-08 0.0007 7.6608e-08 0 7.6802e-08 0 7.6805e-08 0.0007 7.6808e-08 0 7.7002e-08 0 7.7005e-08 0.0007 7.7008e-08 0 7.7202e-08 0 7.7205e-08 0.0007 7.7208e-08 0 7.7402e-08 0 7.7405e-08 0.0007 7.7408e-08 0 7.7602e-08 0 7.7605e-08 0.0007 7.7608e-08 0 7.7802e-08 0 7.7805e-08 0.0007 7.7808e-08 0 7.8002e-08 0 7.8005e-08 0.0007 7.8008e-08 0 7.8202e-08 0 7.8205e-08 0.0007 7.8208e-08 0 7.8402e-08 0 7.8405e-08 0.0007 7.8408e-08 0 7.8602e-08 0 7.8605e-08 0.0007 7.8608e-08 0 7.8802e-08 0 7.8805e-08 0.0007 7.8808e-08 0 7.9002e-08 0 7.9005e-08 0.0007 7.9008e-08 0 7.9202e-08 0 7.9205e-08 0.0007 7.9208e-08 0 7.9402e-08 0 7.9405e-08 0.0007 7.9408e-08 0 7.9602e-08 0 7.9605e-08 0.0007 7.9608e-08 0)
BBUF_G2_2_TMP|1 BUF_G2_2_TMP|1 BUF_G2_2_TMP|2 JJMIT AREA=2.5
BBUF_G2_2_TMP|2 BUF_G2_2_TMP|4 BUF_G2_2_TMP|5 JJMIT AREA=2.5
BBUF_G2_2_TMP|3 BUF_G2_2_TMP|7 BUF_G2_2_TMP|8 JJMIT AREA=2.5
BBUF_G2_2_TMP|4 BUF_G2_2_TMP|10 BUF_G2_2_TMP|11 JJMIT AREA=2.5
IBUF_G2_2_TMP|B1 0 BUF_G2_2_TMP|3  PWL(0 0 5e-12 0.000175)
IBUF_G2_2_TMP|B2 0 BUF_G2_2_TMP|6  PWL(0 0 5e-12 0.0002375)
IBUF_G2_2_TMP|B3 0 BUF_G2_2_TMP|9  PWL(0 0 5e-12 0.0002375)
IBUF_G2_2_TMP|B4 0 BUF_G2_2_TMP|12  PWL(0 0 5e-12 0.000175)
LBUF_G2_2_TMP|1 G2_2 BUF_G2_2_TMP|1  2.067833848e-12
LBUF_G2_2_TMP|2 BUF_G2_2_TMP|1 BUF_G2_2_TMP|4  4.135667696e-12
LBUF_G2_2_TMP|3 BUF_G2_2_TMP|4 BUF_G2_2_TMP|7  4.135667696e-12
LBUF_G2_2_TMP|4 BUF_G2_2_TMP|7 BUF_G2_2_TMP|10  4.135667696e-12
LBUF_G2_2_TMP|5 BUF_G2_2_TMP|10 G2_2_TMP  2.067833848e-12
LBUF_G2_2_TMP|P1 BUF_G2_2_TMP|2 0  5e-13
LBUF_G2_2_TMP|P2 BUF_G2_2_TMP|5 0  5e-13
LBUF_G2_2_TMP|P3 BUF_G2_2_TMP|8 0  5e-13
LBUF_G2_2_TMP|P4 BUF_G2_2_TMP|11 0  5e-13
LBUF_G2_2_TMP|B1 BUF_G2_2_TMP|1 BUF_G2_2_TMP|3  2e-12
LBUF_G2_2_TMP|B2 BUF_G2_2_TMP|4 BUF_G2_2_TMP|6  2e-12
LBUF_G2_2_TMP|B3 BUF_G2_2_TMP|7 BUF_G2_2_TMP|9  2e-12
LBUF_G2_2_TMP|B4 BUF_G2_2_TMP|10 BUF_G2_2_TMP|12  2e-12
RBUF_G2_2_TMP|B1 BUF_G2_2_TMP|1 BUF_G2_2_TMP|101  2.7439617672
RBUF_G2_2_TMP|B2 BUF_G2_2_TMP|4 BUF_G2_2_TMP|104  2.7439617672
RBUF_G2_2_TMP|B3 BUF_G2_2_TMP|7 BUF_G2_2_TMP|107  2.7439617672
RBUF_G2_2_TMP|B4 BUF_G2_2_TMP|10 BUF_G2_2_TMP|110  2.7439617672
LBUF_G2_2_TMP|RB1 BUF_G2_2_TMP|101 0  2.050338398468e-12
LBUF_G2_2_TMP|RB2 BUF_G2_2_TMP|104 0  2.050338398468e-12
LBUF_G2_2_TMP|RB3 BUF_G2_2_TMP|107 0  2.050338398468e-12
LBUF_G2_2_TMP|RB4 BUF_G2_2_TMP|110 0  2.050338398468e-12
LBUF_G2_2|1 G2_2_TMP BUF_G2_2|1  2.067833848e-12
LBUF_G2_2|2 BUF_G2_2|1 BUF_G2_2|4  2.067833848e-12
LBUF_G2_2|3 BUF_G2_2|4 BUF_G2_2|6  2.067833848e-12
LBUF_G2_2|4 BUF_G2_2|6 G2_2_BUF  2.067833848e-12
L_S3|A1 G2_2_TMP _S3|A1  2.067833848e-12
L_S3|A2 _S3|A1 _S3|A2  4.135667696e-12
L_S3|A3 _S3|A3 _S3|AB  8.271335392e-12
L_S3|B1 IP3_2_OUT _S3|B1  2.067833848e-12
L_S3|B2 _S3|B1 _S3|B2  4.135667696e-12
L_S3|B3 _S3|B3 _S3|AB  8.271335392e-12
L_S3|T1 T15 _S3|T1  2.067833848e-12
L_S3|T2 _S3|T1 _S3|T2  4.135667696e-12
L_S3|Q2 _S3|ABTQ _S3|Q1  4.135667696e-12
L_S3|Q1 _S3|Q1 S3  2.067833848e-12
IT16|T 0 T16  PWL(0 0 2e-12 0 5e-12 0.0007 8e-12 0 2.02e-10 0 2.05e-10 0.0007 2.08e-10 0 4.02e-10 0 4.05e-10 0.0007 4.08e-10 0 6.02e-10 0 6.05e-10 0.0007 6.08e-10 0 8.02e-10 0 8.05e-10 0.0007 8.08e-10 0 1.002e-09 0 1.005e-09 0.0007 1.008e-09 0 1.202e-09 0 1.205e-09 0.0007 1.208e-09 0 1.402e-09 0 1.405e-09 0.0007 1.408e-09 0 1.602e-09 0 1.605e-09 0.0007 1.608e-09 0 1.802e-09 0 1.805e-09 0.0007 1.808e-09 0 2.002e-09 0 2.005e-09 0.0007 2.008e-09 0 2.202e-09 0 2.205e-09 0.0007 2.208e-09 0 2.402e-09 0 2.405e-09 0.0007 2.408e-09 0 2.602e-09 0 2.605e-09 0.0007 2.608e-09 0 2.802e-09 0 2.805e-09 0.0007 2.808e-09 0 3.002e-09 0 3.005e-09 0.0007 3.008e-09 0 3.202e-09 0 3.205e-09 0.0007 3.208e-09 0 3.402e-09 0 3.405e-09 0.0007 3.408e-09 0 3.602e-09 0 3.605e-09 0.0007 3.608e-09 0 3.802e-09 0 3.805e-09 0.0007 3.808e-09 0 4.002e-09 0 4.005e-09 0.0007 4.008e-09 0 4.202e-09 0 4.205e-09 0.0007 4.208e-09 0 4.402e-09 0 4.405e-09 0.0007 4.408e-09 0 4.602e-09 0 4.605e-09 0.0007 4.608e-09 0 4.802e-09 0 4.805e-09 0.0007 4.808e-09 0 5.002e-09 0 5.005e-09 0.0007 5.008e-09 0 5.202e-09 0 5.205e-09 0.0007 5.208e-09 0 5.402e-09 0 5.405e-09 0.0007 5.408e-09 0 5.602e-09 0 5.605e-09 0.0007 5.608e-09 0 5.802e-09 0 5.805e-09 0.0007 5.808e-09 0 6.002e-09 0 6.005e-09 0.0007 6.008e-09 0 6.202e-09 0 6.205e-09 0.0007 6.208e-09 0 6.402e-09 0 6.405e-09 0.0007 6.408e-09 0 6.602e-09 0 6.605e-09 0.0007 6.608e-09 0 6.802e-09 0 6.805e-09 0.0007 6.808e-09 0 7.002e-09 0 7.005e-09 0.0007 7.008e-09 0 7.202e-09 0 7.205e-09 0.0007 7.208e-09 0 7.402e-09 0 7.405e-09 0.0007 7.408e-09 0 7.602e-09 0 7.605e-09 0.0007 7.608e-09 0 7.802e-09 0 7.805e-09 0.0007 7.808e-09 0 8.002e-09 0 8.005e-09 0.0007 8.008e-09 0 8.202e-09 0 8.205e-09 0.0007 8.208e-09 0 8.402e-09 0 8.405e-09 0.0007 8.408e-09 0 8.602e-09 0 8.605e-09 0.0007 8.608e-09 0 8.802e-09 0 8.805e-09 0.0007 8.808e-09 0 9.002e-09 0 9.005e-09 0.0007 9.008e-09 0 9.202e-09 0 9.205e-09 0.0007 9.208e-09 0 9.402e-09 0 9.405e-09 0.0007 9.408e-09 0 9.602e-09 0 9.605e-09 0.0007 9.608e-09 0 9.802e-09 0 9.805e-09 0.0007 9.808e-09 0 1.0002e-08 0 1.0005e-08 0.0007 1.0008e-08 0 1.0202e-08 0 1.0205e-08 0.0007 1.0208e-08 0 1.0402e-08 0 1.0405e-08 0.0007 1.0408e-08 0 1.0602e-08 0 1.0605e-08 0.0007 1.0608e-08 0 1.0802e-08 0 1.0805e-08 0.0007 1.0808e-08 0 1.1002e-08 0 1.1005e-08 0.0007 1.1008e-08 0 1.1202e-08 0 1.1205e-08 0.0007 1.1208e-08 0 1.1402e-08 0 1.1405e-08 0.0007 1.1408e-08 0 1.1602e-08 0 1.1605e-08 0.0007 1.1608e-08 0 1.1802e-08 0 1.1805e-08 0.0007 1.1808e-08 0 1.2002e-08 0 1.2005e-08 0.0007 1.2008e-08 0 1.2202e-08 0 1.2205e-08 0.0007 1.2208e-08 0 1.2402e-08 0 1.2405e-08 0.0007 1.2408e-08 0 1.2602e-08 0 1.2605e-08 0.0007 1.2608e-08 0 1.2802e-08 0 1.2805e-08 0.0007 1.2808e-08 0 1.3002e-08 0 1.3005e-08 0.0007 1.3008e-08 0 1.3202e-08 0 1.3205e-08 0.0007 1.3208e-08 0 1.3402e-08 0 1.3405e-08 0.0007 1.3408e-08 0 1.3602e-08 0 1.3605e-08 0.0007 1.3608e-08 0 1.3802e-08 0 1.3805e-08 0.0007 1.3808e-08 0 1.4002e-08 0 1.4005e-08 0.0007 1.4008e-08 0 1.4202e-08 0 1.4205e-08 0.0007 1.4208e-08 0 1.4402e-08 0 1.4405e-08 0.0007 1.4408e-08 0 1.4602e-08 0 1.4605e-08 0.0007 1.4608e-08 0 1.4802e-08 0 1.4805e-08 0.0007 1.4808e-08 0 1.5002e-08 0 1.5005e-08 0.0007 1.5008e-08 0 1.5202e-08 0 1.5205e-08 0.0007 1.5208e-08 0 1.5402e-08 0 1.5405e-08 0.0007 1.5408e-08 0 1.5602e-08 0 1.5605e-08 0.0007 1.5608e-08 0 1.5802e-08 0 1.5805e-08 0.0007 1.5808e-08 0 1.6002e-08 0 1.6005e-08 0.0007 1.6008e-08 0 1.6202e-08 0 1.6205e-08 0.0007 1.6208e-08 0 1.6402e-08 0 1.6405e-08 0.0007 1.6408e-08 0 1.6602e-08 0 1.6605e-08 0.0007 1.6608e-08 0 1.6802e-08 0 1.6805e-08 0.0007 1.6808e-08 0 1.7002e-08 0 1.7005e-08 0.0007 1.7008e-08 0 1.7202e-08 0 1.7205e-08 0.0007 1.7208e-08 0 1.7402e-08 0 1.7405e-08 0.0007 1.7408e-08 0 1.7602e-08 0 1.7605e-08 0.0007 1.7608e-08 0 1.7802e-08 0 1.7805e-08 0.0007 1.7808e-08 0 1.8002e-08 0 1.8005e-08 0.0007 1.8008e-08 0 1.8202e-08 0 1.8205e-08 0.0007 1.8208e-08 0 1.8402e-08 0 1.8405e-08 0.0007 1.8408e-08 0 1.8602e-08 0 1.8605e-08 0.0007 1.8608e-08 0 1.8802e-08 0 1.8805e-08 0.0007 1.8808e-08 0 1.9002e-08 0 1.9005e-08 0.0007 1.9008e-08 0 1.9202e-08 0 1.9205e-08 0.0007 1.9208e-08 0 1.9402e-08 0 1.9405e-08 0.0007 1.9408e-08 0 1.9602e-08 0 1.9605e-08 0.0007 1.9608e-08 0 1.9802e-08 0 1.9805e-08 0.0007 1.9808e-08 0 2.0002e-08 0 2.0005e-08 0.0007 2.0008e-08 0 2.0202e-08 0 2.0205e-08 0.0007 2.0208e-08 0 2.0402e-08 0 2.0405e-08 0.0007 2.0408e-08 0 2.0602e-08 0 2.0605e-08 0.0007 2.0608e-08 0 2.0802e-08 0 2.0805e-08 0.0007 2.0808e-08 0 2.1002e-08 0 2.1005e-08 0.0007 2.1008e-08 0 2.1202e-08 0 2.1205e-08 0.0007 2.1208e-08 0 2.1402e-08 0 2.1405e-08 0.0007 2.1408e-08 0 2.1602e-08 0 2.1605e-08 0.0007 2.1608e-08 0 2.1802e-08 0 2.1805e-08 0.0007 2.1808e-08 0 2.2002e-08 0 2.2005e-08 0.0007 2.2008e-08 0 2.2202e-08 0 2.2205e-08 0.0007 2.2208e-08 0 2.2402e-08 0 2.2405e-08 0.0007 2.2408e-08 0 2.2602e-08 0 2.2605e-08 0.0007 2.2608e-08 0 2.2802e-08 0 2.2805e-08 0.0007 2.2808e-08 0 2.3002e-08 0 2.3005e-08 0.0007 2.3008e-08 0 2.3202e-08 0 2.3205e-08 0.0007 2.3208e-08 0 2.3402e-08 0 2.3405e-08 0.0007 2.3408e-08 0 2.3602e-08 0 2.3605e-08 0.0007 2.3608e-08 0 2.3802e-08 0 2.3805e-08 0.0007 2.3808e-08 0 2.4002e-08 0 2.4005e-08 0.0007 2.4008e-08 0 2.4202e-08 0 2.4205e-08 0.0007 2.4208e-08 0 2.4402e-08 0 2.4405e-08 0.0007 2.4408e-08 0 2.4602e-08 0 2.4605e-08 0.0007 2.4608e-08 0 2.4802e-08 0 2.4805e-08 0.0007 2.4808e-08 0 2.5002e-08 0 2.5005e-08 0.0007 2.5008e-08 0 2.5202e-08 0 2.5205e-08 0.0007 2.5208e-08 0 2.5402e-08 0 2.5405e-08 0.0007 2.5408e-08 0 2.5602e-08 0 2.5605e-08 0.0007 2.5608e-08 0 2.5802e-08 0 2.5805e-08 0.0007 2.5808e-08 0 2.6002e-08 0 2.6005e-08 0.0007 2.6008e-08 0 2.6202e-08 0 2.6205e-08 0.0007 2.6208e-08 0 2.6402e-08 0 2.6405e-08 0.0007 2.6408e-08 0 2.6602e-08 0 2.6605e-08 0.0007 2.6608e-08 0 2.6802e-08 0 2.6805e-08 0.0007 2.6808e-08 0 2.7002e-08 0 2.7005e-08 0.0007 2.7008e-08 0 2.7202e-08 0 2.7205e-08 0.0007 2.7208e-08 0 2.7402e-08 0 2.7405e-08 0.0007 2.7408e-08 0 2.7602e-08 0 2.7605e-08 0.0007 2.7608e-08 0 2.7802e-08 0 2.7805e-08 0.0007 2.7808e-08 0 2.8002e-08 0 2.8005e-08 0.0007 2.8008e-08 0 2.8202e-08 0 2.8205e-08 0.0007 2.8208e-08 0 2.8402e-08 0 2.8405e-08 0.0007 2.8408e-08 0 2.8602e-08 0 2.8605e-08 0.0007 2.8608e-08 0 2.8802e-08 0 2.8805e-08 0.0007 2.8808e-08 0 2.9002e-08 0 2.9005e-08 0.0007 2.9008e-08 0 2.9202e-08 0 2.9205e-08 0.0007 2.9208e-08 0 2.9402e-08 0 2.9405e-08 0.0007 2.9408e-08 0 2.9602e-08 0 2.9605e-08 0.0007 2.9608e-08 0 2.9802e-08 0 2.9805e-08 0.0007 2.9808e-08 0 3.0002e-08 0 3.0005e-08 0.0007 3.0008e-08 0 3.0202e-08 0 3.0205e-08 0.0007 3.0208e-08 0 3.0402e-08 0 3.0405e-08 0.0007 3.0408e-08 0 3.0602e-08 0 3.0605e-08 0.0007 3.0608e-08 0 3.0802e-08 0 3.0805e-08 0.0007 3.0808e-08 0 3.1002e-08 0 3.1005e-08 0.0007 3.1008e-08 0 3.1202e-08 0 3.1205e-08 0.0007 3.1208e-08 0 3.1402e-08 0 3.1405e-08 0.0007 3.1408e-08 0 3.1602e-08 0 3.1605e-08 0.0007 3.1608e-08 0 3.1802e-08 0 3.1805e-08 0.0007 3.1808e-08 0 3.2002e-08 0 3.2005e-08 0.0007 3.2008e-08 0 3.2202e-08 0 3.2205e-08 0.0007 3.2208e-08 0 3.2402e-08 0 3.2405e-08 0.0007 3.2408e-08 0 3.2602e-08 0 3.2605e-08 0.0007 3.2608e-08 0 3.2802e-08 0 3.2805e-08 0.0007 3.2808e-08 0 3.3002e-08 0 3.3005e-08 0.0007 3.3008e-08 0 3.3202e-08 0 3.3205e-08 0.0007 3.3208e-08 0 3.3402e-08 0 3.3405e-08 0.0007 3.3408e-08 0 3.3602e-08 0 3.3605e-08 0.0007 3.3608e-08 0 3.3802e-08 0 3.3805e-08 0.0007 3.3808e-08 0 3.4002e-08 0 3.4005e-08 0.0007 3.4008e-08 0 3.4202e-08 0 3.4205e-08 0.0007 3.4208e-08 0 3.4402e-08 0 3.4405e-08 0.0007 3.4408e-08 0 3.4602e-08 0 3.4605e-08 0.0007 3.4608e-08 0 3.4802e-08 0 3.4805e-08 0.0007 3.4808e-08 0 3.5002e-08 0 3.5005e-08 0.0007 3.5008e-08 0 3.5202e-08 0 3.5205e-08 0.0007 3.5208e-08 0 3.5402e-08 0 3.5405e-08 0.0007 3.5408e-08 0 3.5602e-08 0 3.5605e-08 0.0007 3.5608e-08 0 3.5802e-08 0 3.5805e-08 0.0007 3.5808e-08 0 3.6002e-08 0 3.6005e-08 0.0007 3.6008e-08 0 3.6202e-08 0 3.6205e-08 0.0007 3.6208e-08 0 3.6402e-08 0 3.6405e-08 0.0007 3.6408e-08 0 3.6602e-08 0 3.6605e-08 0.0007 3.6608e-08 0 3.6802e-08 0 3.6805e-08 0.0007 3.6808e-08 0 3.7002e-08 0 3.7005e-08 0.0007 3.7008e-08 0 3.7202e-08 0 3.7205e-08 0.0007 3.7208e-08 0 3.7402e-08 0 3.7405e-08 0.0007 3.7408e-08 0 3.7602e-08 0 3.7605e-08 0.0007 3.7608e-08 0 3.7802e-08 0 3.7805e-08 0.0007 3.7808e-08 0 3.8002e-08 0 3.8005e-08 0.0007 3.8008e-08 0 3.8202e-08 0 3.8205e-08 0.0007 3.8208e-08 0 3.8402e-08 0 3.8405e-08 0.0007 3.8408e-08 0 3.8602e-08 0 3.8605e-08 0.0007 3.8608e-08 0 3.8802e-08 0 3.8805e-08 0.0007 3.8808e-08 0 3.9002e-08 0 3.9005e-08 0.0007 3.9008e-08 0 3.9202e-08 0 3.9205e-08 0.0007 3.9208e-08 0 3.9402e-08 0 3.9405e-08 0.0007 3.9408e-08 0 3.9602e-08 0 3.9605e-08 0.0007 3.9608e-08 0 3.9802e-08 0 3.9805e-08 0.0007 3.9808e-08 0 4.0002e-08 0 4.0005e-08 0.0007 4.0008e-08 0 4.0202e-08 0 4.0205e-08 0.0007 4.0208e-08 0 4.0402e-08 0 4.0405e-08 0.0007 4.0408e-08 0 4.0602e-08 0 4.0605e-08 0.0007 4.0608e-08 0 4.0802e-08 0 4.0805e-08 0.0007 4.0808e-08 0 4.1002e-08 0 4.1005e-08 0.0007 4.1008e-08 0 4.1202e-08 0 4.1205e-08 0.0007 4.1208e-08 0 4.1402e-08 0 4.1405e-08 0.0007 4.1408e-08 0 4.1602e-08 0 4.1605e-08 0.0007 4.1608e-08 0 4.1802e-08 0 4.1805e-08 0.0007 4.1808e-08 0 4.2002e-08 0 4.2005e-08 0.0007 4.2008e-08 0 4.2202e-08 0 4.2205e-08 0.0007 4.2208e-08 0 4.2402e-08 0 4.2405e-08 0.0007 4.2408e-08 0 4.2602e-08 0 4.2605e-08 0.0007 4.2608e-08 0 4.2802e-08 0 4.2805e-08 0.0007 4.2808e-08 0 4.3002e-08 0 4.3005e-08 0.0007 4.3008e-08 0 4.3202e-08 0 4.3205e-08 0.0007 4.3208e-08 0 4.3402e-08 0 4.3405e-08 0.0007 4.3408e-08 0 4.3602e-08 0 4.3605e-08 0.0007 4.3608e-08 0 4.3802e-08 0 4.3805e-08 0.0007 4.3808e-08 0 4.4002e-08 0 4.4005e-08 0.0007 4.4008e-08 0 4.4202e-08 0 4.4205e-08 0.0007 4.4208e-08 0 4.4402e-08 0 4.4405e-08 0.0007 4.4408e-08 0 4.4602e-08 0 4.4605e-08 0.0007 4.4608e-08 0 4.4802e-08 0 4.4805e-08 0.0007 4.4808e-08 0 4.5002e-08 0 4.5005e-08 0.0007 4.5008e-08 0 4.5202e-08 0 4.5205e-08 0.0007 4.5208e-08 0 4.5402e-08 0 4.5405e-08 0.0007 4.5408e-08 0 4.5602e-08 0 4.5605e-08 0.0007 4.5608e-08 0 4.5802e-08 0 4.5805e-08 0.0007 4.5808e-08 0 4.6002e-08 0 4.6005e-08 0.0007 4.6008e-08 0 4.6202e-08 0 4.6205e-08 0.0007 4.6208e-08 0 4.6402e-08 0 4.6405e-08 0.0007 4.6408e-08 0 4.6602e-08 0 4.6605e-08 0.0007 4.6608e-08 0 4.6802e-08 0 4.6805e-08 0.0007 4.6808e-08 0 4.7002e-08 0 4.7005e-08 0.0007 4.7008e-08 0 4.7202e-08 0 4.7205e-08 0.0007 4.7208e-08 0 4.7402e-08 0 4.7405e-08 0.0007 4.7408e-08 0 4.7602e-08 0 4.7605e-08 0.0007 4.7608e-08 0 4.7802e-08 0 4.7805e-08 0.0007 4.7808e-08 0 4.8002e-08 0 4.8005e-08 0.0007 4.8008e-08 0 4.8202e-08 0 4.8205e-08 0.0007 4.8208e-08 0 4.8402e-08 0 4.8405e-08 0.0007 4.8408e-08 0 4.8602e-08 0 4.8605e-08 0.0007 4.8608e-08 0 4.8802e-08 0 4.8805e-08 0.0007 4.8808e-08 0 4.9002e-08 0 4.9005e-08 0.0007 4.9008e-08 0 4.9202e-08 0 4.9205e-08 0.0007 4.9208e-08 0 4.9402e-08 0 4.9405e-08 0.0007 4.9408e-08 0 4.9602e-08 0 4.9605e-08 0.0007 4.9608e-08 0 4.9802e-08 0 4.9805e-08 0.0007 4.9808e-08 0 5.0002e-08 0 5.0005e-08 0.0007 5.0008e-08 0 5.0202e-08 0 5.0205e-08 0.0007 5.0208e-08 0 5.0402e-08 0 5.0405e-08 0.0007 5.0408e-08 0 5.0602e-08 0 5.0605e-08 0.0007 5.0608e-08 0 5.0802e-08 0 5.0805e-08 0.0007 5.0808e-08 0 5.1002e-08 0 5.1005e-08 0.0007 5.1008e-08 0 5.1202e-08 0 5.1205e-08 0.0007 5.1208e-08 0 5.1402e-08 0 5.1405e-08 0.0007 5.1408e-08 0 5.1602e-08 0 5.1605e-08 0.0007 5.1608e-08 0 5.1802e-08 0 5.1805e-08 0.0007 5.1808e-08 0 5.2002e-08 0 5.2005e-08 0.0007 5.2008e-08 0 5.2202e-08 0 5.2205e-08 0.0007 5.2208e-08 0 5.2402e-08 0 5.2405e-08 0.0007 5.2408e-08 0 5.2602e-08 0 5.2605e-08 0.0007 5.2608e-08 0 5.2802e-08 0 5.2805e-08 0.0007 5.2808e-08 0 5.3002e-08 0 5.3005e-08 0.0007 5.3008e-08 0 5.3202e-08 0 5.3205e-08 0.0007 5.3208e-08 0 5.3402e-08 0 5.3405e-08 0.0007 5.3408e-08 0 5.3602e-08 0 5.3605e-08 0.0007 5.3608e-08 0 5.3802e-08 0 5.3805e-08 0.0007 5.3808e-08 0 5.4002e-08 0 5.4005e-08 0.0007 5.4008e-08 0 5.4202e-08 0 5.4205e-08 0.0007 5.4208e-08 0 5.4402e-08 0 5.4405e-08 0.0007 5.4408e-08 0 5.4602e-08 0 5.4605e-08 0.0007 5.4608e-08 0 5.4802e-08 0 5.4805e-08 0.0007 5.4808e-08 0 5.5002e-08 0 5.5005e-08 0.0007 5.5008e-08 0 5.5202e-08 0 5.5205e-08 0.0007 5.5208e-08 0 5.5402e-08 0 5.5405e-08 0.0007 5.5408e-08 0 5.5602e-08 0 5.5605e-08 0.0007 5.5608e-08 0 5.5802e-08 0 5.5805e-08 0.0007 5.5808e-08 0 5.6002e-08 0 5.6005e-08 0.0007 5.6008e-08 0 5.6202e-08 0 5.6205e-08 0.0007 5.6208e-08 0 5.6402e-08 0 5.6405e-08 0.0007 5.6408e-08 0 5.6602e-08 0 5.6605e-08 0.0007 5.6608e-08 0 5.6802e-08 0 5.6805e-08 0.0007 5.6808e-08 0 5.7002e-08 0 5.7005e-08 0.0007 5.7008e-08 0 5.7202e-08 0 5.7205e-08 0.0007 5.7208e-08 0 5.7402e-08 0 5.7405e-08 0.0007 5.7408e-08 0 5.7602e-08 0 5.7605e-08 0.0007 5.7608e-08 0 5.7802e-08 0 5.7805e-08 0.0007 5.7808e-08 0 5.8002e-08 0 5.8005e-08 0.0007 5.8008e-08 0 5.8202e-08 0 5.8205e-08 0.0007 5.8208e-08 0 5.8402e-08 0 5.8405e-08 0.0007 5.8408e-08 0 5.8602e-08 0 5.8605e-08 0.0007 5.8608e-08 0 5.8802e-08 0 5.8805e-08 0.0007 5.8808e-08 0 5.9002e-08 0 5.9005e-08 0.0007 5.9008e-08 0 5.9202e-08 0 5.9205e-08 0.0007 5.9208e-08 0 5.9402e-08 0 5.9405e-08 0.0007 5.9408e-08 0 5.9602e-08 0 5.9605e-08 0.0007 5.9608e-08 0 5.9802e-08 0 5.9805e-08 0.0007 5.9808e-08 0 6.0002e-08 0 6.0005e-08 0.0007 6.0008e-08 0 6.0202e-08 0 6.0205e-08 0.0007 6.0208e-08 0 6.0402e-08 0 6.0405e-08 0.0007 6.0408e-08 0 6.0602e-08 0 6.0605e-08 0.0007 6.0608e-08 0 6.0802e-08 0 6.0805e-08 0.0007 6.0808e-08 0 6.1002e-08 0 6.1005e-08 0.0007 6.1008e-08 0 6.1202e-08 0 6.1205e-08 0.0007 6.1208e-08 0 6.1402e-08 0 6.1405e-08 0.0007 6.1408e-08 0 6.1602e-08 0 6.1605e-08 0.0007 6.1608e-08 0 6.1802e-08 0 6.1805e-08 0.0007 6.1808e-08 0 6.2002e-08 0 6.2005e-08 0.0007 6.2008e-08 0 6.2202e-08 0 6.2205e-08 0.0007 6.2208e-08 0 6.2402e-08 0 6.2405e-08 0.0007 6.2408e-08 0 6.2602e-08 0 6.2605e-08 0.0007 6.2608e-08 0 6.2802e-08 0 6.2805e-08 0.0007 6.2808e-08 0 6.3002e-08 0 6.3005e-08 0.0007 6.3008e-08 0 6.3202e-08 0 6.3205e-08 0.0007 6.3208e-08 0 6.3402e-08 0 6.3405e-08 0.0007 6.3408e-08 0 6.3602e-08 0 6.3605e-08 0.0007 6.3608e-08 0 6.3802e-08 0 6.3805e-08 0.0007 6.3808e-08 0 6.4002e-08 0 6.4005e-08 0.0007 6.4008e-08 0 6.4202e-08 0 6.4205e-08 0.0007 6.4208e-08 0 6.4402e-08 0 6.4405e-08 0.0007 6.4408e-08 0 6.4602e-08 0 6.4605e-08 0.0007 6.4608e-08 0 6.4802e-08 0 6.4805e-08 0.0007 6.4808e-08 0 6.5002e-08 0 6.5005e-08 0.0007 6.5008e-08 0 6.5202e-08 0 6.5205e-08 0.0007 6.5208e-08 0 6.5402e-08 0 6.5405e-08 0.0007 6.5408e-08 0 6.5602e-08 0 6.5605e-08 0.0007 6.5608e-08 0 6.5802e-08 0 6.5805e-08 0.0007 6.5808e-08 0 6.6002e-08 0 6.6005e-08 0.0007 6.6008e-08 0 6.6202e-08 0 6.6205e-08 0.0007 6.6208e-08 0 6.6402e-08 0 6.6405e-08 0.0007 6.6408e-08 0 6.6602e-08 0 6.6605e-08 0.0007 6.6608e-08 0 6.6802e-08 0 6.6805e-08 0.0007 6.6808e-08 0 6.7002e-08 0 6.7005e-08 0.0007 6.7008e-08 0 6.7202e-08 0 6.7205e-08 0.0007 6.7208e-08 0 6.7402e-08 0 6.7405e-08 0.0007 6.7408e-08 0 6.7602e-08 0 6.7605e-08 0.0007 6.7608e-08 0 6.7802e-08 0 6.7805e-08 0.0007 6.7808e-08 0 6.8002e-08 0 6.8005e-08 0.0007 6.8008e-08 0 6.8202e-08 0 6.8205e-08 0.0007 6.8208e-08 0 6.8402e-08 0 6.8405e-08 0.0007 6.8408e-08 0 6.8602e-08 0 6.8605e-08 0.0007 6.8608e-08 0 6.8802e-08 0 6.8805e-08 0.0007 6.8808e-08 0 6.9002e-08 0 6.9005e-08 0.0007 6.9008e-08 0 6.9202e-08 0 6.9205e-08 0.0007 6.9208e-08 0 6.9402e-08 0 6.9405e-08 0.0007 6.9408e-08 0 6.9602e-08 0 6.9605e-08 0.0007 6.9608e-08 0 6.9802e-08 0 6.9805e-08 0.0007 6.9808e-08 0 7.0002e-08 0 7.0005e-08 0.0007 7.0008e-08 0 7.0202e-08 0 7.0205e-08 0.0007 7.0208e-08 0 7.0402e-08 0 7.0405e-08 0.0007 7.0408e-08 0 7.0602e-08 0 7.0605e-08 0.0007 7.0608e-08 0 7.0802e-08 0 7.0805e-08 0.0007 7.0808e-08 0 7.1002e-08 0 7.1005e-08 0.0007 7.1008e-08 0 7.1202e-08 0 7.1205e-08 0.0007 7.1208e-08 0 7.1402e-08 0 7.1405e-08 0.0007 7.1408e-08 0 7.1602e-08 0 7.1605e-08 0.0007 7.1608e-08 0 7.1802e-08 0 7.1805e-08 0.0007 7.1808e-08 0 7.2002e-08 0 7.2005e-08 0.0007 7.2008e-08 0 7.2202e-08 0 7.2205e-08 0.0007 7.2208e-08 0 7.2402e-08 0 7.2405e-08 0.0007 7.2408e-08 0 7.2602e-08 0 7.2605e-08 0.0007 7.2608e-08 0 7.2802e-08 0 7.2805e-08 0.0007 7.2808e-08 0 7.3002e-08 0 7.3005e-08 0.0007 7.3008e-08 0 7.3202e-08 0 7.3205e-08 0.0007 7.3208e-08 0 7.3402e-08 0 7.3405e-08 0.0007 7.3408e-08 0 7.3602e-08 0 7.3605e-08 0.0007 7.3608e-08 0 7.3802e-08 0 7.3805e-08 0.0007 7.3808e-08 0 7.4002e-08 0 7.4005e-08 0.0007 7.4008e-08 0 7.4202e-08 0 7.4205e-08 0.0007 7.4208e-08 0 7.4402e-08 0 7.4405e-08 0.0007 7.4408e-08 0 7.4602e-08 0 7.4605e-08 0.0007 7.4608e-08 0 7.4802e-08 0 7.4805e-08 0.0007 7.4808e-08 0 7.5002e-08 0 7.5005e-08 0.0007 7.5008e-08 0 7.5202e-08 0 7.5205e-08 0.0007 7.5208e-08 0 7.5402e-08 0 7.5405e-08 0.0007 7.5408e-08 0 7.5602e-08 0 7.5605e-08 0.0007 7.5608e-08 0 7.5802e-08 0 7.5805e-08 0.0007 7.5808e-08 0 7.6002e-08 0 7.6005e-08 0.0007 7.6008e-08 0 7.6202e-08 0 7.6205e-08 0.0007 7.6208e-08 0 7.6402e-08 0 7.6405e-08 0.0007 7.6408e-08 0 7.6602e-08 0 7.6605e-08 0.0007 7.6608e-08 0 7.6802e-08 0 7.6805e-08 0.0007 7.6808e-08 0 7.7002e-08 0 7.7005e-08 0.0007 7.7008e-08 0 7.7202e-08 0 7.7205e-08 0.0007 7.7208e-08 0 7.7402e-08 0 7.7405e-08 0.0007 7.7408e-08 0 7.7602e-08 0 7.7605e-08 0.0007 7.7608e-08 0 7.7802e-08 0 7.7805e-08 0.0007 7.7808e-08 0 7.8002e-08 0 7.8005e-08 0.0007 7.8008e-08 0 7.8202e-08 0 7.8205e-08 0.0007 7.8208e-08 0 7.8402e-08 0 7.8405e-08 0.0007 7.8408e-08 0 7.8602e-08 0 7.8605e-08 0.0007 7.8608e-08 0 7.8802e-08 0 7.8805e-08 0.0007 7.8808e-08 0 7.9002e-08 0 7.9005e-08 0.0007 7.9008e-08 0 7.9202e-08 0 7.9205e-08 0.0007 7.9208e-08 0 7.9402e-08 0 7.9405e-08 0.0007 7.9408e-08 0 7.9602e-08 0 7.9605e-08 0.0007 7.9608e-08 0)
L_S4|1 G3_2 _S4|A1  2.067833848e-12
L_S4|2 _S4|A1 _S4|A2  4.135667696e-12
L_S4|3 _S4|A3 _S4|A4  8.271335392e-12
L_S4|T T16 _S4|T1  2.067833848e-12
L_S4|4 _S4|T1 _S4|T2  4.135667696e-12
L_S4|5 _S4|A4 _S4|Q1  4.135667696e-12
L_S4|6 _S4|Q1 S4  2.067833848e-12
LI0|_SPL_A|1 A0 I0|_SPL_A|D1  2e-12
LI0|_SPL_A|2 I0|_SPL_A|D1 I0|_SPL_A|D2  4.135667696e-12
LI0|_SPL_A|3 I0|_SPL_A|D2 I0|_SPL_A|JCT  9.84682784761905e-13
LI0|_SPL_A|4 I0|_SPL_A|JCT I0|_SPL_A|QA1  9.84682784761905e-13
LI0|_SPL_A|5 I0|_SPL_A|QA1 I0|A1  2e-12
LI0|_SPL_A|6 I0|_SPL_A|JCT I0|_SPL_A|QB1  9.84682784761905e-13
LI0|_SPL_A|7 I0|_SPL_A|QB1 I0|A2  2e-12
LI0|_SPL_B|1 B0 I0|_SPL_B|D1  2e-12
LI0|_SPL_B|2 I0|_SPL_B|D1 I0|_SPL_B|D2  4.135667696e-12
LI0|_SPL_B|3 I0|_SPL_B|D2 I0|_SPL_B|JCT  9.84682784761905e-13
LI0|_SPL_B|4 I0|_SPL_B|JCT I0|_SPL_B|QA1  9.84682784761905e-13
LI0|_SPL_B|5 I0|_SPL_B|QA1 I0|B1  2e-12
LI0|_SPL_B|6 I0|_SPL_B|JCT I0|_SPL_B|QB1  9.84682784761905e-13
LI0|_SPL_B|7 I0|_SPL_B|QB1 I0|B2  2e-12
LI0|_DFF_A|1 I0|A1 I0|_DFF_A|A1  2.067833848e-12
LI0|_DFF_A|2 I0|_DFF_A|A1 I0|_DFF_A|A2  4.135667696e-12
LI0|_DFF_A|3 I0|_DFF_A|A3 I0|_DFF_A|A4  8.271335392e-12
LI0|_DFF_A|T T00 I0|_DFF_A|T1  2.067833848e-12
LI0|_DFF_A|4 I0|_DFF_A|T1 I0|_DFF_A|T2  4.135667696e-12
LI0|_DFF_A|5 I0|_DFF_A|A4 I0|_DFF_A|Q1  4.135667696e-12
LI0|_DFF_A|6 I0|_DFF_A|Q1 I0|A1_SYNC  2.067833848e-12
LI0|_DFF_B|1 I0|B1 I0|_DFF_B|A1  2.067833848e-12
LI0|_DFF_B|2 I0|_DFF_B|A1 I0|_DFF_B|A2  4.135667696e-12
LI0|_DFF_B|3 I0|_DFF_B|A3 I0|_DFF_B|A4  8.271335392e-12
LI0|_DFF_B|T T00 I0|_DFF_B|T1  2.067833848e-12
LI0|_DFF_B|4 I0|_DFF_B|T1 I0|_DFF_B|T2  4.135667696e-12
LI0|_DFF_B|5 I0|_DFF_B|A4 I0|_DFF_B|Q1  4.135667696e-12
LI0|_DFF_B|6 I0|_DFF_B|Q1 I0|B1_SYNC  2.067833848e-12
LI0|_XOR|A1 I0|A2 I0|_XOR|A1  2.067833848e-12
LI0|_XOR|A2 I0|_XOR|A1 I0|_XOR|A2  4.135667696e-12
LI0|_XOR|A3 I0|_XOR|A3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|B1 I0|B2 I0|_XOR|B1  2.067833848e-12
LI0|_XOR|B2 I0|_XOR|B1 I0|_XOR|B2  4.135667696e-12
LI0|_XOR|B3 I0|_XOR|B3 I0|_XOR|AB  8.271335392e-12
LI0|_XOR|T1 T00 I0|_XOR|T1  2.067833848e-12
LI0|_XOR|T2 I0|_XOR|T1 I0|_XOR|T2  4.135667696e-12
LI0|_XOR|Q2 I0|_XOR|ABTQ I0|_XOR|Q1  4.135667696e-12
LI0|_XOR|Q1 I0|_XOR|Q1 IP0_0  2.067833848e-12
LI0|_AND|A1 I0|A1_SYNC I0|_AND|A1  2.067833848e-12
LI0|_AND|A2 I0|_AND|A1 I0|_AND|A2  4.135667696e-12
LI0|_AND|A3 I0|_AND|A3 I0|_AND|Q3  1.2e-12
LI0|_AND|B1 I0|B1_SYNC I0|_AND|B1  2.067833848e-12
LI0|_AND|B2 I0|_AND|B1 I0|_AND|B2  4.135667696e-12
LI0|_AND|B3 I0|_AND|B3 I0|_AND|Q3  1.2e-12
LI0|_AND|Q3 I0|_AND|Q3 I0|_AND|Q2  4.135667696e-12
LI0|_AND|Q2 I0|_AND|Q2 I0|_AND|Q1  4.135667696e-12
LI0|_AND|Q1 I0|_AND|Q1 IG0_0  2.067833848e-12
LI1|_SPL_A|1 A1 I1|_SPL_A|D1  2e-12
LI1|_SPL_A|2 I1|_SPL_A|D1 I1|_SPL_A|D2  4.135667696e-12
LI1|_SPL_A|3 I1|_SPL_A|D2 I1|_SPL_A|JCT  9.84682784761905e-13
LI1|_SPL_A|4 I1|_SPL_A|JCT I1|_SPL_A|QA1  9.84682784761905e-13
LI1|_SPL_A|5 I1|_SPL_A|QA1 I1|A1  2e-12
LI1|_SPL_A|6 I1|_SPL_A|JCT I1|_SPL_A|QB1  9.84682784761905e-13
LI1|_SPL_A|7 I1|_SPL_A|QB1 I1|A2  2e-12
LI1|_SPL_B|1 B1 I1|_SPL_B|D1  2e-12
LI1|_SPL_B|2 I1|_SPL_B|D1 I1|_SPL_B|D2  4.135667696e-12
LI1|_SPL_B|3 I1|_SPL_B|D2 I1|_SPL_B|JCT  9.84682784761905e-13
LI1|_SPL_B|4 I1|_SPL_B|JCT I1|_SPL_B|QA1  9.84682784761905e-13
LI1|_SPL_B|5 I1|_SPL_B|QA1 I1|B1  2e-12
LI1|_SPL_B|6 I1|_SPL_B|JCT I1|_SPL_B|QB1  9.84682784761905e-13
LI1|_SPL_B|7 I1|_SPL_B|QB1 I1|B2  2e-12
LI1|_DFF_A|1 I1|A1 I1|_DFF_A|A1  2.067833848e-12
LI1|_DFF_A|2 I1|_DFF_A|A1 I1|_DFF_A|A2  4.135667696e-12
LI1|_DFF_A|3 I1|_DFF_A|A3 I1|_DFF_A|A4  8.271335392e-12
LI1|_DFF_A|T T01 I1|_DFF_A|T1  2.067833848e-12
LI1|_DFF_A|4 I1|_DFF_A|T1 I1|_DFF_A|T2  4.135667696e-12
LI1|_DFF_A|5 I1|_DFF_A|A4 I1|_DFF_A|Q1  4.135667696e-12
LI1|_DFF_A|6 I1|_DFF_A|Q1 I1|A1_SYNC  2.067833848e-12
LI1|_DFF_B|1 I1|B1 I1|_DFF_B|A1  2.067833848e-12
LI1|_DFF_B|2 I1|_DFF_B|A1 I1|_DFF_B|A2  4.135667696e-12
LI1|_DFF_B|3 I1|_DFF_B|A3 I1|_DFF_B|A4  8.271335392e-12
LI1|_DFF_B|T T01 I1|_DFF_B|T1  2.067833848e-12
LI1|_DFF_B|4 I1|_DFF_B|T1 I1|_DFF_B|T2  4.135667696e-12
LI1|_DFF_B|5 I1|_DFF_B|A4 I1|_DFF_B|Q1  4.135667696e-12
LI1|_DFF_B|6 I1|_DFF_B|Q1 I1|B1_SYNC  2.067833848e-12
LI1|_XOR|A1 I1|A2 I1|_XOR|A1  2.067833848e-12
LI1|_XOR|A2 I1|_XOR|A1 I1|_XOR|A2  4.135667696e-12
LI1|_XOR|A3 I1|_XOR|A3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|B1 I1|B2 I1|_XOR|B1  2.067833848e-12
LI1|_XOR|B2 I1|_XOR|B1 I1|_XOR|B2  4.135667696e-12
LI1|_XOR|B3 I1|_XOR|B3 I1|_XOR|AB  8.271335392e-12
LI1|_XOR|T1 T01 I1|_XOR|T1  2.067833848e-12
LI1|_XOR|T2 I1|_XOR|T1 I1|_XOR|T2  4.135667696e-12
LI1|_XOR|Q2 I1|_XOR|ABTQ I1|_XOR|Q1  4.135667696e-12
LI1|_XOR|Q1 I1|_XOR|Q1 IP1_0  2.067833848e-12
LI1|_AND|A1 I1|A1_SYNC I1|_AND|A1  2.067833848e-12
LI1|_AND|A2 I1|_AND|A1 I1|_AND|A2  4.135667696e-12
LI1|_AND|A3 I1|_AND|A3 I1|_AND|Q3  1.2e-12
LI1|_AND|B1 I1|B1_SYNC I1|_AND|B1  2.067833848e-12
LI1|_AND|B2 I1|_AND|B1 I1|_AND|B2  4.135667696e-12
LI1|_AND|B3 I1|_AND|B3 I1|_AND|Q3  1.2e-12
LI1|_AND|Q3 I1|_AND|Q3 I1|_AND|Q2  4.135667696e-12
LI1|_AND|Q2 I1|_AND|Q2 I1|_AND|Q1  4.135667696e-12
LI1|_AND|Q1 I1|_AND|Q1 IG1_0  2.067833848e-12
LI2|_SPL_A|1 A2 I2|_SPL_A|D1  2e-12
LI2|_SPL_A|2 I2|_SPL_A|D1 I2|_SPL_A|D2  4.135667696e-12
LI2|_SPL_A|3 I2|_SPL_A|D2 I2|_SPL_A|JCT  9.84682784761905e-13
LI2|_SPL_A|4 I2|_SPL_A|JCT I2|_SPL_A|QA1  9.84682784761905e-13
LI2|_SPL_A|5 I2|_SPL_A|QA1 I2|A1  2e-12
LI2|_SPL_A|6 I2|_SPL_A|JCT I2|_SPL_A|QB1  9.84682784761905e-13
LI2|_SPL_A|7 I2|_SPL_A|QB1 I2|A2  2e-12
LI2|_SPL_B|1 B2 I2|_SPL_B|D1  2e-12
LI2|_SPL_B|2 I2|_SPL_B|D1 I2|_SPL_B|D2  4.135667696e-12
LI2|_SPL_B|3 I2|_SPL_B|D2 I2|_SPL_B|JCT  9.84682784761905e-13
LI2|_SPL_B|4 I2|_SPL_B|JCT I2|_SPL_B|QA1  9.84682784761905e-13
LI2|_SPL_B|5 I2|_SPL_B|QA1 I2|B1  2e-12
LI2|_SPL_B|6 I2|_SPL_B|JCT I2|_SPL_B|QB1  9.84682784761905e-13
LI2|_SPL_B|7 I2|_SPL_B|QB1 I2|B2  2e-12
LI2|_DFF_A|1 I2|A1 I2|_DFF_A|A1  2.067833848e-12
LI2|_DFF_A|2 I2|_DFF_A|A1 I2|_DFF_A|A2  4.135667696e-12
LI2|_DFF_A|3 I2|_DFF_A|A3 I2|_DFF_A|A4  8.271335392e-12
LI2|_DFF_A|T T02 I2|_DFF_A|T1  2.067833848e-12
LI2|_DFF_A|4 I2|_DFF_A|T1 I2|_DFF_A|T2  4.135667696e-12
LI2|_DFF_A|5 I2|_DFF_A|A4 I2|_DFF_A|Q1  4.135667696e-12
LI2|_DFF_A|6 I2|_DFF_A|Q1 I2|A1_SYNC  2.067833848e-12
LI2|_DFF_B|1 I2|B1 I2|_DFF_B|A1  2.067833848e-12
LI2|_DFF_B|2 I2|_DFF_B|A1 I2|_DFF_B|A2  4.135667696e-12
LI2|_DFF_B|3 I2|_DFF_B|A3 I2|_DFF_B|A4  8.271335392e-12
LI2|_DFF_B|T T02 I2|_DFF_B|T1  2.067833848e-12
LI2|_DFF_B|4 I2|_DFF_B|T1 I2|_DFF_B|T2  4.135667696e-12
LI2|_DFF_B|5 I2|_DFF_B|A4 I2|_DFF_B|Q1  4.135667696e-12
LI2|_DFF_B|6 I2|_DFF_B|Q1 I2|B1_SYNC  2.067833848e-12
LI2|_XOR|A1 I2|A2 I2|_XOR|A1  2.067833848e-12
LI2|_XOR|A2 I2|_XOR|A1 I2|_XOR|A2  4.135667696e-12
LI2|_XOR|A3 I2|_XOR|A3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|B1 I2|B2 I2|_XOR|B1  2.067833848e-12
LI2|_XOR|B2 I2|_XOR|B1 I2|_XOR|B2  4.135667696e-12
LI2|_XOR|B3 I2|_XOR|B3 I2|_XOR|AB  8.271335392e-12
LI2|_XOR|T1 T02 I2|_XOR|T1  2.067833848e-12
LI2|_XOR|T2 I2|_XOR|T1 I2|_XOR|T2  4.135667696e-12
LI2|_XOR|Q2 I2|_XOR|ABTQ I2|_XOR|Q1  4.135667696e-12
LI2|_XOR|Q1 I2|_XOR|Q1 IP2_0  2.067833848e-12
LI2|_AND|A1 I2|A1_SYNC I2|_AND|A1  2.067833848e-12
LI2|_AND|A2 I2|_AND|A1 I2|_AND|A2  4.135667696e-12
LI2|_AND|A3 I2|_AND|A3 I2|_AND|Q3  1.2e-12
LI2|_AND|B1 I2|B1_SYNC I2|_AND|B1  2.067833848e-12
LI2|_AND|B2 I2|_AND|B1 I2|_AND|B2  4.135667696e-12
LI2|_AND|B3 I2|_AND|B3 I2|_AND|Q3  1.2e-12
LI2|_AND|Q3 I2|_AND|Q3 I2|_AND|Q2  4.135667696e-12
LI2|_AND|Q2 I2|_AND|Q2 I2|_AND|Q1  4.135667696e-12
LI2|_AND|Q1 I2|_AND|Q1 IG2_0  2.067833848e-12
LI3|_SPL_A|1 A3 I3|_SPL_A|D1  2e-12
LI3|_SPL_A|2 I3|_SPL_A|D1 I3|_SPL_A|D2  4.135667696e-12
LI3|_SPL_A|3 I3|_SPL_A|D2 I3|_SPL_A|JCT  9.84682784761905e-13
LI3|_SPL_A|4 I3|_SPL_A|JCT I3|_SPL_A|QA1  9.84682784761905e-13
LI3|_SPL_A|5 I3|_SPL_A|QA1 I3|A1  2e-12
LI3|_SPL_A|6 I3|_SPL_A|JCT I3|_SPL_A|QB1  9.84682784761905e-13
LI3|_SPL_A|7 I3|_SPL_A|QB1 I3|A2  2e-12
LI3|_SPL_B|1 B3 I3|_SPL_B|D1  2e-12
LI3|_SPL_B|2 I3|_SPL_B|D1 I3|_SPL_B|D2  4.135667696e-12
LI3|_SPL_B|3 I3|_SPL_B|D2 I3|_SPL_B|JCT  9.84682784761905e-13
LI3|_SPL_B|4 I3|_SPL_B|JCT I3|_SPL_B|QA1  9.84682784761905e-13
LI3|_SPL_B|5 I3|_SPL_B|QA1 I3|B1  2e-12
LI3|_SPL_B|6 I3|_SPL_B|JCT I3|_SPL_B|QB1  9.84682784761905e-13
LI3|_SPL_B|7 I3|_SPL_B|QB1 I3|B2  2e-12
LI3|_DFF_A|1 I3|A1 I3|_DFF_A|A1  2.067833848e-12
LI3|_DFF_A|2 I3|_DFF_A|A1 I3|_DFF_A|A2  4.135667696e-12
LI3|_DFF_A|3 I3|_DFF_A|A3 I3|_DFF_A|A4  8.271335392e-12
LI3|_DFF_A|T T03 I3|_DFF_A|T1  2.067833848e-12
LI3|_DFF_A|4 I3|_DFF_A|T1 I3|_DFF_A|T2  4.135667696e-12
LI3|_DFF_A|5 I3|_DFF_A|A4 I3|_DFF_A|Q1  4.135667696e-12
LI3|_DFF_A|6 I3|_DFF_A|Q1 I3|A1_SYNC  2.067833848e-12
LI3|_DFF_B|1 I3|B1 I3|_DFF_B|A1  2.067833848e-12
LI3|_DFF_B|2 I3|_DFF_B|A1 I3|_DFF_B|A2  4.135667696e-12
LI3|_DFF_B|3 I3|_DFF_B|A3 I3|_DFF_B|A4  8.271335392e-12
LI3|_DFF_B|T T03 I3|_DFF_B|T1  2.067833848e-12
LI3|_DFF_B|4 I3|_DFF_B|T1 I3|_DFF_B|T2  4.135667696e-12
LI3|_DFF_B|5 I3|_DFF_B|A4 I3|_DFF_B|Q1  4.135667696e-12
LI3|_DFF_B|6 I3|_DFF_B|Q1 I3|B1_SYNC  2.067833848e-12
LI3|_XOR|A1 I3|A2 I3|_XOR|A1  2.067833848e-12
LI3|_XOR|A2 I3|_XOR|A1 I3|_XOR|A2  4.135667696e-12
LI3|_XOR|A3 I3|_XOR|A3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|B1 I3|B2 I3|_XOR|B1  2.067833848e-12
LI3|_XOR|B2 I3|_XOR|B1 I3|_XOR|B2  4.135667696e-12
LI3|_XOR|B3 I3|_XOR|B3 I3|_XOR|AB  8.271335392e-12
LI3|_XOR|T1 T03 I3|_XOR|T1  2.067833848e-12
LI3|_XOR|T2 I3|_XOR|T1 I3|_XOR|T2  4.135667696e-12
LI3|_XOR|Q2 I3|_XOR|ABTQ I3|_XOR|Q1  4.135667696e-12
LI3|_XOR|Q1 I3|_XOR|Q1 IP3_0  2.067833848e-12
LI3|_AND|A1 I3|A1_SYNC I3|_AND|A1  2.067833848e-12
LI3|_AND|A2 I3|_AND|A1 I3|_AND|A2  4.135667696e-12
LI3|_AND|A3 I3|_AND|A3 I3|_AND|Q3  1.2e-12
LI3|_AND|B1 I3|B1_SYNC I3|_AND|B1  2.067833848e-12
LI3|_AND|B2 I3|_AND|B1 I3|_AND|B2  4.135667696e-12
LI3|_AND|B3 I3|_AND|B3 I3|_AND|Q3  1.2e-12
LI3|_AND|Q3 I3|_AND|Q3 I3|_AND|Q2  4.135667696e-12
LI3|_AND|Q2 I3|_AND|Q2 I3|_AND|Q1  4.135667696e-12
LI3|_AND|Q1 I3|_AND|Q1 IG3_0  2.067833848e-12
LSPL_IG0_0|I_D1|B SPL_IG0_0|D1 SPL_IG0_0|I_D1|MID  2e-12
ISPL_IG0_0|I_D1|B 0 SPL_IG0_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_D2|B SPL_IG0_0|D2 SPL_IG0_0|I_D2|MID  2e-12
ISPL_IG0_0|I_D2|B 0 SPL_IG0_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG0_0|I_Q1|B SPL_IG0_0|QA1 SPL_IG0_0|I_Q1|MID  2e-12
ISPL_IG0_0|I_Q1|B 0 SPL_IG0_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG0_0|I_Q2|B SPL_IG0_0|QB1 SPL_IG0_0|I_Q2|MID  2e-12
ISPL_IG0_0|I_Q2|B 0 SPL_IG0_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG0_0|1|1 SPL_IG0_0|D1 SPL_IG0_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|1|P SPL_IG0_0|1|MID_SERIES 0  2e-13
RSPL_IG0_0|1|B SPL_IG0_0|D1 SPL_IG0_0|1|MID_SHUNT  2.7439617672
LSPL_IG0_0|1|RB SPL_IG0_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|2|1 SPL_IG0_0|D2 SPL_IG0_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|2|P SPL_IG0_0|2|MID_SERIES 0  2e-13
RSPL_IG0_0|2|B SPL_IG0_0|D2 SPL_IG0_0|2|MID_SHUNT  2.7439617672
LSPL_IG0_0|2|RB SPL_IG0_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|A|1 SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|A|P SPL_IG0_0|A|MID_SERIES 0  2e-13
RSPL_IG0_0|A|B SPL_IG0_0|QA1 SPL_IG0_0|A|MID_SHUNT  2.7439617672
LSPL_IG0_0|A|RB SPL_IG0_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG0_0|B|1 SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG0_0|B|P SPL_IG0_0|B|MID_SERIES 0  2e-13
RSPL_IG0_0|B|B SPL_IG0_0|QB1 SPL_IG0_0|B|MID_SHUNT  2.7439617672
LSPL_IG0_0|B|RB SPL_IG0_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP1_0|I_D1|B SPL_IP1_0|D1 SPL_IP1_0|I_D1|MID  2e-12
ISPL_IP1_0|I_D1|B 0 SPL_IP1_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_D2|B SPL_IP1_0|D2 SPL_IP1_0|I_D2|MID  2e-12
ISPL_IP1_0|I_D2|B 0 SPL_IP1_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP1_0|I_Q1|B SPL_IP1_0|QA1 SPL_IP1_0|I_Q1|MID  2e-12
ISPL_IP1_0|I_Q1|B 0 SPL_IP1_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP1_0|I_Q2|B SPL_IP1_0|QB1 SPL_IP1_0|I_Q2|MID  2e-12
ISPL_IP1_0|I_Q2|B 0 SPL_IP1_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP1_0|1|1 SPL_IP1_0|D1 SPL_IP1_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|1|P SPL_IP1_0|1|MID_SERIES 0  2e-13
RSPL_IP1_0|1|B SPL_IP1_0|D1 SPL_IP1_0|1|MID_SHUNT  2.7439617672
LSPL_IP1_0|1|RB SPL_IP1_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|2|1 SPL_IP1_0|D2 SPL_IP1_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|2|P SPL_IP1_0|2|MID_SERIES 0  2e-13
RSPL_IP1_0|2|B SPL_IP1_0|D2 SPL_IP1_0|2|MID_SHUNT  2.7439617672
LSPL_IP1_0|2|RB SPL_IP1_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|A|1 SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|A|P SPL_IP1_0|A|MID_SERIES 0  2e-13
RSPL_IP1_0|A|B SPL_IP1_0|QA1 SPL_IP1_0|A|MID_SHUNT  2.7439617672
LSPL_IP1_0|A|RB SPL_IP1_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP1_0|B|1 SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP1_0|B|P SPL_IP1_0|B|MID_SERIES 0  2e-13
RSPL_IP1_0|B|B SPL_IP1_0|QB1 SPL_IP1_0|B|MID_SHUNT  2.7439617672
LSPL_IP1_0|B|RB SPL_IP1_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|1 IP2_0 SPL_IP2_0|SPL1|D1  2e-12
LSPL_IP2_0|SPL1|2 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|D2  4.135667696e-12
LSPL_IP2_0|SPL1|3 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL1|4 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL1|5 SPL_IP2_0|SPL1|QA1 IP2_0_TO2  2e-12
LSPL_IP2_0|SPL1|6 SPL_IP2_0|SPL1|JCT SPL_IP2_0|SPL1|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL1|7 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|QTMP  2e-12
LSPL_IP2_0|SPL2|1 SPL_IP2_0|QTMP SPL_IP2_0|SPL2|D1  2e-12
LSPL_IP2_0|SPL2|2 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|D2  4.135667696e-12
LSPL_IP2_0|SPL2|3 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|JCT  9.84682784761905e-13
LSPL_IP2_0|SPL2|4 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QA1  9.84682784761905e-13
LSPL_IP2_0|SPL2|5 SPL_IP2_0|SPL2|QA1 IP2_0_TO3  2e-12
LSPL_IP2_0|SPL2|6 SPL_IP2_0|SPL2|JCT SPL_IP2_0|SPL2|QB1  9.84682784761905e-13
LSPL_IP2_0|SPL2|7 SPL_IP2_0|SPL2|QB1 IP2_0_OUT  2e-12
LSPL_IG2_0|I_D1|B SPL_IG2_0|D1 SPL_IG2_0|I_D1|MID  2e-12
ISPL_IG2_0|I_D1|B 0 SPL_IG2_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_D2|B SPL_IG2_0|D2 SPL_IG2_0|I_D2|MID  2e-12
ISPL_IG2_0|I_D2|B 0 SPL_IG2_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IG2_0|I_Q1|B SPL_IG2_0|QA1 SPL_IG2_0|I_Q1|MID  2e-12
ISPL_IG2_0|I_Q1|B 0 SPL_IG2_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IG2_0|I_Q2|B SPL_IG2_0|QB1 SPL_IG2_0|I_Q2|MID  2e-12
ISPL_IG2_0|I_Q2|B 0 SPL_IG2_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IG2_0|1|1 SPL_IG2_0|D1 SPL_IG2_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|1|P SPL_IG2_0|1|MID_SERIES 0  2e-13
RSPL_IG2_0|1|B SPL_IG2_0|D1 SPL_IG2_0|1|MID_SHUNT  2.7439617672
LSPL_IG2_0|1|RB SPL_IG2_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|2|1 SPL_IG2_0|D2 SPL_IG2_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|2|P SPL_IG2_0|2|MID_SERIES 0  2e-13
RSPL_IG2_0|2|B SPL_IG2_0|D2 SPL_IG2_0|2|MID_SHUNT  2.7439617672
LSPL_IG2_0|2|RB SPL_IG2_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|A|1 SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|A|P SPL_IG2_0|A|MID_SERIES 0  2e-13
RSPL_IG2_0|A|B SPL_IG2_0|QA1 SPL_IG2_0|A|MID_SHUNT  2.7439617672
LSPL_IG2_0|A|RB SPL_IG2_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IG2_0|B|1 SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IG2_0|B|P SPL_IG2_0|B|MID_SERIES 0  2e-13
RSPL_IG2_0|B|B SPL_IG2_0|QB1 SPL_IG2_0|B|MID_SHUNT  2.7439617672
LSPL_IG2_0|B|RB SPL_IG2_0|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP3_0|I_D1|B SPL_IP3_0|D1 SPL_IP3_0|I_D1|MID  2e-12
ISPL_IP3_0|I_D1|B 0 SPL_IP3_0|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_D2|B SPL_IP3_0|D2 SPL_IP3_0|I_D2|MID  2e-12
ISPL_IP3_0|I_D2|B 0 SPL_IP3_0|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LSPL_IP3_0|I_Q1|B SPL_IP3_0|QA1 SPL_IP3_0|I_Q1|MID  2e-12
ISPL_IP3_0|I_Q1|B 0 SPL_IP3_0|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LSPL_IP3_0|I_Q2|B SPL_IP3_0|QB1 SPL_IP3_0|I_Q2|MID  2e-12
ISPL_IP3_0|I_Q2|B 0 SPL_IP3_0|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BSPL_IP3_0|1|1 SPL_IP3_0|D1 SPL_IP3_0|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|1|P SPL_IP3_0|1|MID_SERIES 0  2e-13
RSPL_IP3_0|1|B SPL_IP3_0|D1 SPL_IP3_0|1|MID_SHUNT  2.7439617672
LSPL_IP3_0|1|RB SPL_IP3_0|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|2|1 SPL_IP3_0|D2 SPL_IP3_0|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|2|P SPL_IP3_0|2|MID_SERIES 0  2e-13
RSPL_IP3_0|2|B SPL_IP3_0|D2 SPL_IP3_0|2|MID_SHUNT  2.7439617672
LSPL_IP3_0|2|RB SPL_IP3_0|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|A|1 SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|A|P SPL_IP3_0|A|MID_SERIES 0  2e-13
RSPL_IP3_0|A|B SPL_IP3_0|QA1 SPL_IP3_0|A|MID_SHUNT  2.7439617672
LSPL_IP3_0|A|RB SPL_IP3_0|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP3_0|B|1 SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP3_0|B|P SPL_IP3_0|B|MID_SERIES 0  2e-13
RSPL_IP3_0|B|B SPL_IP3_0|QB1 SPL_IP3_0|B|MID_SHUNT  2.7439617672
LSPL_IP3_0|B|RB SPL_IP3_0|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|1 IP0_0 _PG0_01|P|A1  2.067833848e-12
L_PG0_01|P|2 _PG0_01|P|A1 _PG0_01|P|A2  4.135667696e-12
L_PG0_01|P|3 _PG0_01|P|A3 _PG0_01|P|A4  8.271335392e-12
L_PG0_01|P|T T04 _PG0_01|P|T1  2.067833848e-12
L_PG0_01|P|4 _PG0_01|P|T1 _PG0_01|P|T2  4.135667696e-12
L_PG0_01|P|5 _PG0_01|P|A4 _PG0_01|P|Q1  4.135667696e-12
L_PG0_01|P|6 _PG0_01|P|Q1 P0_1  2.067833848e-12
L_PG0_01|G|1 IG0_0_TO0 _PG0_01|G|A1  2.067833848e-12
L_PG0_01|G|2 _PG0_01|G|A1 _PG0_01|G|A2  4.135667696e-12
L_PG0_01|G|3 _PG0_01|G|A3 _PG0_01|G|A4  8.271335392e-12
L_PG0_01|G|T T04 _PG0_01|G|T1  2.067833848e-12
L_PG0_01|G|4 _PG0_01|G|T1 _PG0_01|G|T2  4.135667696e-12
L_PG0_01|G|5 _PG0_01|G|A4 _PG0_01|G|Q1  4.135667696e-12
L_PG0_01|G|6 _PG0_01|G|Q1 G0_1  2.067833848e-12
L_PG1_01|_SPL_G1|1 IG1_0 _PG1_01|_SPL_G1|D1  2e-12
L_PG1_01|_SPL_G1|2 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|D2  4.135667696e-12
L_PG1_01|_SPL_G1|3 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG1_01|_SPL_G1|4 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG1_01|_SPL_G1|5 _PG1_01|_SPL_G1|QA1 _PG1_01|G1_COPY_1  2e-12
L_PG1_01|_SPL_G1|6 _PG1_01|_SPL_G1|JCT _PG1_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG1_01|_SPL_G1|7 _PG1_01|_SPL_G1|QB1 _PG1_01|G1_COPY_2  2e-12
L_PG1_01|_PG|A1 IP1_0_TO1 _PG1_01|_PG|A1  2.067833848e-12
L_PG1_01|_PG|A2 _PG1_01|_PG|A1 _PG1_01|_PG|A2  4.135667696e-12
L_PG1_01|_PG|A3 _PG1_01|_PG|A3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|B1 _PG1_01|G1_COPY_1 _PG1_01|_PG|B1  2.067833848e-12
L_PG1_01|_PG|B2 _PG1_01|_PG|B1 _PG1_01|_PG|B2  4.135667696e-12
L_PG1_01|_PG|B3 _PG1_01|_PG|B3 _PG1_01|_PG|Q3  1.2e-12
L_PG1_01|_PG|Q3 _PG1_01|_PG|Q3 _PG1_01|_PG|Q2  4.135667696e-12
L_PG1_01|_PG|Q2 _PG1_01|_PG|Q2 _PG1_01|_PG|Q1  4.135667696e-12
L_PG1_01|_PG|Q1 _PG1_01|_PG|Q1 _PG1_01|PG  2.067833848e-12
L_PG1_01|_GG|A1 IG0_0_TO1 _PG1_01|_GG|A1  2.067833848e-12
L_PG1_01|_GG|A2 _PG1_01|_GG|A1 _PG1_01|_GG|A2  4.135667696e-12
L_PG1_01|_GG|A3 _PG1_01|_GG|A3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|B1 _PG1_01|G1_COPY_2 _PG1_01|_GG|B1  2.067833848e-12
L_PG1_01|_GG|B2 _PG1_01|_GG|B1 _PG1_01|_GG|B2  4.135667696e-12
L_PG1_01|_GG|B3 _PG1_01|_GG|B3 _PG1_01|_GG|Q3  1.2e-12
L_PG1_01|_GG|Q3 _PG1_01|_GG|Q3 _PG1_01|_GG|Q2  4.135667696e-12
L_PG1_01|_GG|Q2 _PG1_01|_GG|Q2 _PG1_01|_GG|Q1  4.135667696e-12
L_PG1_01|_GG|Q1 _PG1_01|_GG|Q1 _PG1_01|GG  2.067833848e-12
L_PG1_01|_DFF_PG|1 _PG1_01|PG _PG1_01|_DFF_PG|A1  2.067833848e-12
L_PG1_01|_DFF_PG|2 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|A2  4.135667696e-12
L_PG1_01|_DFF_PG|3 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|A4  8.271335392e-12
L_PG1_01|_DFF_PG|T T05 _PG1_01|_DFF_PG|T1  2.067833848e-12
L_PG1_01|_DFF_PG|4 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T2  4.135667696e-12
L_PG1_01|_DFF_PG|5 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|Q1  4.135667696e-12
L_PG1_01|_DFF_PG|6 _PG1_01|_DFF_PG|Q1 _PG1_01|PG_SYNC  2.067833848e-12
L_PG1_01|_DFF_GG|1 _PG1_01|GG _PG1_01|_DFF_GG|A1  2.067833848e-12
L_PG1_01|_DFF_GG|2 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|A2  4.135667696e-12
L_PG1_01|_DFF_GG|3 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|A4  8.271335392e-12
L_PG1_01|_DFF_GG|T T05 _PG1_01|_DFF_GG|T1  2.067833848e-12
L_PG1_01|_DFF_GG|4 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T2  4.135667696e-12
L_PG1_01|_DFF_GG|5 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|Q1  4.135667696e-12
L_PG1_01|_DFF_GG|6 _PG1_01|_DFF_GG|Q1 _PG1_01|GG_SYNC  2.067833848e-12
L_PG1_01|_AND_G|A1 _PG1_01|PG_SYNC _PG1_01|_AND_G|A1  2.067833848e-12
L_PG1_01|_AND_G|A2 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A2  4.135667696e-12
L_PG1_01|_AND_G|A3 _PG1_01|_AND_G|A3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|B1 _PG1_01|GG_SYNC _PG1_01|_AND_G|B1  2.067833848e-12
L_PG1_01|_AND_G|B2 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B2  4.135667696e-12
L_PG1_01|_AND_G|B3 _PG1_01|_AND_G|B3 _PG1_01|_AND_G|Q3  1.2e-12
L_PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|Q2  4.135667696e-12
L_PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q1  4.135667696e-12
L_PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1 G1_1  2.067833848e-12
L_PG2_01|P|1 IP2_0_TO2 _PG2_01|P|A1  2.067833848e-12
L_PG2_01|P|2 _PG2_01|P|A1 _PG2_01|P|A2  4.135667696e-12
L_PG2_01|P|3 _PG2_01|P|A3 _PG2_01|P|A4  8.271335392e-12
L_PG2_01|P|T T06 _PG2_01|P|T1  2.067833848e-12
L_PG2_01|P|4 _PG2_01|P|T1 _PG2_01|P|T2  4.135667696e-12
L_PG2_01|P|5 _PG2_01|P|A4 _PG2_01|P|Q1  4.135667696e-12
L_PG2_01|P|6 _PG2_01|P|Q1 P2_1  2.067833848e-12
L_PG2_01|G|1 IG2_0_TO2 _PG2_01|G|A1  2.067833848e-12
L_PG2_01|G|2 _PG2_01|G|A1 _PG2_01|G|A2  4.135667696e-12
L_PG2_01|G|3 _PG2_01|G|A3 _PG2_01|G|A4  8.271335392e-12
L_PG2_01|G|T T06 _PG2_01|G|T1  2.067833848e-12
L_PG2_01|G|4 _PG2_01|G|T1 _PG2_01|G|T2  4.135667696e-12
L_PG2_01|G|5 _PG2_01|G|A4 _PG2_01|G|Q1  4.135667696e-12
L_PG2_01|G|6 _PG2_01|G|Q1 G2_1  2.067833848e-12
L_PG3_01|_SPL_G1|1 IG3_0 _PG3_01|_SPL_G1|D1  2e-12
L_PG3_01|_SPL_G1|2 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|D2  4.135667696e-12
L_PG3_01|_SPL_G1|3 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_G1|4 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_G1|5 _PG3_01|_SPL_G1|QA1 _PG3_01|G1_COPY_1  2e-12
L_PG3_01|_SPL_G1|6 _PG3_01|_SPL_G1|JCT _PG3_01|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_G1|7 _PG3_01|_SPL_G1|QB1 _PG3_01|G1_COPY_2  2e-12
L_PG3_01|_SPL_P1|1 IP3_0_TO1 _PG3_01|_SPL_P1|D1  2e-12
L_PG3_01|_SPL_P1|2 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|D2  4.135667696e-12
L_PG3_01|_SPL_P1|3 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|JCT  9.84682784761905e-13
L_PG3_01|_SPL_P1|4 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QA1  9.84682784761905e-13
L_PG3_01|_SPL_P1|5 _PG3_01|_SPL_P1|QA1 _PG3_01|P1_COPY_1  2e-12
L_PG3_01|_SPL_P1|6 _PG3_01|_SPL_P1|JCT _PG3_01|_SPL_P1|QB1  9.84682784761905e-13
L_PG3_01|_SPL_P1|7 _PG3_01|_SPL_P1|QB1 _PG3_01|P1_COPY_2  2e-12
L_PG3_01|_PG|A1 _PG3_01|P1_COPY_1 _PG3_01|_PG|A1  2.067833848e-12
L_PG3_01|_PG|A2 _PG3_01|_PG|A1 _PG3_01|_PG|A2  4.135667696e-12
L_PG3_01|_PG|A3 _PG3_01|_PG|A3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|B1 _PG3_01|G1_COPY_1 _PG3_01|_PG|B1  2.067833848e-12
L_PG3_01|_PG|B2 _PG3_01|_PG|B1 _PG3_01|_PG|B2  4.135667696e-12
L_PG3_01|_PG|B3 _PG3_01|_PG|B3 _PG3_01|_PG|Q3  1.2e-12
L_PG3_01|_PG|Q3 _PG3_01|_PG|Q3 _PG3_01|_PG|Q2  4.135667696e-12
L_PG3_01|_PG|Q2 _PG3_01|_PG|Q2 _PG3_01|_PG|Q1  4.135667696e-12
L_PG3_01|_PG|Q1 _PG3_01|_PG|Q1 _PG3_01|PG  2.067833848e-12
L_PG3_01|_GG|A1 IG2_0_TO3 _PG3_01|_GG|A1  2.067833848e-12
L_PG3_01|_GG|A2 _PG3_01|_GG|A1 _PG3_01|_GG|A2  4.135667696e-12
L_PG3_01|_GG|A3 _PG3_01|_GG|A3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|B1 _PG3_01|G1_COPY_2 _PG3_01|_GG|B1  2.067833848e-12
L_PG3_01|_GG|B2 _PG3_01|_GG|B1 _PG3_01|_GG|B2  4.135667696e-12
L_PG3_01|_GG|B3 _PG3_01|_GG|B3 _PG3_01|_GG|Q3  1.2e-12
L_PG3_01|_GG|Q3 _PG3_01|_GG|Q3 _PG3_01|_GG|Q2  4.135667696e-12
L_PG3_01|_GG|Q2 _PG3_01|_GG|Q2 _PG3_01|_GG|Q1  4.135667696e-12
L_PG3_01|_GG|Q1 _PG3_01|_GG|Q1 _PG3_01|GG  2.067833848e-12
L_PG3_01|_DFF_P0|1 IP2_0_TO3 _PG3_01|_DFF_P0|A1  2.067833848e-12
L_PG3_01|_DFF_P0|2 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|A2  4.135667696e-12
L_PG3_01|_DFF_P0|3 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|A4  8.271335392e-12
L_PG3_01|_DFF_P0|T T07 _PG3_01|_DFF_P0|T1  2.067833848e-12
L_PG3_01|_DFF_P0|4 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T2  4.135667696e-12
L_PG3_01|_DFF_P0|5 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|Q1  4.135667696e-12
L_PG3_01|_DFF_P0|6 _PG3_01|_DFF_P0|Q1 _PG3_01|P0_SYNC  2.067833848e-12
L_PG3_01|_DFF_P1|1 _PG3_01|P1_COPY_2 _PG3_01|_DFF_P1|A1  2.067833848e-12
L_PG3_01|_DFF_P1|2 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|A2  4.135667696e-12
L_PG3_01|_DFF_P1|3 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|A4  8.271335392e-12
L_PG3_01|_DFF_P1|T T07 _PG3_01|_DFF_P1|T1  2.067833848e-12
L_PG3_01|_DFF_P1|4 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T2  4.135667696e-12
L_PG3_01|_DFF_P1|5 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|Q1  4.135667696e-12
L_PG3_01|_DFF_P1|6 _PG3_01|_DFF_P1|Q1 _PG3_01|P1_SYNC  2.067833848e-12
L_PG3_01|_DFF_PG|1 _PG3_01|PG _PG3_01|_DFF_PG|A1  2.067833848e-12
L_PG3_01|_DFF_PG|2 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|A2  4.135667696e-12
L_PG3_01|_DFF_PG|3 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|A4  8.271335392e-12
L_PG3_01|_DFF_PG|T T07 _PG3_01|_DFF_PG|T1  2.067833848e-12
L_PG3_01|_DFF_PG|4 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T2  4.135667696e-12
L_PG3_01|_DFF_PG|5 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|Q1  4.135667696e-12
L_PG3_01|_DFF_PG|6 _PG3_01|_DFF_PG|Q1 _PG3_01|PG_SYNC  2.067833848e-12
L_PG3_01|_DFF_GG|1 _PG3_01|GG _PG3_01|_DFF_GG|A1  2.067833848e-12
L_PG3_01|_DFF_GG|2 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|A2  4.135667696e-12
L_PG3_01|_DFF_GG|3 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|A4  8.271335392e-12
L_PG3_01|_DFF_GG|T T07 _PG3_01|_DFF_GG|T1  2.067833848e-12
L_PG3_01|_DFF_GG|4 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T2  4.135667696e-12
L_PG3_01|_DFF_GG|5 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|Q1  4.135667696e-12
L_PG3_01|_DFF_GG|6 _PG3_01|_DFF_GG|Q1 _PG3_01|GG_SYNC  2.067833848e-12
L_PG3_01|_AND_G|A1 _PG3_01|PG_SYNC _PG3_01|_AND_G|A1  2.067833848e-12
L_PG3_01|_AND_G|A2 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A2  4.135667696e-12
L_PG3_01|_AND_G|A3 _PG3_01|_AND_G|A3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|B1 _PG3_01|GG_SYNC _PG3_01|_AND_G|B1  2.067833848e-12
L_PG3_01|_AND_G|B2 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B2  4.135667696e-12
L_PG3_01|_AND_G|B3 _PG3_01|_AND_G|B3 _PG3_01|_AND_G|Q3  1.2e-12
L_PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|Q2  4.135667696e-12
L_PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q1  4.135667696e-12
L_PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1 G3_1  2.067833848e-12
L_PG3_01|_AND_P|A1 _PG3_01|P0_SYNC _PG3_01|_AND_P|A1  2.067833848e-12
L_PG3_01|_AND_P|A2 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A2  4.135667696e-12
L_PG3_01|_AND_P|A3 _PG3_01|_AND_P|A3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|B1 _PG3_01|P1_SYNC _PG3_01|_AND_P|B1  2.067833848e-12
L_PG3_01|_AND_P|B2 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B2  4.135667696e-12
L_PG3_01|_AND_P|B3 _PG3_01|_AND_P|B3 _PG3_01|_AND_P|Q3  1.2e-12
L_PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|Q2  4.135667696e-12
L_PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q1  4.135667696e-12
L_PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1 P3_1  2.067833848e-12
L_DFF_IP1_01|I_1|B _DFF_IP1_01|A1 _DFF_IP1_01|I_1|MID  2e-12
I_DFF_IP1_01|I_1|B 0 _DFF_IP1_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_3|B _DFF_IP1_01|A3 _DFF_IP1_01|I_3|MID  2e-12
I_DFF_IP1_01|I_3|B 0 _DFF_IP1_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_01|I_T|B _DFF_IP1_01|T1 _DFF_IP1_01|I_T|MID  2e-12
I_DFF_IP1_01|I_T|B 0 _DFF_IP1_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_01|I_6|B _DFF_IP1_01|Q1 _DFF_IP1_01|I_6|MID  2e-12
I_DFF_IP1_01|I_6|B 0 _DFF_IP1_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_01|1|1 _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|1|P _DFF_IP1_01|1|MID_SERIES 0  2e-13
R_DFF_IP1_01|1|B _DFF_IP1_01|A1 _DFF_IP1_01|1|MID_SHUNT  2.7439617672
L_DFF_IP1_01|1|RB _DFF_IP1_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|23|1 _DFF_IP1_01|A2 _DFF_IP1_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|23|B _DFF_IP1_01|A2 _DFF_IP1_01|23|MID_SHUNT  3.84154647408
L_DFF_IP1_01|23|RB _DFF_IP1_01|23|MID_SHUNT _DFF_IP1_01|A3  2.1704737578552e-12
B_DFF_IP1_01|3|1 _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|3|P _DFF_IP1_01|3|MID_SERIES 0  2e-13
R_DFF_IP1_01|3|B _DFF_IP1_01|A3 _DFF_IP1_01|3|MID_SHUNT  2.7439617672
L_DFF_IP1_01|3|RB _DFF_IP1_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|4|1 _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|4|P _DFF_IP1_01|4|MID_SERIES 0  2e-13
R_DFF_IP1_01|4|B _DFF_IP1_01|A4 _DFF_IP1_01|4|MID_SHUNT  2.7439617672
L_DFF_IP1_01|4|RB _DFF_IP1_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|T|1 _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|T|P _DFF_IP1_01|T|MID_SERIES 0  2e-13
R_DFF_IP1_01|T|B _DFF_IP1_01|T1 _DFF_IP1_01|T|MID_SHUNT  2.7439617672
L_DFF_IP1_01|T|RB _DFF_IP1_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_01|45|1 _DFF_IP1_01|T2 _DFF_IP1_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_01|45|B _DFF_IP1_01|T2 _DFF_IP1_01|45|MID_SHUNT  3.84154647408
L_DFF_IP1_01|45|RB _DFF_IP1_01|45|MID_SHUNT _DFF_IP1_01|A4  2.1704737578552e-12
B_DFF_IP1_01|6|1 _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_01|6|P _DFF_IP1_01|6|MID_SERIES 0  2e-13
R_DFF_IP1_01|6|B _DFF_IP1_01|Q1 _DFF_IP1_01|6|MID_SHUNT  2.7439617672
L_DFF_IP1_01|6|RB _DFF_IP1_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_01|I_1|B _DFF_IP2_01|A1 _DFF_IP2_01|I_1|MID  2e-12
I_DFF_IP2_01|I_1|B 0 _DFF_IP2_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_3|B _DFF_IP2_01|A3 _DFF_IP2_01|I_3|MID  2e-12
I_DFF_IP2_01|I_3|B 0 _DFF_IP2_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_01|I_T|B _DFF_IP2_01|T1 _DFF_IP2_01|I_T|MID  2e-12
I_DFF_IP2_01|I_T|B 0 _DFF_IP2_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_01|I_6|B _DFF_IP2_01|Q1 _DFF_IP2_01|I_6|MID  2e-12
I_DFF_IP2_01|I_6|B 0 _DFF_IP2_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_01|1|1 _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|1|P _DFF_IP2_01|1|MID_SERIES 0  2e-13
R_DFF_IP2_01|1|B _DFF_IP2_01|A1 _DFF_IP2_01|1|MID_SHUNT  2.7439617672
L_DFF_IP2_01|1|RB _DFF_IP2_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|23|1 _DFF_IP2_01|A2 _DFF_IP2_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|23|B _DFF_IP2_01|A2 _DFF_IP2_01|23|MID_SHUNT  3.84154647408
L_DFF_IP2_01|23|RB _DFF_IP2_01|23|MID_SHUNT _DFF_IP2_01|A3  2.1704737578552e-12
B_DFF_IP2_01|3|1 _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|3|P _DFF_IP2_01|3|MID_SERIES 0  2e-13
R_DFF_IP2_01|3|B _DFF_IP2_01|A3 _DFF_IP2_01|3|MID_SHUNT  2.7439617672
L_DFF_IP2_01|3|RB _DFF_IP2_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|4|1 _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|4|P _DFF_IP2_01|4|MID_SERIES 0  2e-13
R_DFF_IP2_01|4|B _DFF_IP2_01|A4 _DFF_IP2_01|4|MID_SHUNT  2.7439617672
L_DFF_IP2_01|4|RB _DFF_IP2_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|T|1 _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|T|P _DFF_IP2_01|T|MID_SERIES 0  2e-13
R_DFF_IP2_01|T|B _DFF_IP2_01|T1 _DFF_IP2_01|T|MID_SHUNT  2.7439617672
L_DFF_IP2_01|T|RB _DFF_IP2_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_01|45|1 _DFF_IP2_01|T2 _DFF_IP2_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_01|45|B _DFF_IP2_01|T2 _DFF_IP2_01|45|MID_SHUNT  3.84154647408
L_DFF_IP2_01|45|RB _DFF_IP2_01|45|MID_SHUNT _DFF_IP2_01|A4  2.1704737578552e-12
B_DFF_IP2_01|6|1 _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_01|6|P _DFF_IP2_01|6|MID_SERIES 0  2e-13
R_DFF_IP2_01|6|B _DFF_IP2_01|Q1 _DFF_IP2_01|6|MID_SHUNT  2.7439617672
L_DFF_IP2_01|6|RB _DFF_IP2_01|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_01|I_1|B _DFF_IP3_01|A1 _DFF_IP3_01|I_1|MID  2e-12
I_DFF_IP3_01|I_1|B 0 _DFF_IP3_01|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_3|B _DFF_IP3_01|A3 _DFF_IP3_01|I_3|MID  2e-12
I_DFF_IP3_01|I_3|B 0 _DFF_IP3_01|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_01|I_T|B _DFF_IP3_01|T1 _DFF_IP3_01|I_T|MID  2e-12
I_DFF_IP3_01|I_T|B 0 _DFF_IP3_01|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_01|I_6|B _DFF_IP3_01|Q1 _DFF_IP3_01|I_6|MID  2e-12
I_DFF_IP3_01|I_6|B 0 _DFF_IP3_01|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_01|1|1 _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|1|P _DFF_IP3_01|1|MID_SERIES 0  2e-13
R_DFF_IP3_01|1|B _DFF_IP3_01|A1 _DFF_IP3_01|1|MID_SHUNT  2.7439617672
L_DFF_IP3_01|1|RB _DFF_IP3_01|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|23|1 _DFF_IP3_01|A2 _DFF_IP3_01|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|23|B _DFF_IP3_01|A2 _DFF_IP3_01|23|MID_SHUNT  3.84154647408
L_DFF_IP3_01|23|RB _DFF_IP3_01|23|MID_SHUNT _DFF_IP3_01|A3  2.1704737578552e-12
B_DFF_IP3_01|3|1 _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|3|P _DFF_IP3_01|3|MID_SERIES 0  2e-13
R_DFF_IP3_01|3|B _DFF_IP3_01|A3 _DFF_IP3_01|3|MID_SHUNT  2.7439617672
L_DFF_IP3_01|3|RB _DFF_IP3_01|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|4|1 _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|4|P _DFF_IP3_01|4|MID_SERIES 0  2e-13
R_DFF_IP3_01|4|B _DFF_IP3_01|A4 _DFF_IP3_01|4|MID_SHUNT  2.7439617672
L_DFF_IP3_01|4|RB _DFF_IP3_01|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|T|1 _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|T|P _DFF_IP3_01|T|MID_SERIES 0  2e-13
R_DFF_IP3_01|T|B _DFF_IP3_01|T1 _DFF_IP3_01|T|MID_SHUNT  2.7439617672
L_DFF_IP3_01|T|RB _DFF_IP3_01|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_01|45|1 _DFF_IP3_01|T2 _DFF_IP3_01|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_01|45|B _DFF_IP3_01|T2 _DFF_IP3_01|45|MID_SHUNT  3.84154647408
L_DFF_IP3_01|45|RB _DFF_IP3_01|45|MID_SHUNT _DFF_IP3_01|A4  2.1704737578552e-12
B_DFF_IP3_01|6|1 _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_01|6|P _DFF_IP3_01|6|MID_SERIES 0  2e-13
R_DFF_IP3_01|6|B _DFF_IP3_01|Q1 _DFF_IP3_01|6|MID_SHUNT  2.7439617672
L_DFF_IP3_01|6|RB _DFF_IP3_01|6|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL1|1 G1_1 SPL_G1_1|SPL1|D1  2e-12
LSPL_G1_1|SPL1|2 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|D2  4.135667696e-12
LSPL_G1_1|SPL1|3 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|JCT  9.84682784761905e-13
LSPL_G1_1|SPL1|4 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QA1  9.84682784761905e-13
LSPL_G1_1|SPL1|5 SPL_G1_1|SPL1|QA1 G1_1_TO1  2e-12
LSPL_G1_1|SPL1|6 SPL_G1_1|SPL1|JCT SPL_G1_1|SPL1|QB1  9.84682784761905e-13
LSPL_G1_1|SPL1|7 SPL_G1_1|SPL1|QB1 SPL_G1_1|QTMP  2e-12
LSPL_G1_1|SPL2|1 SPL_G1_1|QTMP SPL_G1_1|SPL2|D1  2e-12
LSPL_G1_1|SPL2|2 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|D2  4.135667696e-12
LSPL_G1_1|SPL2|3 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|JCT  9.84682784761905e-13
LSPL_G1_1|SPL2|4 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QA1  9.84682784761905e-13
LSPL_G1_1|SPL2|5 SPL_G1_1|SPL2|QA1 G1_1_TO2  2e-12
LSPL_G1_1|SPL2|6 SPL_G1_1|SPL2|JCT SPL_G1_1|SPL2|QB1  9.84682784761905e-13
LSPL_G1_1|SPL2|7 SPL_G1_1|SPL2|QB1 G1_1_TO3  2e-12
L_PG0_12|P|1 P0_1 _PG0_12|P|A1  2.067833848e-12
L_PG0_12|P|2 _PG0_12|P|A1 _PG0_12|P|A2  4.135667696e-12
L_PG0_12|P|3 _PG0_12|P|A3 _PG0_12|P|A4  8.271335392e-12
L_PG0_12|P|T T08 _PG0_12|P|T1  2.067833848e-12
L_PG0_12|P|4 _PG0_12|P|T1 _PG0_12|P|T2  4.135667696e-12
L_PG0_12|P|5 _PG0_12|P|A4 _PG0_12|P|Q1  4.135667696e-12
L_PG0_12|P|6 _PG0_12|P|Q1 P0_2  2.067833848e-12
L_PG0_12|G|1 G0_1 _PG0_12|G|A1  2.067833848e-12
L_PG0_12|G|2 _PG0_12|G|A1 _PG0_12|G|A2  4.135667696e-12
L_PG0_12|G|3 _PG0_12|G|A3 _PG0_12|G|A4  8.271335392e-12
L_PG0_12|G|T T08 _PG0_12|G|T1  2.067833848e-12
L_PG0_12|G|4 _PG0_12|G|T1 _PG0_12|G|T2  4.135667696e-12
L_PG0_12|G|5 _PG0_12|G|A4 _PG0_12|G|Q1  4.135667696e-12
L_PG0_12|G|6 _PG0_12|G|Q1 G0_2  2.067833848e-12
L_PG1_12|I_1|B _PG1_12|A1 _PG1_12|I_1|MID  2e-12
I_PG1_12|I_1|B 0 _PG1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_3|B _PG1_12|A3 _PG1_12|I_3|MID  2e-12
I_PG1_12|I_3|B 0 _PG1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_12|I_T|B _PG1_12|T1 _PG1_12|I_T|MID  2e-12
I_PG1_12|I_T|B 0 _PG1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_12|I_6|B _PG1_12|Q1 _PG1_12|I_6|MID  2e-12
I_PG1_12|I_6|B 0 _PG1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_12|1|1 _PG1_12|A1 _PG1_12|1|MID_SERIES JJMIT AREA=2.5
L_PG1_12|1|P _PG1_12|1|MID_SERIES 0  2e-13
R_PG1_12|1|B _PG1_12|A1 _PG1_12|1|MID_SHUNT  2.7439617672
L_PG1_12|1|RB _PG1_12|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|23|1 _PG1_12|A2 _PG1_12|A3 JJMIT AREA=1.7857142857142858
R_PG1_12|23|B _PG1_12|A2 _PG1_12|23|MID_SHUNT  3.84154647408
L_PG1_12|23|RB _PG1_12|23|MID_SHUNT _PG1_12|A3  2.1704737578552e-12
B_PG1_12|3|1 _PG1_12|A3 _PG1_12|3|MID_SERIES JJMIT AREA=2.5
L_PG1_12|3|P _PG1_12|3|MID_SERIES 0  2e-13
R_PG1_12|3|B _PG1_12|A3 _PG1_12|3|MID_SHUNT  2.7439617672
L_PG1_12|3|RB _PG1_12|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|4|1 _PG1_12|A4 _PG1_12|4|MID_SERIES JJMIT AREA=2.5
L_PG1_12|4|P _PG1_12|4|MID_SERIES 0  2e-13
R_PG1_12|4|B _PG1_12|A4 _PG1_12|4|MID_SHUNT  2.7439617672
L_PG1_12|4|RB _PG1_12|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|T|1 _PG1_12|T1 _PG1_12|T|MID_SERIES JJMIT AREA=2.5
L_PG1_12|T|P _PG1_12|T|MID_SERIES 0  2e-13
R_PG1_12|T|B _PG1_12|T1 _PG1_12|T|MID_SHUNT  2.7439617672
L_PG1_12|T|RB _PG1_12|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_12|45|1 _PG1_12|T2 _PG1_12|A4 JJMIT AREA=1.7857142857142858
R_PG1_12|45|B _PG1_12|T2 _PG1_12|45|MID_SHUNT  3.84154647408
L_PG1_12|45|RB _PG1_12|45|MID_SHUNT _PG1_12|A4  2.1704737578552e-12
B_PG1_12|6|1 _PG1_12|Q1 _PG1_12|6|MID_SERIES JJMIT AREA=2.5
L_PG1_12|6|P _PG1_12|6|MID_SERIES 0  2e-13
R_PG1_12|6|B _PG1_12|Q1 _PG1_12|6|MID_SHUNT  2.7439617672
L_PG1_12|6|RB _PG1_12|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|1 G2_1 _PG2_12|_SPL_G1|D1  2e-12
L_PG2_12|_SPL_G1|2 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|D2  4.135667696e-12
L_PG2_12|_SPL_G1|3 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG2_12|_SPL_G1|4 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG2_12|_SPL_G1|5 _PG2_12|_SPL_G1|QA1 _PG2_12|G1_COPY_1  2e-12
L_PG2_12|_SPL_G1|6 _PG2_12|_SPL_G1|JCT _PG2_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG2_12|_SPL_G1|7 _PG2_12|_SPL_G1|QB1 _PG2_12|G1_COPY_2  2e-12
L_PG2_12|_PG|A1 P2_1 _PG2_12|_PG|A1  2.067833848e-12
L_PG2_12|_PG|A2 _PG2_12|_PG|A1 _PG2_12|_PG|A2  4.135667696e-12
L_PG2_12|_PG|A3 _PG2_12|_PG|A3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|B1 _PG2_12|G1_COPY_1 _PG2_12|_PG|B1  2.067833848e-12
L_PG2_12|_PG|B2 _PG2_12|_PG|B1 _PG2_12|_PG|B2  4.135667696e-12
L_PG2_12|_PG|B3 _PG2_12|_PG|B3 _PG2_12|_PG|Q3  1.2e-12
L_PG2_12|_PG|Q3 _PG2_12|_PG|Q3 _PG2_12|_PG|Q2  4.135667696e-12
L_PG2_12|_PG|Q2 _PG2_12|_PG|Q2 _PG2_12|_PG|Q1  4.135667696e-12
L_PG2_12|_PG|Q1 _PG2_12|_PG|Q1 _PG2_12|PG  2.067833848e-12
L_PG2_12|_GG|A1 G1_1_TO2 _PG2_12|_GG|A1  2.067833848e-12
L_PG2_12|_GG|A2 _PG2_12|_GG|A1 _PG2_12|_GG|A2  4.135667696e-12
L_PG2_12|_GG|A3 _PG2_12|_GG|A3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|B1 _PG2_12|G1_COPY_2 _PG2_12|_GG|B1  2.067833848e-12
L_PG2_12|_GG|B2 _PG2_12|_GG|B1 _PG2_12|_GG|B2  4.135667696e-12
L_PG2_12|_GG|B3 _PG2_12|_GG|B3 _PG2_12|_GG|Q3  1.2e-12
L_PG2_12|_GG|Q3 _PG2_12|_GG|Q3 _PG2_12|_GG|Q2  4.135667696e-12
L_PG2_12|_GG|Q2 _PG2_12|_GG|Q2 _PG2_12|_GG|Q1  4.135667696e-12
L_PG2_12|_GG|Q1 _PG2_12|_GG|Q1 _PG2_12|GG  2.067833848e-12
L_PG2_12|_DFF_PG|1 _PG2_12|PG _PG2_12|_DFF_PG|A1  2.067833848e-12
L_PG2_12|_DFF_PG|2 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|A2  4.135667696e-12
L_PG2_12|_DFF_PG|3 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|A4  8.271335392e-12
L_PG2_12|_DFF_PG|T T10 _PG2_12|_DFF_PG|T1  2.067833848e-12
L_PG2_12|_DFF_PG|4 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T2  4.135667696e-12
L_PG2_12|_DFF_PG|5 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|Q1  4.135667696e-12
L_PG2_12|_DFF_PG|6 _PG2_12|_DFF_PG|Q1 _PG2_12|PG_SYNC  2.067833848e-12
L_PG2_12|_DFF_GG|1 _PG2_12|GG _PG2_12|_DFF_GG|A1  2.067833848e-12
L_PG2_12|_DFF_GG|2 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|A2  4.135667696e-12
L_PG2_12|_DFF_GG|3 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|A4  8.271335392e-12
L_PG2_12|_DFF_GG|T T10 _PG2_12|_DFF_GG|T1  2.067833848e-12
L_PG2_12|_DFF_GG|4 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T2  4.135667696e-12
L_PG2_12|_DFF_GG|5 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|Q1  4.135667696e-12
L_PG2_12|_DFF_GG|6 _PG2_12|_DFF_GG|Q1 _PG2_12|GG_SYNC  2.067833848e-12
L_PG2_12|_AND_G|A1 _PG2_12|PG_SYNC _PG2_12|_AND_G|A1  2.067833848e-12
L_PG2_12|_AND_G|A2 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A2  4.135667696e-12
L_PG2_12|_AND_G|A3 _PG2_12|_AND_G|A3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|B1 _PG2_12|GG_SYNC _PG2_12|_AND_G|B1  2.067833848e-12
L_PG2_12|_AND_G|B2 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B2  4.135667696e-12
L_PG2_12|_AND_G|B3 _PG2_12|_AND_G|B3 _PG2_12|_AND_G|Q3  1.2e-12
L_PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|Q2  4.135667696e-12
L_PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q1  4.135667696e-12
L_PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1 G2_2  2.067833848e-12
L_PG3_12|_SPL_G1|1 G3_1 _PG3_12|_SPL_G1|D1  2e-12
L_PG3_12|_SPL_G1|2 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|D2  4.135667696e-12
L_PG3_12|_SPL_G1|3 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|JCT  9.84682784761905e-13
L_PG3_12|_SPL_G1|4 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QA1  9.84682784761905e-13
L_PG3_12|_SPL_G1|5 _PG3_12|_SPL_G1|QA1 _PG3_12|G1_COPY_1  2e-12
L_PG3_12|_SPL_G1|6 _PG3_12|_SPL_G1|JCT _PG3_12|_SPL_G1|QB1  9.84682784761905e-13
L_PG3_12|_SPL_G1|7 _PG3_12|_SPL_G1|QB1 _PG3_12|G1_COPY_2  2e-12
L_PG3_12|_PG|A1 P3_1 _PG3_12|_PG|A1  2.067833848e-12
L_PG3_12|_PG|A2 _PG3_12|_PG|A1 _PG3_12|_PG|A2  4.135667696e-12
L_PG3_12|_PG|A3 _PG3_12|_PG|A3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|B1 _PG3_12|G1_COPY_1 _PG3_12|_PG|B1  2.067833848e-12
L_PG3_12|_PG|B2 _PG3_12|_PG|B1 _PG3_12|_PG|B2  4.135667696e-12
L_PG3_12|_PG|B3 _PG3_12|_PG|B3 _PG3_12|_PG|Q3  1.2e-12
L_PG3_12|_PG|Q3 _PG3_12|_PG|Q3 _PG3_12|_PG|Q2  4.135667696e-12
L_PG3_12|_PG|Q2 _PG3_12|_PG|Q2 _PG3_12|_PG|Q1  4.135667696e-12
L_PG3_12|_PG|Q1 _PG3_12|_PG|Q1 _PG3_12|PG  2.067833848e-12
L_PG3_12|_GG|A1 G1_1_TO3 _PG3_12|_GG|A1  2.067833848e-12
L_PG3_12|_GG|A2 _PG3_12|_GG|A1 _PG3_12|_GG|A2  4.135667696e-12
L_PG3_12|_GG|A3 _PG3_12|_GG|A3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|B1 _PG3_12|G1_COPY_2 _PG3_12|_GG|B1  2.067833848e-12
L_PG3_12|_GG|B2 _PG3_12|_GG|B1 _PG3_12|_GG|B2  4.135667696e-12
L_PG3_12|_GG|B3 _PG3_12|_GG|B3 _PG3_12|_GG|Q3  1.2e-12
L_PG3_12|_GG|Q3 _PG3_12|_GG|Q3 _PG3_12|_GG|Q2  4.135667696e-12
L_PG3_12|_GG|Q2 _PG3_12|_GG|Q2 _PG3_12|_GG|Q1  4.135667696e-12
L_PG3_12|_GG|Q1 _PG3_12|_GG|Q1 _PG3_12|GG  2.067833848e-12
L_PG3_12|_DFF_PG|1 _PG3_12|PG _PG3_12|_DFF_PG|A1  2.067833848e-12
L_PG3_12|_DFF_PG|2 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|A2  4.135667696e-12
L_PG3_12|_DFF_PG|3 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|A4  8.271335392e-12
L_PG3_12|_DFF_PG|T T11 _PG3_12|_DFF_PG|T1  2.067833848e-12
L_PG3_12|_DFF_PG|4 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T2  4.135667696e-12
L_PG3_12|_DFF_PG|5 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|Q1  4.135667696e-12
L_PG3_12|_DFF_PG|6 _PG3_12|_DFF_PG|Q1 _PG3_12|PG_SYNC  2.067833848e-12
L_PG3_12|_DFF_GG|1 _PG3_12|GG _PG3_12|_DFF_GG|A1  2.067833848e-12
L_PG3_12|_DFF_GG|2 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|A2  4.135667696e-12
L_PG3_12|_DFF_GG|3 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|A4  8.271335392e-12
L_PG3_12|_DFF_GG|T T11 _PG3_12|_DFF_GG|T1  2.067833848e-12
L_PG3_12|_DFF_GG|4 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T2  4.135667696e-12
L_PG3_12|_DFF_GG|5 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|Q1  4.135667696e-12
L_PG3_12|_DFF_GG|6 _PG3_12|_DFF_GG|Q1 _PG3_12|GG_SYNC  2.067833848e-12
L_PG3_12|_AND_G|A1 _PG3_12|PG_SYNC _PG3_12|_AND_G|A1  2.067833848e-12
L_PG3_12|_AND_G|A2 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A2  4.135667696e-12
L_PG3_12|_AND_G|A3 _PG3_12|_AND_G|A3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|B1 _PG3_12|GG_SYNC _PG3_12|_AND_G|B1  2.067833848e-12
L_PG3_12|_AND_G|B2 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B2  4.135667696e-12
L_PG3_12|_AND_G|B3 _PG3_12|_AND_G|B3 _PG3_12|_AND_G|Q3  1.2e-12
L_PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|Q2  4.135667696e-12
L_PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q1  4.135667696e-12
L_PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1 G3_2  2.067833848e-12
L_DFF_IP1_12|I_1|B _DFF_IP1_12|A1 _DFF_IP1_12|I_1|MID  2e-12
I_DFF_IP1_12|I_1|B 0 _DFF_IP1_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_3|B _DFF_IP1_12|A3 _DFF_IP1_12|I_3|MID  2e-12
I_DFF_IP1_12|I_3|B 0 _DFF_IP1_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP1_12|I_T|B _DFF_IP1_12|T1 _DFF_IP1_12|I_T|MID  2e-12
I_DFF_IP1_12|I_T|B 0 _DFF_IP1_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP1_12|I_6|B _DFF_IP1_12|Q1 _DFF_IP1_12|I_6|MID  2e-12
I_DFF_IP1_12|I_6|B 0 _DFF_IP1_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP1_12|1|1 _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|1|P _DFF_IP1_12|1|MID_SERIES 0  2e-13
R_DFF_IP1_12|1|B _DFF_IP1_12|A1 _DFF_IP1_12|1|MID_SHUNT  2.7439617672
L_DFF_IP1_12|1|RB _DFF_IP1_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|23|1 _DFF_IP1_12|A2 _DFF_IP1_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|23|B _DFF_IP1_12|A2 _DFF_IP1_12|23|MID_SHUNT  3.84154647408
L_DFF_IP1_12|23|RB _DFF_IP1_12|23|MID_SHUNT _DFF_IP1_12|A3  2.1704737578552e-12
B_DFF_IP1_12|3|1 _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|3|P _DFF_IP1_12|3|MID_SERIES 0  2e-13
R_DFF_IP1_12|3|B _DFF_IP1_12|A3 _DFF_IP1_12|3|MID_SHUNT  2.7439617672
L_DFF_IP1_12|3|RB _DFF_IP1_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|4|1 _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|4|P _DFF_IP1_12|4|MID_SERIES 0  2e-13
R_DFF_IP1_12|4|B _DFF_IP1_12|A4 _DFF_IP1_12|4|MID_SHUNT  2.7439617672
L_DFF_IP1_12|4|RB _DFF_IP1_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|T|1 _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|T|P _DFF_IP1_12|T|MID_SERIES 0  2e-13
R_DFF_IP1_12|T|B _DFF_IP1_12|T1 _DFF_IP1_12|T|MID_SHUNT  2.7439617672
L_DFF_IP1_12|T|RB _DFF_IP1_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP1_12|45|1 _DFF_IP1_12|T2 _DFF_IP1_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP1_12|45|B _DFF_IP1_12|T2 _DFF_IP1_12|45|MID_SHUNT  3.84154647408
L_DFF_IP1_12|45|RB _DFF_IP1_12|45|MID_SHUNT _DFF_IP1_12|A4  2.1704737578552e-12
B_DFF_IP1_12|6|1 _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP1_12|6|P _DFF_IP1_12|6|MID_SERIES 0  2e-13
R_DFF_IP1_12|6|B _DFF_IP1_12|Q1 _DFF_IP1_12|6|MID_SHUNT  2.7439617672
L_DFF_IP1_12|6|RB _DFF_IP1_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP2_12|I_1|B _DFF_IP2_12|A1 _DFF_IP2_12|I_1|MID  2e-12
I_DFF_IP2_12|I_1|B 0 _DFF_IP2_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_3|B _DFF_IP2_12|A3 _DFF_IP2_12|I_3|MID  2e-12
I_DFF_IP2_12|I_3|B 0 _DFF_IP2_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP2_12|I_T|B _DFF_IP2_12|T1 _DFF_IP2_12|I_T|MID  2e-12
I_DFF_IP2_12|I_T|B 0 _DFF_IP2_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP2_12|I_6|B _DFF_IP2_12|Q1 _DFF_IP2_12|I_6|MID  2e-12
I_DFF_IP2_12|I_6|B 0 _DFF_IP2_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP2_12|1|1 _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|1|P _DFF_IP2_12|1|MID_SERIES 0  2e-13
R_DFF_IP2_12|1|B _DFF_IP2_12|A1 _DFF_IP2_12|1|MID_SHUNT  2.7439617672
L_DFF_IP2_12|1|RB _DFF_IP2_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|23|1 _DFF_IP2_12|A2 _DFF_IP2_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|23|B _DFF_IP2_12|A2 _DFF_IP2_12|23|MID_SHUNT  3.84154647408
L_DFF_IP2_12|23|RB _DFF_IP2_12|23|MID_SHUNT _DFF_IP2_12|A3  2.1704737578552e-12
B_DFF_IP2_12|3|1 _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|3|P _DFF_IP2_12|3|MID_SERIES 0  2e-13
R_DFF_IP2_12|3|B _DFF_IP2_12|A3 _DFF_IP2_12|3|MID_SHUNT  2.7439617672
L_DFF_IP2_12|3|RB _DFF_IP2_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|4|1 _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|4|P _DFF_IP2_12|4|MID_SERIES 0  2e-13
R_DFF_IP2_12|4|B _DFF_IP2_12|A4 _DFF_IP2_12|4|MID_SHUNT  2.7439617672
L_DFF_IP2_12|4|RB _DFF_IP2_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|T|1 _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|T|P _DFF_IP2_12|T|MID_SERIES 0  2e-13
R_DFF_IP2_12|T|B _DFF_IP2_12|T1 _DFF_IP2_12|T|MID_SHUNT  2.7439617672
L_DFF_IP2_12|T|RB _DFF_IP2_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP2_12|45|1 _DFF_IP2_12|T2 _DFF_IP2_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP2_12|45|B _DFF_IP2_12|T2 _DFF_IP2_12|45|MID_SHUNT  3.84154647408
L_DFF_IP2_12|45|RB _DFF_IP2_12|45|MID_SHUNT _DFF_IP2_12|A4  2.1704737578552e-12
B_DFF_IP2_12|6|1 _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP2_12|6|P _DFF_IP2_12|6|MID_SERIES 0  2e-13
R_DFF_IP2_12|6|B _DFF_IP2_12|Q1 _DFF_IP2_12|6|MID_SHUNT  2.7439617672
L_DFF_IP2_12|6|RB _DFF_IP2_12|6|MID_SHUNT 0  1.550338398468e-12
L_DFF_IP3_12|I_1|B _DFF_IP3_12|A1 _DFF_IP3_12|I_1|MID  2e-12
I_DFF_IP3_12|I_1|B 0 _DFF_IP3_12|I_1|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_3|B _DFF_IP3_12|A3 _DFF_IP3_12|I_3|MID  2e-12
I_DFF_IP3_12|I_3|B 0 _DFF_IP3_12|I_3|MID  PWL(0 0 5e-12 0.00025)
L_DFF_IP3_12|I_T|B _DFF_IP3_12|T1 _DFF_IP3_12|I_T|MID  2e-12
I_DFF_IP3_12|I_T|B 0 _DFF_IP3_12|I_T|MID  PWL(0 0 5e-12 0.000175)
L_DFF_IP3_12|I_6|B _DFF_IP3_12|Q1 _DFF_IP3_12|I_6|MID  2e-12
I_DFF_IP3_12|I_6|B 0 _DFF_IP3_12|I_6|MID  PWL(0 0 5e-12 0.000175)
B_DFF_IP3_12|1|1 _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|1|P _DFF_IP3_12|1|MID_SERIES 0  2e-13
R_DFF_IP3_12|1|B _DFF_IP3_12|A1 _DFF_IP3_12|1|MID_SHUNT  2.7439617672
L_DFF_IP3_12|1|RB _DFF_IP3_12|1|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|23|1 _DFF_IP3_12|A2 _DFF_IP3_12|A3 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|23|B _DFF_IP3_12|A2 _DFF_IP3_12|23|MID_SHUNT  3.84154647408
L_DFF_IP3_12|23|RB _DFF_IP3_12|23|MID_SHUNT _DFF_IP3_12|A3  2.1704737578552e-12
B_DFF_IP3_12|3|1 _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|3|P _DFF_IP3_12|3|MID_SERIES 0  2e-13
R_DFF_IP3_12|3|B _DFF_IP3_12|A3 _DFF_IP3_12|3|MID_SHUNT  2.7439617672
L_DFF_IP3_12|3|RB _DFF_IP3_12|3|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|4|1 _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|4|P _DFF_IP3_12|4|MID_SERIES 0  2e-13
R_DFF_IP3_12|4|B _DFF_IP3_12|A4 _DFF_IP3_12|4|MID_SHUNT  2.7439617672
L_DFF_IP3_12|4|RB _DFF_IP3_12|4|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|T|1 _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|T|P _DFF_IP3_12|T|MID_SERIES 0  2e-13
R_DFF_IP3_12|T|B _DFF_IP3_12|T1 _DFF_IP3_12|T|MID_SHUNT  2.7439617672
L_DFF_IP3_12|T|RB _DFF_IP3_12|T|MID_SHUNT 0  1.550338398468e-12
B_DFF_IP3_12|45|1 _DFF_IP3_12|T2 _DFF_IP3_12|A4 JJMIT AREA=1.7857142857142858
R_DFF_IP3_12|45|B _DFF_IP3_12|T2 _DFF_IP3_12|45|MID_SHUNT  3.84154647408
L_DFF_IP3_12|45|RB _DFF_IP3_12|45|MID_SHUNT _DFF_IP3_12|A4  2.1704737578552e-12
B_DFF_IP3_12|6|1 _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SERIES JJMIT AREA=2.5
L_DFF_IP3_12|6|P _DFF_IP3_12|6|MID_SERIES 0  2e-13
R_DFF_IP3_12|6|B _DFF_IP3_12|Q1 _DFF_IP3_12|6|MID_SHUNT  2.7439617672
L_DFF_IP3_12|6|RB _DFF_IP3_12|6|MID_SHUNT 0  1.550338398468e-12
L_S0|I_1|B _S0|A1 _S0|I_1|MID  2e-12
I_S0|I_1|B 0 _S0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_3|B _S0|A3 _S0|I_3|MID  2e-12
I_S0|I_3|B 0 _S0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S0|I_T|B _S0|T1 _S0|I_T|MID  2e-12
I_S0|I_T|B 0 _S0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S0|I_6|B _S0|Q1 _S0|I_6|MID  2e-12
I_S0|I_6|B 0 _S0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S0|1|1 _S0|A1 _S0|1|MID_SERIES JJMIT AREA=2.5
L_S0|1|P _S0|1|MID_SERIES 0  2e-13
R_S0|1|B _S0|A1 _S0|1|MID_SHUNT  2.7439617672
L_S0|1|RB _S0|1|MID_SHUNT 0  1.550338398468e-12
B_S0|23|1 _S0|A2 _S0|A3 JJMIT AREA=1.7857142857142858
R_S0|23|B _S0|A2 _S0|23|MID_SHUNT  3.84154647408
L_S0|23|RB _S0|23|MID_SHUNT _S0|A3  2.1704737578552e-12
B_S0|3|1 _S0|A3 _S0|3|MID_SERIES JJMIT AREA=2.5
L_S0|3|P _S0|3|MID_SERIES 0  2e-13
R_S0|3|B _S0|A3 _S0|3|MID_SHUNT  2.7439617672
L_S0|3|RB _S0|3|MID_SHUNT 0  1.550338398468e-12
B_S0|4|1 _S0|A4 _S0|4|MID_SERIES JJMIT AREA=2.5
L_S0|4|P _S0|4|MID_SERIES 0  2e-13
R_S0|4|B _S0|A4 _S0|4|MID_SHUNT  2.7439617672
L_S0|4|RB _S0|4|MID_SHUNT 0  1.550338398468e-12
B_S0|T|1 _S0|T1 _S0|T|MID_SERIES JJMIT AREA=2.5
L_S0|T|P _S0|T|MID_SERIES 0  2e-13
R_S0|T|B _S0|T1 _S0|T|MID_SHUNT  2.7439617672
L_S0|T|RB _S0|T|MID_SHUNT 0  1.550338398468e-12
B_S0|45|1 _S0|T2 _S0|A4 JJMIT AREA=1.7857142857142858
R_S0|45|B _S0|T2 _S0|45|MID_SHUNT  3.84154647408
L_S0|45|RB _S0|45|MID_SHUNT _S0|A4  2.1704737578552e-12
B_S0|6|1 _S0|Q1 _S0|6|MID_SERIES JJMIT AREA=2.5
L_S0|6|P _S0|6|MID_SERIES 0  2e-13
R_S0|6|B _S0|Q1 _S0|6|MID_SHUNT  2.7439617672
L_S0|6|RB _S0|6|MID_SHUNT 0  1.550338398468e-12
BBUF_G0_2|1|1 BUF_G0_2|1 BUF_G0_2|1|MID_SERIES JJMIT AREA=2.5
LBUF_G0_2|1|P BUF_G0_2|1|MID_SERIES 0  2e-13
RBUF_G0_2|1|B BUF_G0_2|1 BUF_G0_2|1|MID_SHUNT  2.7439617672
LBUF_G0_2|1|RB BUF_G0_2|1|MID_SHUNT 0  1.750338398468e-12
LBUF_G0_2|B|B BUF_G0_2|4 BUF_G0_2|B|MID  2e-12
IBUF_G0_2|B|B 0 BUF_G0_2|B|MID  PWL(0 0 5e-12 0.0005)
BBUF_G0_2|2|1 BUF_G0_2|6 BUF_G0_2|2|MID_SERIES JJMIT AREA=2.5
LBUF_G0_2|2|P BUF_G0_2|2|MID_SERIES 0  2e-13
RBUF_G0_2|2|B BUF_G0_2|6 BUF_G0_2|2|MID_SHUNT  2.7439617672
LBUF_G0_2|2|RB BUF_G0_2|2|MID_SHUNT 0  1.750338398468e-12
BBUF_IP1_2|1|1 BUF_IP1_2|1 BUF_IP1_2|1|MID_SERIES JJMIT AREA=2.5
LBUF_IP1_2|1|P BUF_IP1_2|1|MID_SERIES 0  2e-13
RBUF_IP1_2|1|B BUF_IP1_2|1 BUF_IP1_2|1|MID_SHUNT  2.7439617672
LBUF_IP1_2|1|RB BUF_IP1_2|1|MID_SHUNT 0  1.750338398468e-12
LBUF_IP1_2|B|B BUF_IP1_2|4 BUF_IP1_2|B|MID  2e-12
IBUF_IP1_2|B|B 0 BUF_IP1_2|B|MID  PWL(0 0 5e-12 0.0005)
BBUF_IP1_2|2|1 BUF_IP1_2|6 BUF_IP1_2|2|MID_SERIES JJMIT AREA=2.5
LBUF_IP1_2|2|P BUF_IP1_2|2|MID_SERIES 0  2e-13
RBUF_IP1_2|2|B BUF_IP1_2|6 BUF_IP1_2|2|MID_SHUNT  2.7439617672
LBUF_IP1_2|2|RB BUF_IP1_2|2|MID_SHUNT 0  1.750338398468e-12
L_S1|I_A1|B _S1|A1 _S1|I_A1|MID  2e-12
I_S1|I_A1|B 0 _S1|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_A3|B _S1|A3 _S1|I_A3|MID  2e-12
I_S1|I_A3|B 0 _S1|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B1|B _S1|B1 _S1|I_B1|MID  2e-12
I_S1|I_B1|B 0 _S1|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_B3|B _S1|B3 _S1|I_B3|MID  2e-12
I_S1|I_B3|B 0 _S1|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S1|I_Q1|B _S1|Q1 _S1|I_Q1|MID  2e-12
I_S1|I_Q1|B 0 _S1|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S1|A1|1 _S1|A1 _S1|A1|MID_SERIES JJMIT AREA=2.5
L_S1|A1|P _S1|A1|MID_SERIES 0  5e-13
R_S1|A1|B _S1|A1 _S1|A1|MID_SHUNT  2.7439617672
L_S1|A1|RB _S1|A1|MID_SHUNT 0  2.050338398468e-12
B_S1|A2|1 _S1|A2 _S1|A2|MID_SERIES JJMIT AREA=2.5
L_S1|A2|P _S1|A2|MID_SERIES 0  5e-13
R_S1|A2|B _S1|A2 _S1|A2|MID_SHUNT  2.7439617672
L_S1|A2|RB _S1|A2|MID_SHUNT 0  2.050338398468e-12
B_S1|A3|1 _S1|A2 _S1|A3|MID_SERIES JJMIT AREA=2.5
L_S1|A3|P _S1|A3|MID_SERIES _S1|A3  1.2e-12
R_S1|A3|B _S1|A2 _S1|A3|MID_SHUNT  2.7439617672
L_S1|A3|RB _S1|A3|MID_SHUNT _S1|A3  2.050338398468e-12
B_S1|B1|1 _S1|B1 _S1|B1|MID_SERIES JJMIT AREA=2.5
L_S1|B1|P _S1|B1|MID_SERIES 0  5e-13
R_S1|B1|B _S1|B1 _S1|B1|MID_SHUNT  2.7439617672
L_S1|B1|RB _S1|B1|MID_SHUNT 0  2.050338398468e-12
B_S1|B2|1 _S1|B2 _S1|B2|MID_SERIES JJMIT AREA=2.5
L_S1|B2|P _S1|B2|MID_SERIES 0  5e-13
R_S1|B2|B _S1|B2 _S1|B2|MID_SHUNT  2.7439617672
L_S1|B2|RB _S1|B2|MID_SHUNT 0  2.050338398468e-12
B_S1|B3|1 _S1|B2 _S1|B3|MID_SERIES JJMIT AREA=2.5
L_S1|B3|P _S1|B3|MID_SERIES _S1|B3  1.2e-12
R_S1|B3|B _S1|B2 _S1|B3|MID_SHUNT  2.7439617672
L_S1|B3|RB _S1|B3|MID_SHUNT _S1|B3  2.050338398468e-12
B_S1|T1|1 _S1|T1 _S1|T1|MID_SERIES JJMIT AREA=2.5
L_S1|T1|P _S1|T1|MID_SERIES 0  5e-13
R_S1|T1|B _S1|T1 _S1|T1|MID_SHUNT  2.7439617672
L_S1|T1|RB _S1|T1|MID_SHUNT 0  2.050338398468e-12
B_S1|T2|1 _S1|T2 _S1|ABTQ JJMIT AREA=2.0
R_S1|T2|B _S1|T2 _S1|T2|MID_SHUNT  3.429952209
L_S1|T2|RB _S1|T2|MID_SHUNT _S1|ABTQ  2.437922998085e-12
B_S1|AB|1 _S1|AB _S1|AB|MID_SERIES JJMIT AREA=1.6
L_S1|AB|P _S1|AB|MID_SERIES _S1|ABTQ  1.2e-12
R_S1|AB|B _S1|AB _S1|AB|MID_SHUNT  4.2874402612499996
L_S1|AB|RB _S1|AB|MID_SHUNT _S1|ABTQ  2.92240374760625e-12
B_S1|ABTQ|1 _S1|ABTQ _S1|ABTQ|MID_SERIES JJMIT AREA=2.0
L_S1|ABTQ|P _S1|ABTQ|MID_SERIES 0  5e-13
R_S1|ABTQ|B _S1|ABTQ _S1|ABTQ|MID_SHUNT  3.429952209
L_S1|ABTQ|RB _S1|ABTQ|MID_SHUNT 0  2.437922998085e-12
B_S1|Q1|1 _S1|Q1 _S1|Q1|MID_SERIES JJMIT AREA=2.5
L_S1|Q1|P _S1|Q1|MID_SERIES 0  5e-13
R_S1|Q1|B _S1|Q1 _S1|Q1|MID_SHUNT  2.7439617672
L_S1|Q1|RB _S1|Q1|MID_SHUNT 0  2.050338398468e-12
BBUF_G1_2|1|1 BUF_G1_2|1 BUF_G1_2|1|MID_SERIES JJMIT AREA=2.5
LBUF_G1_2|1|P BUF_G1_2|1|MID_SERIES 0  2e-13
RBUF_G1_2|1|B BUF_G1_2|1 BUF_G1_2|1|MID_SHUNT  2.7439617672
LBUF_G1_2|1|RB BUF_G1_2|1|MID_SHUNT 0  1.750338398468e-12
LBUF_G1_2|B|B BUF_G1_2|4 BUF_G1_2|B|MID  2e-12
IBUF_G1_2|B|B 0 BUF_G1_2|B|MID  PWL(0 0 5e-12 0.0005)
BBUF_G1_2|2|1 BUF_G1_2|6 BUF_G1_2|2|MID_SERIES JJMIT AREA=2.5
LBUF_G1_2|2|P BUF_G1_2|2|MID_SERIES 0  2e-13
RBUF_G1_2|2|B BUF_G1_2|6 BUF_G1_2|2|MID_SHUNT  2.7439617672
LBUF_G1_2|2|RB BUF_G1_2|2|MID_SHUNT 0  1.750338398468e-12
BBUF_IP2_2|1|1 BUF_IP2_2|1 BUF_IP2_2|1|MID_SERIES JJMIT AREA=2.5
LBUF_IP2_2|1|P BUF_IP2_2|1|MID_SERIES 0  2e-13
RBUF_IP2_2|1|B BUF_IP2_2|1 BUF_IP2_2|1|MID_SHUNT  2.7439617672
LBUF_IP2_2|1|RB BUF_IP2_2|1|MID_SHUNT 0  1.750338398468e-12
LBUF_IP2_2|B|B BUF_IP2_2|4 BUF_IP2_2|B|MID  2e-12
IBUF_IP2_2|B|B 0 BUF_IP2_2|B|MID  PWL(0 0 5e-12 0.0005)
BBUF_IP2_2|2|1 BUF_IP2_2|6 BUF_IP2_2|2|MID_SERIES JJMIT AREA=2.5
LBUF_IP2_2|2|P BUF_IP2_2|2|MID_SERIES 0  2e-13
RBUF_IP2_2|2|B BUF_IP2_2|6 BUF_IP2_2|2|MID_SHUNT  2.7439617672
LBUF_IP2_2|2|RB BUF_IP2_2|2|MID_SHUNT 0  1.750338398468e-12
L_S2|I_A1|B _S2|A1 _S2|I_A1|MID  2e-12
I_S2|I_A1|B 0 _S2|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_A3|B _S2|A3 _S2|I_A3|MID  2e-12
I_S2|I_A3|B 0 _S2|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B1|B _S2|B1 _S2|I_B1|MID  2e-12
I_S2|I_B1|B 0 _S2|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_B3|B _S2|B3 _S2|I_B3|MID  2e-12
I_S2|I_B3|B 0 _S2|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S2|I_Q1|B _S2|Q1 _S2|I_Q1|MID  2e-12
I_S2|I_Q1|B 0 _S2|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S2|A1|1 _S2|A1 _S2|A1|MID_SERIES JJMIT AREA=2.5
L_S2|A1|P _S2|A1|MID_SERIES 0  5e-13
R_S2|A1|B _S2|A1 _S2|A1|MID_SHUNT  2.7439617672
L_S2|A1|RB _S2|A1|MID_SHUNT 0  2.050338398468e-12
B_S2|A2|1 _S2|A2 _S2|A2|MID_SERIES JJMIT AREA=2.5
L_S2|A2|P _S2|A2|MID_SERIES 0  5e-13
R_S2|A2|B _S2|A2 _S2|A2|MID_SHUNT  2.7439617672
L_S2|A2|RB _S2|A2|MID_SHUNT 0  2.050338398468e-12
B_S2|A3|1 _S2|A2 _S2|A3|MID_SERIES JJMIT AREA=2.5
L_S2|A3|P _S2|A3|MID_SERIES _S2|A3  1.2e-12
R_S2|A3|B _S2|A2 _S2|A3|MID_SHUNT  2.7439617672
L_S2|A3|RB _S2|A3|MID_SHUNT _S2|A3  2.050338398468e-12
B_S2|B1|1 _S2|B1 _S2|B1|MID_SERIES JJMIT AREA=2.5
L_S2|B1|P _S2|B1|MID_SERIES 0  5e-13
R_S2|B1|B _S2|B1 _S2|B1|MID_SHUNT  2.7439617672
L_S2|B1|RB _S2|B1|MID_SHUNT 0  2.050338398468e-12
B_S2|B2|1 _S2|B2 _S2|B2|MID_SERIES JJMIT AREA=2.5
L_S2|B2|P _S2|B2|MID_SERIES 0  5e-13
R_S2|B2|B _S2|B2 _S2|B2|MID_SHUNT  2.7439617672
L_S2|B2|RB _S2|B2|MID_SHUNT 0  2.050338398468e-12
B_S2|B3|1 _S2|B2 _S2|B3|MID_SERIES JJMIT AREA=2.5
L_S2|B3|P _S2|B3|MID_SERIES _S2|B3  1.2e-12
R_S2|B3|B _S2|B2 _S2|B3|MID_SHUNT  2.7439617672
L_S2|B3|RB _S2|B3|MID_SHUNT _S2|B3  2.050338398468e-12
B_S2|T1|1 _S2|T1 _S2|T1|MID_SERIES JJMIT AREA=2.5
L_S2|T1|P _S2|T1|MID_SERIES 0  5e-13
R_S2|T1|B _S2|T1 _S2|T1|MID_SHUNT  2.7439617672
L_S2|T1|RB _S2|T1|MID_SHUNT 0  2.050338398468e-12
B_S2|T2|1 _S2|T2 _S2|ABTQ JJMIT AREA=2.0
R_S2|T2|B _S2|T2 _S2|T2|MID_SHUNT  3.429952209
L_S2|T2|RB _S2|T2|MID_SHUNT _S2|ABTQ  2.437922998085e-12
B_S2|AB|1 _S2|AB _S2|AB|MID_SERIES JJMIT AREA=1.6
L_S2|AB|P _S2|AB|MID_SERIES _S2|ABTQ  1.2e-12
R_S2|AB|B _S2|AB _S2|AB|MID_SHUNT  4.2874402612499996
L_S2|AB|RB _S2|AB|MID_SHUNT _S2|ABTQ  2.92240374760625e-12
B_S2|ABTQ|1 _S2|ABTQ _S2|ABTQ|MID_SERIES JJMIT AREA=2.0
L_S2|ABTQ|P _S2|ABTQ|MID_SERIES 0  5e-13
R_S2|ABTQ|B _S2|ABTQ _S2|ABTQ|MID_SHUNT  3.429952209
L_S2|ABTQ|RB _S2|ABTQ|MID_SHUNT 0  2.437922998085e-12
B_S2|Q1|1 _S2|Q1 _S2|Q1|MID_SERIES JJMIT AREA=2.5
L_S2|Q1|P _S2|Q1|MID_SERIES 0  5e-13
R_S2|Q1|B _S2|Q1 _S2|Q1|MID_SHUNT  2.7439617672
L_S2|Q1|RB _S2|Q1|MID_SHUNT 0  2.050338398468e-12
BBUF_G2_2|1|1 BUF_G2_2|1 BUF_G2_2|1|MID_SERIES JJMIT AREA=2.5
LBUF_G2_2|1|P BUF_G2_2|1|MID_SERIES 0  2e-13
RBUF_G2_2|1|B BUF_G2_2|1 BUF_G2_2|1|MID_SHUNT  2.7439617672
LBUF_G2_2|1|RB BUF_G2_2|1|MID_SHUNT 0  1.750338398468e-12
LBUF_G2_2|B|B BUF_G2_2|4 BUF_G2_2|B|MID  2e-12
IBUF_G2_2|B|B 0 BUF_G2_2|B|MID  PWL(0 0 5e-12 0.0005)
BBUF_G2_2|2|1 BUF_G2_2|6 BUF_G2_2|2|MID_SERIES JJMIT AREA=2.5
LBUF_G2_2|2|P BUF_G2_2|2|MID_SERIES 0  2e-13
RBUF_G2_2|2|B BUF_G2_2|6 BUF_G2_2|2|MID_SHUNT  2.7439617672
LBUF_G2_2|2|RB BUF_G2_2|2|MID_SHUNT 0  1.750338398468e-12
L_S3|I_A1|B _S3|A1 _S3|I_A1|MID  2e-12
I_S3|I_A1|B 0 _S3|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_A3|B _S3|A3 _S3|I_A3|MID  2e-12
I_S3|I_A3|B 0 _S3|I_A3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B1|B _S3|B1 _S3|I_B1|MID  2e-12
I_S3|I_B1|B 0 _S3|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_B3|B _S3|B3 _S3|I_B3|MID  2e-12
I_S3|I_B3|B 0 _S3|I_B3|MID  PWL(0 0 5e-12 0.000175)
L_S3|I_Q1|B _S3|Q1 _S3|I_Q1|MID  2e-12
I_S3|I_Q1|B 0 _S3|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_S3|A1|1 _S3|A1 _S3|A1|MID_SERIES JJMIT AREA=2.5
L_S3|A1|P _S3|A1|MID_SERIES 0  5e-13
R_S3|A1|B _S3|A1 _S3|A1|MID_SHUNT  2.7439617672
L_S3|A1|RB _S3|A1|MID_SHUNT 0  2.050338398468e-12
B_S3|A2|1 _S3|A2 _S3|A2|MID_SERIES JJMIT AREA=2.5
L_S3|A2|P _S3|A2|MID_SERIES 0  5e-13
R_S3|A2|B _S3|A2 _S3|A2|MID_SHUNT  2.7439617672
L_S3|A2|RB _S3|A2|MID_SHUNT 0  2.050338398468e-12
B_S3|A3|1 _S3|A2 _S3|A3|MID_SERIES JJMIT AREA=2.5
L_S3|A3|P _S3|A3|MID_SERIES _S3|A3  1.2e-12
R_S3|A3|B _S3|A2 _S3|A3|MID_SHUNT  2.7439617672
L_S3|A3|RB _S3|A3|MID_SHUNT _S3|A3  2.050338398468e-12
B_S3|B1|1 _S3|B1 _S3|B1|MID_SERIES JJMIT AREA=2.5
L_S3|B1|P _S3|B1|MID_SERIES 0  5e-13
R_S3|B1|B _S3|B1 _S3|B1|MID_SHUNT  2.7439617672
L_S3|B1|RB _S3|B1|MID_SHUNT 0  2.050338398468e-12
B_S3|B2|1 _S3|B2 _S3|B2|MID_SERIES JJMIT AREA=2.5
L_S3|B2|P _S3|B2|MID_SERIES 0  5e-13
R_S3|B2|B _S3|B2 _S3|B2|MID_SHUNT  2.7439617672
L_S3|B2|RB _S3|B2|MID_SHUNT 0  2.050338398468e-12
B_S3|B3|1 _S3|B2 _S3|B3|MID_SERIES JJMIT AREA=2.5
L_S3|B3|P _S3|B3|MID_SERIES _S3|B3  1.2e-12
R_S3|B3|B _S3|B2 _S3|B3|MID_SHUNT  2.7439617672
L_S3|B3|RB _S3|B3|MID_SHUNT _S3|B3  2.050338398468e-12
B_S3|T1|1 _S3|T1 _S3|T1|MID_SERIES JJMIT AREA=2.5
L_S3|T1|P _S3|T1|MID_SERIES 0  5e-13
R_S3|T1|B _S3|T1 _S3|T1|MID_SHUNT  2.7439617672
L_S3|T1|RB _S3|T1|MID_SHUNT 0  2.050338398468e-12
B_S3|T2|1 _S3|T2 _S3|ABTQ JJMIT AREA=2.0
R_S3|T2|B _S3|T2 _S3|T2|MID_SHUNT  3.429952209
L_S3|T2|RB _S3|T2|MID_SHUNT _S3|ABTQ  2.437922998085e-12
B_S3|AB|1 _S3|AB _S3|AB|MID_SERIES JJMIT AREA=1.8
L_S3|AB|P _S3|AB|MID_SERIES _S3|ABTQ  1.2e-12
R_S3|AB|B _S3|AB _S3|AB|MID_SHUNT  3.81105801
L_S3|AB|RB _S3|AB|MID_SHUNT _S3|ABTQ  2.65324777565e-12
B_S3|ABTQ|1 _S3|ABTQ _S3|ABTQ|MID_SERIES JJMIT AREA=2.25
L_S3|ABTQ|P _S3|ABTQ|MID_SERIES 0  5e-13
R_S3|ABTQ|B _S3|ABTQ _S3|ABTQ|MID_SHUNT  3.048846408
L_S3|ABTQ|RB _S3|ABTQ|MID_SHUNT 0  2.2225982205200003e-12
B_S3|Q1|1 _S3|Q1 _S3|Q1|MID_SERIES JJMIT AREA=2.5
L_S3|Q1|P _S3|Q1|MID_SERIES 0  5e-13
R_S3|Q1|B _S3|Q1 _S3|Q1|MID_SHUNT  2.7439617672
L_S3|Q1|RB _S3|Q1|MID_SHUNT 0  2.050338398468e-12
L_S4|I_1|B _S4|A1 _S4|I_1|MID  2e-12
I_S4|I_1|B 0 _S4|I_1|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_3|B _S4|A3 _S4|I_3|MID  2e-12
I_S4|I_3|B 0 _S4|I_3|MID  PWL(0 0 5e-12 0.00025)
L_S4|I_T|B _S4|T1 _S4|I_T|MID  2e-12
I_S4|I_T|B 0 _S4|I_T|MID  PWL(0 0 5e-12 0.000175)
L_S4|I_6|B _S4|Q1 _S4|I_6|MID  2e-12
I_S4|I_6|B 0 _S4|I_6|MID  PWL(0 0 5e-12 0.000175)
B_S4|1|1 _S4|A1 _S4|1|MID_SERIES JJMIT AREA=2.5
L_S4|1|P _S4|1|MID_SERIES 0  2e-13
R_S4|1|B _S4|A1 _S4|1|MID_SHUNT  2.7439617672
L_S4|1|RB _S4|1|MID_SHUNT 0  1.550338398468e-12
B_S4|23|1 _S4|A2 _S4|A3 JJMIT AREA=1.7857142857142858
R_S4|23|B _S4|A2 _S4|23|MID_SHUNT  3.84154647408
L_S4|23|RB _S4|23|MID_SHUNT _S4|A3  2.1704737578552e-12
B_S4|3|1 _S4|A3 _S4|3|MID_SERIES JJMIT AREA=2.5
L_S4|3|P _S4|3|MID_SERIES 0  2e-13
R_S4|3|B _S4|A3 _S4|3|MID_SHUNT  2.7439617672
L_S4|3|RB _S4|3|MID_SHUNT 0  1.550338398468e-12
B_S4|4|1 _S4|A4 _S4|4|MID_SERIES JJMIT AREA=2.5
L_S4|4|P _S4|4|MID_SERIES 0  2e-13
R_S4|4|B _S4|A4 _S4|4|MID_SHUNT  2.7439617672
L_S4|4|RB _S4|4|MID_SHUNT 0  1.550338398468e-12
B_S4|T|1 _S4|T1 _S4|T|MID_SERIES JJMIT AREA=2.5
L_S4|T|P _S4|T|MID_SERIES 0  2e-13
R_S4|T|B _S4|T1 _S4|T|MID_SHUNT  2.7439617672
L_S4|T|RB _S4|T|MID_SHUNT 0  1.550338398468e-12
B_S4|45|1 _S4|T2 _S4|A4 JJMIT AREA=1.7857142857142858
R_S4|45|B _S4|T2 _S4|45|MID_SHUNT  3.84154647408
L_S4|45|RB _S4|45|MID_SHUNT _S4|A4  2.1704737578552e-12
B_S4|6|1 _S4|Q1 _S4|6|MID_SERIES JJMIT AREA=2.5
L_S4|6|P _S4|6|MID_SERIES 0  2e-13
R_S4|6|B _S4|Q1 _S4|6|MID_SHUNT  2.7439617672
L_S4|6|RB _S4|6|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_A|I_D1|B I0|_SPL_A|D1 I0|_SPL_A|I_D1|MID  2e-12
II0|_SPL_A|I_D1|B 0 I0|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_D2|B I0|_SPL_A|D2 I0|_SPL_A|I_D2|MID  2e-12
II0|_SPL_A|I_D2|B 0 I0|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_A|I_Q1|B I0|_SPL_A|QA1 I0|_SPL_A|I_Q1|MID  2e-12
II0|_SPL_A|I_Q1|B 0 I0|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_A|I_Q2|B I0|_SPL_A|QB1 I0|_SPL_A|I_Q2|MID  2e-12
II0|_SPL_A|I_Q2|B 0 I0|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_A|1|1 I0|_SPL_A|D1 I0|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|1|P I0|_SPL_A|1|MID_SERIES 0  2e-13
RI0|_SPL_A|1|B I0|_SPL_A|D1 I0|_SPL_A|1|MID_SHUNT  2.7439617672
LI0|_SPL_A|1|RB I0|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|2|1 I0|_SPL_A|D2 I0|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|2|P I0|_SPL_A|2|MID_SERIES 0  2e-13
RI0|_SPL_A|2|B I0|_SPL_A|D2 I0|_SPL_A|2|MID_SHUNT  2.7439617672
LI0|_SPL_A|2|RB I0|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|A|1 I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|A|P I0|_SPL_A|A|MID_SERIES 0  2e-13
RI0|_SPL_A|A|B I0|_SPL_A|QA1 I0|_SPL_A|A|MID_SHUNT  2.7439617672
LI0|_SPL_A|A|RB I0|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_A|B|1 I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_A|B|P I0|_SPL_A|B|MID_SERIES 0  2e-13
RI0|_SPL_A|B|B I0|_SPL_A|QB1 I0|_SPL_A|B|MID_SHUNT  2.7439617672
LI0|_SPL_A|B|RB I0|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI0|_SPL_B|I_D1|B I0|_SPL_B|D1 I0|_SPL_B|I_D1|MID  2e-12
II0|_SPL_B|I_D1|B 0 I0|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_D2|B I0|_SPL_B|D2 I0|_SPL_B|I_D2|MID  2e-12
II0|_SPL_B|I_D2|B 0 I0|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI0|_SPL_B|I_Q1|B I0|_SPL_B|QA1 I0|_SPL_B|I_Q1|MID  2e-12
II0|_SPL_B|I_Q1|B 0 I0|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI0|_SPL_B|I_Q2|B I0|_SPL_B|QB1 I0|_SPL_B|I_Q2|MID  2e-12
II0|_SPL_B|I_Q2|B 0 I0|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI0|_SPL_B|1|1 I0|_SPL_B|D1 I0|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|1|P I0|_SPL_B|1|MID_SERIES 0  2e-13
RI0|_SPL_B|1|B I0|_SPL_B|D1 I0|_SPL_B|1|MID_SHUNT  2.7439617672
LI0|_SPL_B|1|RB I0|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|2|1 I0|_SPL_B|D2 I0|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|2|P I0|_SPL_B|2|MID_SERIES 0  2e-13
RI0|_SPL_B|2|B I0|_SPL_B|D2 I0|_SPL_B|2|MID_SHUNT  2.7439617672
LI0|_SPL_B|2|RB I0|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|A|1 I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|A|P I0|_SPL_B|A|MID_SERIES 0  2e-13
RI0|_SPL_B|A|B I0|_SPL_B|QA1 I0|_SPL_B|A|MID_SHUNT  2.7439617672
LI0|_SPL_B|A|RB I0|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI0|_SPL_B|B|1 I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI0|_SPL_B|B|P I0|_SPL_B|B|MID_SERIES 0  2e-13
RI0|_SPL_B|B|B I0|_SPL_B|QB1 I0|_SPL_B|B|MID_SHUNT  2.7439617672
LI0|_SPL_B|B|RB I0|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_A|I_1|B I0|_DFF_A|A1 I0|_DFF_A|I_1|MID  2e-12
II0|_DFF_A|I_1|B 0 I0|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_3|B I0|_DFF_A|A3 I0|_DFF_A|I_3|MID  2e-12
II0|_DFF_A|I_3|B 0 I0|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_A|I_T|B I0|_DFF_A|T1 I0|_DFF_A|I_T|MID  2e-12
II0|_DFF_A|I_T|B 0 I0|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_A|I_6|B I0|_DFF_A|Q1 I0|_DFF_A|I_6|MID  2e-12
II0|_DFF_A|I_6|B 0 I0|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_A|1|1 I0|_DFF_A|A1 I0|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|1|P I0|_DFF_A|1|MID_SERIES 0  2e-13
RI0|_DFF_A|1|B I0|_DFF_A|A1 I0|_DFF_A|1|MID_SHUNT  2.7439617672
LI0|_DFF_A|1|RB I0|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|23|1 I0|_DFF_A|A2 I0|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|23|B I0|_DFF_A|A2 I0|_DFF_A|23|MID_SHUNT  3.84154647408
LI0|_DFF_A|23|RB I0|_DFF_A|23|MID_SHUNT I0|_DFF_A|A3  2.1704737578552e-12
BI0|_DFF_A|3|1 I0|_DFF_A|A3 I0|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|3|P I0|_DFF_A|3|MID_SERIES 0  2e-13
RI0|_DFF_A|3|B I0|_DFF_A|A3 I0|_DFF_A|3|MID_SHUNT  2.7439617672
LI0|_DFF_A|3|RB I0|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|4|1 I0|_DFF_A|A4 I0|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|4|P I0|_DFF_A|4|MID_SERIES 0  2e-13
RI0|_DFF_A|4|B I0|_DFF_A|A4 I0|_DFF_A|4|MID_SHUNT  2.7439617672
LI0|_DFF_A|4|RB I0|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|T|1 I0|_DFF_A|T1 I0|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|T|P I0|_DFF_A|T|MID_SERIES 0  2e-13
RI0|_DFF_A|T|B I0|_DFF_A|T1 I0|_DFF_A|T|MID_SHUNT  2.7439617672
LI0|_DFF_A|T|RB I0|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_A|45|1 I0|_DFF_A|T2 I0|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_A|45|B I0|_DFF_A|T2 I0|_DFF_A|45|MID_SHUNT  3.84154647408
LI0|_DFF_A|45|RB I0|_DFF_A|45|MID_SHUNT I0|_DFF_A|A4  2.1704737578552e-12
BI0|_DFF_A|6|1 I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_A|6|P I0|_DFF_A|6|MID_SERIES 0  2e-13
RI0|_DFF_A|6|B I0|_DFF_A|Q1 I0|_DFF_A|6|MID_SHUNT  2.7439617672
LI0|_DFF_A|6|RB I0|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI0|_DFF_B|I_1|B I0|_DFF_B|A1 I0|_DFF_B|I_1|MID  2e-12
II0|_DFF_B|I_1|B 0 I0|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_3|B I0|_DFF_B|A3 I0|_DFF_B|I_3|MID  2e-12
II0|_DFF_B|I_3|B 0 I0|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI0|_DFF_B|I_T|B I0|_DFF_B|T1 I0|_DFF_B|I_T|MID  2e-12
II0|_DFF_B|I_T|B 0 I0|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI0|_DFF_B|I_6|B I0|_DFF_B|Q1 I0|_DFF_B|I_6|MID  2e-12
II0|_DFF_B|I_6|B 0 I0|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI0|_DFF_B|1|1 I0|_DFF_B|A1 I0|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|1|P I0|_DFF_B|1|MID_SERIES 0  2e-13
RI0|_DFF_B|1|B I0|_DFF_B|A1 I0|_DFF_B|1|MID_SHUNT  2.7439617672
LI0|_DFF_B|1|RB I0|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|23|1 I0|_DFF_B|A2 I0|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|23|B I0|_DFF_B|A2 I0|_DFF_B|23|MID_SHUNT  3.84154647408
LI0|_DFF_B|23|RB I0|_DFF_B|23|MID_SHUNT I0|_DFF_B|A3  2.1704737578552e-12
BI0|_DFF_B|3|1 I0|_DFF_B|A3 I0|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|3|P I0|_DFF_B|3|MID_SERIES 0  2e-13
RI0|_DFF_B|3|B I0|_DFF_B|A3 I0|_DFF_B|3|MID_SHUNT  2.7439617672
LI0|_DFF_B|3|RB I0|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|4|1 I0|_DFF_B|A4 I0|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|4|P I0|_DFF_B|4|MID_SERIES 0  2e-13
RI0|_DFF_B|4|B I0|_DFF_B|A4 I0|_DFF_B|4|MID_SHUNT  2.7439617672
LI0|_DFF_B|4|RB I0|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|T|1 I0|_DFF_B|T1 I0|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|T|P I0|_DFF_B|T|MID_SERIES 0  2e-13
RI0|_DFF_B|T|B I0|_DFF_B|T1 I0|_DFF_B|T|MID_SHUNT  2.7439617672
LI0|_DFF_B|T|RB I0|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI0|_DFF_B|45|1 I0|_DFF_B|T2 I0|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI0|_DFF_B|45|B I0|_DFF_B|T2 I0|_DFF_B|45|MID_SHUNT  3.84154647408
LI0|_DFF_B|45|RB I0|_DFF_B|45|MID_SHUNT I0|_DFF_B|A4  2.1704737578552e-12
BI0|_DFF_B|6|1 I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI0|_DFF_B|6|P I0|_DFF_B|6|MID_SERIES 0  2e-13
RI0|_DFF_B|6|B I0|_DFF_B|Q1 I0|_DFF_B|6|MID_SHUNT  2.7439617672
LI0|_DFF_B|6|RB I0|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI0|_XOR|I_A1|B I0|_XOR|A1 I0|_XOR|I_A1|MID  2e-12
II0|_XOR|I_A1|B 0 I0|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_A3|B I0|_XOR|A3 I0|_XOR|I_A3|MID  2e-12
II0|_XOR|I_A3|B 0 I0|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B1|B I0|_XOR|B1 I0|_XOR|I_B1|MID  2e-12
II0|_XOR|I_B1|B 0 I0|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_B3|B I0|_XOR|B3 I0|_XOR|I_B3|MID  2e-12
II0|_XOR|I_B3|B 0 I0|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI0|_XOR|I_Q1|B I0|_XOR|Q1 I0|_XOR|I_Q1|MID  2e-12
II0|_XOR|I_Q1|B 0 I0|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_XOR|A1|1 I0|_XOR|A1 I0|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A1|P I0|_XOR|A1|MID_SERIES 0  5e-13
RI0|_XOR|A1|B I0|_XOR|A1 I0|_XOR|A1|MID_SHUNT  2.7439617672
LI0|_XOR|A1|RB I0|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A2|1 I0|_XOR|A2 I0|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A2|P I0|_XOR|A2|MID_SERIES 0  5e-13
RI0|_XOR|A2|B I0|_XOR|A2 I0|_XOR|A2|MID_SHUNT  2.7439617672
LI0|_XOR|A2|RB I0|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|A3|1 I0|_XOR|A2 I0|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|A3|P I0|_XOR|A3|MID_SERIES I0|_XOR|A3  1.2e-12
RI0|_XOR|A3|B I0|_XOR|A2 I0|_XOR|A3|MID_SHUNT  2.7439617672
LI0|_XOR|A3|RB I0|_XOR|A3|MID_SHUNT I0|_XOR|A3  2.050338398468e-12
BI0|_XOR|B1|1 I0|_XOR|B1 I0|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B1|P I0|_XOR|B1|MID_SERIES 0  5e-13
RI0|_XOR|B1|B I0|_XOR|B1 I0|_XOR|B1|MID_SHUNT  2.7439617672
LI0|_XOR|B1|RB I0|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B2|1 I0|_XOR|B2 I0|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B2|P I0|_XOR|B2|MID_SERIES 0  5e-13
RI0|_XOR|B2|B I0|_XOR|B2 I0|_XOR|B2|MID_SHUNT  2.7439617672
LI0|_XOR|B2|RB I0|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|B3|1 I0|_XOR|B2 I0|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|B3|P I0|_XOR|B3|MID_SERIES I0|_XOR|B3  1.2e-12
RI0|_XOR|B3|B I0|_XOR|B2 I0|_XOR|B3|MID_SHUNT  2.7439617672
LI0|_XOR|B3|RB I0|_XOR|B3|MID_SHUNT I0|_XOR|B3  2.050338398468e-12
BI0|_XOR|T1|1 I0|_XOR|T1 I0|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|T1|P I0|_XOR|T1|MID_SERIES 0  5e-13
RI0|_XOR|T1|B I0|_XOR|T1 I0|_XOR|T1|MID_SHUNT  2.7439617672
LI0|_XOR|T1|RB I0|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|T2|1 I0|_XOR|T2 I0|_XOR|ABTQ JJMIT AREA=2.0
RI0|_XOR|T2|B I0|_XOR|T2 I0|_XOR|T2|MID_SHUNT  3.429952209
LI0|_XOR|T2|RB I0|_XOR|T2|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|AB|1 I0|_XOR|AB I0|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI0|_XOR|AB|P I0|_XOR|AB|MID_SERIES I0|_XOR|ABTQ  1.2e-12
RI0|_XOR|AB|B I0|_XOR|AB I0|_XOR|AB|MID_SHUNT  3.429952209
LI0|_XOR|AB|RB I0|_XOR|AB|MID_SHUNT I0|_XOR|ABTQ  2.437922998085e-12
BI0|_XOR|ABTQ|1 I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|ABTQ|P I0|_XOR|ABTQ|MID_SERIES 0  5e-13
RI0|_XOR|ABTQ|B I0|_XOR|ABTQ I0|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI0|_XOR|ABTQ|RB I0|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI0|_XOR|Q1|1 I0|_XOR|Q1 I0|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_XOR|Q1|P I0|_XOR|Q1|MID_SERIES 0  5e-13
RI0|_XOR|Q1|B I0|_XOR|Q1 I0|_XOR|Q1|MID_SHUNT  2.7439617672
LI0|_XOR|Q1|RB I0|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI0|_AND|I_A1|B I0|_AND|A1 I0|_AND|I_A1|MID  2e-12
II0|_AND|I_A1|B 0 I0|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_B1|B I0|_AND|B1 I0|_AND|I_B1|MID  2e-12
II0|_AND|I_B1|B 0 I0|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q3|B I0|_AND|Q3 I0|_AND|I_Q3|MID  2e-12
II0|_AND|I_Q3|B 0 I0|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI0|_AND|I_Q2|B I0|_AND|Q2 I0|_AND|I_Q2|MID  2e-12
II0|_AND|I_Q2|B 0 I0|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI0|_AND|I_Q1|B I0|_AND|Q1 I0|_AND|I_Q1|MID  2e-12
II0|_AND|I_Q1|B 0 I0|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI0|_AND|A1|1 I0|_AND|A1 I0|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A1|P I0|_AND|A1|MID_SERIES 0  2e-13
RI0|_AND|A1|B I0|_AND|A1 I0|_AND|A1|MID_SHUNT  2.7439617672
LI0|_AND|A1|RB I0|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A2|1 I0|_AND|A2 I0|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|A2|P I0|_AND|A2|MID_SERIES 0  2e-13
RI0|_AND|A2|B I0|_AND|A2 I0|_AND|A2|MID_SHUNT  2.7439617672
LI0|_AND|A2|RB I0|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|A12|1 I0|_AND|A2 I0|_AND|A3 JJMIT AREA=1.7857142857142858
RI0|_AND|A12|B I0|_AND|A2 I0|_AND|A12|MID_SHUNT  3.84154647408
LI0|_AND|A12|RB I0|_AND|A12|MID_SHUNT I0|_AND|A3  2.1704737578552e-12
BI0|_AND|B1|1 I0|_AND|B1 I0|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B1|P I0|_AND|B1|MID_SERIES 0  2e-13
RI0|_AND|B1|B I0|_AND|B1 I0|_AND|B1|MID_SHUNT  2.7439617672
LI0|_AND|B1|RB I0|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B2|1 I0|_AND|B2 I0|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|B2|P I0|_AND|B2|MID_SERIES 0  2e-13
RI0|_AND|B2|B I0|_AND|B2 I0|_AND|B2|MID_SHUNT  2.7439617672
LI0|_AND|B2|RB I0|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|B12|1 I0|_AND|B2 I0|_AND|B3 JJMIT AREA=1.7857142857142858
RI0|_AND|B12|B I0|_AND|B2 I0|_AND|B12|MID_SHUNT  3.84154647408
LI0|_AND|B12|RB I0|_AND|B12|MID_SHUNT I0|_AND|B3  2.1704737578552e-12
BI0|_AND|Q2|1 I0|_AND|Q2 I0|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q2|P I0|_AND|Q2|MID_SERIES 0  2e-13
RI0|_AND|Q2|B I0|_AND|Q2 I0|_AND|Q2|MID_SHUNT  2.7439617672
LI0|_AND|Q2|RB I0|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI0|_AND|Q1|1 I0|_AND|Q1 I0|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI0|_AND|Q1|P I0|_AND|Q1|MID_SERIES 0  2e-13
RI0|_AND|Q1|B I0|_AND|Q1 I0|_AND|Q1|MID_SHUNT  2.7439617672
LI0|_AND|Q1|RB I0|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_A|I_D1|B I1|_SPL_A|D1 I1|_SPL_A|I_D1|MID  2e-12
II1|_SPL_A|I_D1|B 0 I1|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_D2|B I1|_SPL_A|D2 I1|_SPL_A|I_D2|MID  2e-12
II1|_SPL_A|I_D2|B 0 I1|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_A|I_Q1|B I1|_SPL_A|QA1 I1|_SPL_A|I_Q1|MID  2e-12
II1|_SPL_A|I_Q1|B 0 I1|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_A|I_Q2|B I1|_SPL_A|QB1 I1|_SPL_A|I_Q2|MID  2e-12
II1|_SPL_A|I_Q2|B 0 I1|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_A|1|1 I1|_SPL_A|D1 I1|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|1|P I1|_SPL_A|1|MID_SERIES 0  2e-13
RI1|_SPL_A|1|B I1|_SPL_A|D1 I1|_SPL_A|1|MID_SHUNT  2.7439617672
LI1|_SPL_A|1|RB I1|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|2|1 I1|_SPL_A|D2 I1|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|2|P I1|_SPL_A|2|MID_SERIES 0  2e-13
RI1|_SPL_A|2|B I1|_SPL_A|D2 I1|_SPL_A|2|MID_SHUNT  2.7439617672
LI1|_SPL_A|2|RB I1|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|A|1 I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|A|P I1|_SPL_A|A|MID_SERIES 0  2e-13
RI1|_SPL_A|A|B I1|_SPL_A|QA1 I1|_SPL_A|A|MID_SHUNT  2.7439617672
LI1|_SPL_A|A|RB I1|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_A|B|1 I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_A|B|P I1|_SPL_A|B|MID_SERIES 0  2e-13
RI1|_SPL_A|B|B I1|_SPL_A|QB1 I1|_SPL_A|B|MID_SHUNT  2.7439617672
LI1|_SPL_A|B|RB I1|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI1|_SPL_B|I_D1|B I1|_SPL_B|D1 I1|_SPL_B|I_D1|MID  2e-12
II1|_SPL_B|I_D1|B 0 I1|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_D2|B I1|_SPL_B|D2 I1|_SPL_B|I_D2|MID  2e-12
II1|_SPL_B|I_D2|B 0 I1|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI1|_SPL_B|I_Q1|B I1|_SPL_B|QA1 I1|_SPL_B|I_Q1|MID  2e-12
II1|_SPL_B|I_Q1|B 0 I1|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI1|_SPL_B|I_Q2|B I1|_SPL_B|QB1 I1|_SPL_B|I_Q2|MID  2e-12
II1|_SPL_B|I_Q2|B 0 I1|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI1|_SPL_B|1|1 I1|_SPL_B|D1 I1|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|1|P I1|_SPL_B|1|MID_SERIES 0  2e-13
RI1|_SPL_B|1|B I1|_SPL_B|D1 I1|_SPL_B|1|MID_SHUNT  2.7439617672
LI1|_SPL_B|1|RB I1|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|2|1 I1|_SPL_B|D2 I1|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|2|P I1|_SPL_B|2|MID_SERIES 0  2e-13
RI1|_SPL_B|2|B I1|_SPL_B|D2 I1|_SPL_B|2|MID_SHUNT  2.7439617672
LI1|_SPL_B|2|RB I1|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|A|1 I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|A|P I1|_SPL_B|A|MID_SERIES 0  2e-13
RI1|_SPL_B|A|B I1|_SPL_B|QA1 I1|_SPL_B|A|MID_SHUNT  2.7439617672
LI1|_SPL_B|A|RB I1|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI1|_SPL_B|B|1 I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI1|_SPL_B|B|P I1|_SPL_B|B|MID_SERIES 0  2e-13
RI1|_SPL_B|B|B I1|_SPL_B|QB1 I1|_SPL_B|B|MID_SHUNT  2.7439617672
LI1|_SPL_B|B|RB I1|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_A|I_1|B I1|_DFF_A|A1 I1|_DFF_A|I_1|MID  2e-12
II1|_DFF_A|I_1|B 0 I1|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_3|B I1|_DFF_A|A3 I1|_DFF_A|I_3|MID  2e-12
II1|_DFF_A|I_3|B 0 I1|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_A|I_T|B I1|_DFF_A|T1 I1|_DFF_A|I_T|MID  2e-12
II1|_DFF_A|I_T|B 0 I1|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_A|I_6|B I1|_DFF_A|Q1 I1|_DFF_A|I_6|MID  2e-12
II1|_DFF_A|I_6|B 0 I1|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_A|1|1 I1|_DFF_A|A1 I1|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|1|P I1|_DFF_A|1|MID_SERIES 0  2e-13
RI1|_DFF_A|1|B I1|_DFF_A|A1 I1|_DFF_A|1|MID_SHUNT  2.7439617672
LI1|_DFF_A|1|RB I1|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|23|1 I1|_DFF_A|A2 I1|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|23|B I1|_DFF_A|A2 I1|_DFF_A|23|MID_SHUNT  3.84154647408
LI1|_DFF_A|23|RB I1|_DFF_A|23|MID_SHUNT I1|_DFF_A|A3  2.1704737578552e-12
BI1|_DFF_A|3|1 I1|_DFF_A|A3 I1|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|3|P I1|_DFF_A|3|MID_SERIES 0  2e-13
RI1|_DFF_A|3|B I1|_DFF_A|A3 I1|_DFF_A|3|MID_SHUNT  2.7439617672
LI1|_DFF_A|3|RB I1|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|4|1 I1|_DFF_A|A4 I1|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|4|P I1|_DFF_A|4|MID_SERIES 0  2e-13
RI1|_DFF_A|4|B I1|_DFF_A|A4 I1|_DFF_A|4|MID_SHUNT  2.7439617672
LI1|_DFF_A|4|RB I1|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|T|1 I1|_DFF_A|T1 I1|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|T|P I1|_DFF_A|T|MID_SERIES 0  2e-13
RI1|_DFF_A|T|B I1|_DFF_A|T1 I1|_DFF_A|T|MID_SHUNT  2.7439617672
LI1|_DFF_A|T|RB I1|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_A|45|1 I1|_DFF_A|T2 I1|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_A|45|B I1|_DFF_A|T2 I1|_DFF_A|45|MID_SHUNT  3.84154647408
LI1|_DFF_A|45|RB I1|_DFF_A|45|MID_SHUNT I1|_DFF_A|A4  2.1704737578552e-12
BI1|_DFF_A|6|1 I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_A|6|P I1|_DFF_A|6|MID_SERIES 0  2e-13
RI1|_DFF_A|6|B I1|_DFF_A|Q1 I1|_DFF_A|6|MID_SHUNT  2.7439617672
LI1|_DFF_A|6|RB I1|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI1|_DFF_B|I_1|B I1|_DFF_B|A1 I1|_DFF_B|I_1|MID  2e-12
II1|_DFF_B|I_1|B 0 I1|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_3|B I1|_DFF_B|A3 I1|_DFF_B|I_3|MID  2e-12
II1|_DFF_B|I_3|B 0 I1|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI1|_DFF_B|I_T|B I1|_DFF_B|T1 I1|_DFF_B|I_T|MID  2e-12
II1|_DFF_B|I_T|B 0 I1|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI1|_DFF_B|I_6|B I1|_DFF_B|Q1 I1|_DFF_B|I_6|MID  2e-12
II1|_DFF_B|I_6|B 0 I1|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI1|_DFF_B|1|1 I1|_DFF_B|A1 I1|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|1|P I1|_DFF_B|1|MID_SERIES 0  2e-13
RI1|_DFF_B|1|B I1|_DFF_B|A1 I1|_DFF_B|1|MID_SHUNT  2.7439617672
LI1|_DFF_B|1|RB I1|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|23|1 I1|_DFF_B|A2 I1|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|23|B I1|_DFF_B|A2 I1|_DFF_B|23|MID_SHUNT  3.84154647408
LI1|_DFF_B|23|RB I1|_DFF_B|23|MID_SHUNT I1|_DFF_B|A3  2.1704737578552e-12
BI1|_DFF_B|3|1 I1|_DFF_B|A3 I1|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|3|P I1|_DFF_B|3|MID_SERIES 0  2e-13
RI1|_DFF_B|3|B I1|_DFF_B|A3 I1|_DFF_B|3|MID_SHUNT  2.7439617672
LI1|_DFF_B|3|RB I1|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|4|1 I1|_DFF_B|A4 I1|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|4|P I1|_DFF_B|4|MID_SERIES 0  2e-13
RI1|_DFF_B|4|B I1|_DFF_B|A4 I1|_DFF_B|4|MID_SHUNT  2.7439617672
LI1|_DFF_B|4|RB I1|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|T|1 I1|_DFF_B|T1 I1|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|T|P I1|_DFF_B|T|MID_SERIES 0  2e-13
RI1|_DFF_B|T|B I1|_DFF_B|T1 I1|_DFF_B|T|MID_SHUNT  2.7439617672
LI1|_DFF_B|T|RB I1|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI1|_DFF_B|45|1 I1|_DFF_B|T2 I1|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI1|_DFF_B|45|B I1|_DFF_B|T2 I1|_DFF_B|45|MID_SHUNT  3.84154647408
LI1|_DFF_B|45|RB I1|_DFF_B|45|MID_SHUNT I1|_DFF_B|A4  2.1704737578552e-12
BI1|_DFF_B|6|1 I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI1|_DFF_B|6|P I1|_DFF_B|6|MID_SERIES 0  2e-13
RI1|_DFF_B|6|B I1|_DFF_B|Q1 I1|_DFF_B|6|MID_SHUNT  2.7439617672
LI1|_DFF_B|6|RB I1|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI1|_XOR|I_A1|B I1|_XOR|A1 I1|_XOR|I_A1|MID  2e-12
II1|_XOR|I_A1|B 0 I1|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_A3|B I1|_XOR|A3 I1|_XOR|I_A3|MID  2e-12
II1|_XOR|I_A3|B 0 I1|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B1|B I1|_XOR|B1 I1|_XOR|I_B1|MID  2e-12
II1|_XOR|I_B1|B 0 I1|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_B3|B I1|_XOR|B3 I1|_XOR|I_B3|MID  2e-12
II1|_XOR|I_B3|B 0 I1|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI1|_XOR|I_Q1|B I1|_XOR|Q1 I1|_XOR|I_Q1|MID  2e-12
II1|_XOR|I_Q1|B 0 I1|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_XOR|A1|1 I1|_XOR|A1 I1|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A1|P I1|_XOR|A1|MID_SERIES 0  5e-13
RI1|_XOR|A1|B I1|_XOR|A1 I1|_XOR|A1|MID_SHUNT  2.7439617672
LI1|_XOR|A1|RB I1|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A2|1 I1|_XOR|A2 I1|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A2|P I1|_XOR|A2|MID_SERIES 0  5e-13
RI1|_XOR|A2|B I1|_XOR|A2 I1|_XOR|A2|MID_SHUNT  2.7439617672
LI1|_XOR|A2|RB I1|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|A3|1 I1|_XOR|A2 I1|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|A3|P I1|_XOR|A3|MID_SERIES I1|_XOR|A3  1.2e-12
RI1|_XOR|A3|B I1|_XOR|A2 I1|_XOR|A3|MID_SHUNT  2.7439617672
LI1|_XOR|A3|RB I1|_XOR|A3|MID_SHUNT I1|_XOR|A3  2.050338398468e-12
BI1|_XOR|B1|1 I1|_XOR|B1 I1|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B1|P I1|_XOR|B1|MID_SERIES 0  5e-13
RI1|_XOR|B1|B I1|_XOR|B1 I1|_XOR|B1|MID_SHUNT  2.7439617672
LI1|_XOR|B1|RB I1|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B2|1 I1|_XOR|B2 I1|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B2|P I1|_XOR|B2|MID_SERIES 0  5e-13
RI1|_XOR|B2|B I1|_XOR|B2 I1|_XOR|B2|MID_SHUNT  2.7439617672
LI1|_XOR|B2|RB I1|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|B3|1 I1|_XOR|B2 I1|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|B3|P I1|_XOR|B3|MID_SERIES I1|_XOR|B3  1.2e-12
RI1|_XOR|B3|B I1|_XOR|B2 I1|_XOR|B3|MID_SHUNT  2.7439617672
LI1|_XOR|B3|RB I1|_XOR|B3|MID_SHUNT I1|_XOR|B3  2.050338398468e-12
BI1|_XOR|T1|1 I1|_XOR|T1 I1|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|T1|P I1|_XOR|T1|MID_SERIES 0  5e-13
RI1|_XOR|T1|B I1|_XOR|T1 I1|_XOR|T1|MID_SHUNT  2.7439617672
LI1|_XOR|T1|RB I1|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|T2|1 I1|_XOR|T2 I1|_XOR|ABTQ JJMIT AREA=2.0
RI1|_XOR|T2|B I1|_XOR|T2 I1|_XOR|T2|MID_SHUNT  3.429952209
LI1|_XOR|T2|RB I1|_XOR|T2|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|AB|1 I1|_XOR|AB I1|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI1|_XOR|AB|P I1|_XOR|AB|MID_SERIES I1|_XOR|ABTQ  1.2e-12
RI1|_XOR|AB|B I1|_XOR|AB I1|_XOR|AB|MID_SHUNT  3.429952209
LI1|_XOR|AB|RB I1|_XOR|AB|MID_SHUNT I1|_XOR|ABTQ  2.437922998085e-12
BI1|_XOR|ABTQ|1 I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|ABTQ|P I1|_XOR|ABTQ|MID_SERIES 0  5e-13
RI1|_XOR|ABTQ|B I1|_XOR|ABTQ I1|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI1|_XOR|ABTQ|RB I1|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI1|_XOR|Q1|1 I1|_XOR|Q1 I1|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_XOR|Q1|P I1|_XOR|Q1|MID_SERIES 0  5e-13
RI1|_XOR|Q1|B I1|_XOR|Q1 I1|_XOR|Q1|MID_SHUNT  2.7439617672
LI1|_XOR|Q1|RB I1|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI1|_AND|I_A1|B I1|_AND|A1 I1|_AND|I_A1|MID  2e-12
II1|_AND|I_A1|B 0 I1|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_B1|B I1|_AND|B1 I1|_AND|I_B1|MID  2e-12
II1|_AND|I_B1|B 0 I1|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q3|B I1|_AND|Q3 I1|_AND|I_Q3|MID  2e-12
II1|_AND|I_Q3|B 0 I1|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI1|_AND|I_Q2|B I1|_AND|Q2 I1|_AND|I_Q2|MID  2e-12
II1|_AND|I_Q2|B 0 I1|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI1|_AND|I_Q1|B I1|_AND|Q1 I1|_AND|I_Q1|MID  2e-12
II1|_AND|I_Q1|B 0 I1|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI1|_AND|A1|1 I1|_AND|A1 I1|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A1|P I1|_AND|A1|MID_SERIES 0  2e-13
RI1|_AND|A1|B I1|_AND|A1 I1|_AND|A1|MID_SHUNT  2.7439617672
LI1|_AND|A1|RB I1|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A2|1 I1|_AND|A2 I1|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|A2|P I1|_AND|A2|MID_SERIES 0  2e-13
RI1|_AND|A2|B I1|_AND|A2 I1|_AND|A2|MID_SHUNT  2.7439617672
LI1|_AND|A2|RB I1|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|A12|1 I1|_AND|A2 I1|_AND|A3 JJMIT AREA=1.7857142857142858
RI1|_AND|A12|B I1|_AND|A2 I1|_AND|A12|MID_SHUNT  3.84154647408
LI1|_AND|A12|RB I1|_AND|A12|MID_SHUNT I1|_AND|A3  2.1704737578552e-12
BI1|_AND|B1|1 I1|_AND|B1 I1|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B1|P I1|_AND|B1|MID_SERIES 0  2e-13
RI1|_AND|B1|B I1|_AND|B1 I1|_AND|B1|MID_SHUNT  2.7439617672
LI1|_AND|B1|RB I1|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B2|1 I1|_AND|B2 I1|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|B2|P I1|_AND|B2|MID_SERIES 0  2e-13
RI1|_AND|B2|B I1|_AND|B2 I1|_AND|B2|MID_SHUNT  2.7439617672
LI1|_AND|B2|RB I1|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|B12|1 I1|_AND|B2 I1|_AND|B3 JJMIT AREA=1.7857142857142858
RI1|_AND|B12|B I1|_AND|B2 I1|_AND|B12|MID_SHUNT  3.84154647408
LI1|_AND|B12|RB I1|_AND|B12|MID_SHUNT I1|_AND|B3  2.1704737578552e-12
BI1|_AND|Q2|1 I1|_AND|Q2 I1|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q2|P I1|_AND|Q2|MID_SERIES 0  2e-13
RI1|_AND|Q2|B I1|_AND|Q2 I1|_AND|Q2|MID_SHUNT  2.7439617672
LI1|_AND|Q2|RB I1|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI1|_AND|Q1|1 I1|_AND|Q1 I1|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI1|_AND|Q1|P I1|_AND|Q1|MID_SERIES 0  2e-13
RI1|_AND|Q1|B I1|_AND|Q1 I1|_AND|Q1|MID_SHUNT  2.7439617672
LI1|_AND|Q1|RB I1|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_A|I_D1|B I2|_SPL_A|D1 I2|_SPL_A|I_D1|MID  2e-12
II2|_SPL_A|I_D1|B 0 I2|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_D2|B I2|_SPL_A|D2 I2|_SPL_A|I_D2|MID  2e-12
II2|_SPL_A|I_D2|B 0 I2|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_A|I_Q1|B I2|_SPL_A|QA1 I2|_SPL_A|I_Q1|MID  2e-12
II2|_SPL_A|I_Q1|B 0 I2|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_A|I_Q2|B I2|_SPL_A|QB1 I2|_SPL_A|I_Q2|MID  2e-12
II2|_SPL_A|I_Q2|B 0 I2|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_A|1|1 I2|_SPL_A|D1 I2|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|1|P I2|_SPL_A|1|MID_SERIES 0  2e-13
RI2|_SPL_A|1|B I2|_SPL_A|D1 I2|_SPL_A|1|MID_SHUNT  2.7439617672
LI2|_SPL_A|1|RB I2|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|2|1 I2|_SPL_A|D2 I2|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|2|P I2|_SPL_A|2|MID_SERIES 0  2e-13
RI2|_SPL_A|2|B I2|_SPL_A|D2 I2|_SPL_A|2|MID_SHUNT  2.7439617672
LI2|_SPL_A|2|RB I2|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|A|1 I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|A|P I2|_SPL_A|A|MID_SERIES 0  2e-13
RI2|_SPL_A|A|B I2|_SPL_A|QA1 I2|_SPL_A|A|MID_SHUNT  2.7439617672
LI2|_SPL_A|A|RB I2|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_A|B|1 I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_A|B|P I2|_SPL_A|B|MID_SERIES 0  2e-13
RI2|_SPL_A|B|B I2|_SPL_A|QB1 I2|_SPL_A|B|MID_SHUNT  2.7439617672
LI2|_SPL_A|B|RB I2|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI2|_SPL_B|I_D1|B I2|_SPL_B|D1 I2|_SPL_B|I_D1|MID  2e-12
II2|_SPL_B|I_D1|B 0 I2|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_D2|B I2|_SPL_B|D2 I2|_SPL_B|I_D2|MID  2e-12
II2|_SPL_B|I_D2|B 0 I2|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI2|_SPL_B|I_Q1|B I2|_SPL_B|QA1 I2|_SPL_B|I_Q1|MID  2e-12
II2|_SPL_B|I_Q1|B 0 I2|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI2|_SPL_B|I_Q2|B I2|_SPL_B|QB1 I2|_SPL_B|I_Q2|MID  2e-12
II2|_SPL_B|I_Q2|B 0 I2|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI2|_SPL_B|1|1 I2|_SPL_B|D1 I2|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|1|P I2|_SPL_B|1|MID_SERIES 0  2e-13
RI2|_SPL_B|1|B I2|_SPL_B|D1 I2|_SPL_B|1|MID_SHUNT  2.7439617672
LI2|_SPL_B|1|RB I2|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|2|1 I2|_SPL_B|D2 I2|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|2|P I2|_SPL_B|2|MID_SERIES 0  2e-13
RI2|_SPL_B|2|B I2|_SPL_B|D2 I2|_SPL_B|2|MID_SHUNT  2.7439617672
LI2|_SPL_B|2|RB I2|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|A|1 I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|A|P I2|_SPL_B|A|MID_SERIES 0  2e-13
RI2|_SPL_B|A|B I2|_SPL_B|QA1 I2|_SPL_B|A|MID_SHUNT  2.7439617672
LI2|_SPL_B|A|RB I2|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI2|_SPL_B|B|1 I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI2|_SPL_B|B|P I2|_SPL_B|B|MID_SERIES 0  2e-13
RI2|_SPL_B|B|B I2|_SPL_B|QB1 I2|_SPL_B|B|MID_SHUNT  2.7439617672
LI2|_SPL_B|B|RB I2|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_A|I_1|B I2|_DFF_A|A1 I2|_DFF_A|I_1|MID  2e-12
II2|_DFF_A|I_1|B 0 I2|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_3|B I2|_DFF_A|A3 I2|_DFF_A|I_3|MID  2e-12
II2|_DFF_A|I_3|B 0 I2|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_A|I_T|B I2|_DFF_A|T1 I2|_DFF_A|I_T|MID  2e-12
II2|_DFF_A|I_T|B 0 I2|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_A|I_6|B I2|_DFF_A|Q1 I2|_DFF_A|I_6|MID  2e-12
II2|_DFF_A|I_6|B 0 I2|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_A|1|1 I2|_DFF_A|A1 I2|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|1|P I2|_DFF_A|1|MID_SERIES 0  2e-13
RI2|_DFF_A|1|B I2|_DFF_A|A1 I2|_DFF_A|1|MID_SHUNT  2.7439617672
LI2|_DFF_A|1|RB I2|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|23|1 I2|_DFF_A|A2 I2|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|23|B I2|_DFF_A|A2 I2|_DFF_A|23|MID_SHUNT  3.84154647408
LI2|_DFF_A|23|RB I2|_DFF_A|23|MID_SHUNT I2|_DFF_A|A3  2.1704737578552e-12
BI2|_DFF_A|3|1 I2|_DFF_A|A3 I2|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|3|P I2|_DFF_A|3|MID_SERIES 0  2e-13
RI2|_DFF_A|3|B I2|_DFF_A|A3 I2|_DFF_A|3|MID_SHUNT  2.7439617672
LI2|_DFF_A|3|RB I2|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|4|1 I2|_DFF_A|A4 I2|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|4|P I2|_DFF_A|4|MID_SERIES 0  2e-13
RI2|_DFF_A|4|B I2|_DFF_A|A4 I2|_DFF_A|4|MID_SHUNT  2.7439617672
LI2|_DFF_A|4|RB I2|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|T|1 I2|_DFF_A|T1 I2|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|T|P I2|_DFF_A|T|MID_SERIES 0  2e-13
RI2|_DFF_A|T|B I2|_DFF_A|T1 I2|_DFF_A|T|MID_SHUNT  2.7439617672
LI2|_DFF_A|T|RB I2|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_A|45|1 I2|_DFF_A|T2 I2|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_A|45|B I2|_DFF_A|T2 I2|_DFF_A|45|MID_SHUNT  3.84154647408
LI2|_DFF_A|45|RB I2|_DFF_A|45|MID_SHUNT I2|_DFF_A|A4  2.1704737578552e-12
BI2|_DFF_A|6|1 I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_A|6|P I2|_DFF_A|6|MID_SERIES 0  2e-13
RI2|_DFF_A|6|B I2|_DFF_A|Q1 I2|_DFF_A|6|MID_SHUNT  2.7439617672
LI2|_DFF_A|6|RB I2|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI2|_DFF_B|I_1|B I2|_DFF_B|A1 I2|_DFF_B|I_1|MID  2e-12
II2|_DFF_B|I_1|B 0 I2|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_3|B I2|_DFF_B|A3 I2|_DFF_B|I_3|MID  2e-12
II2|_DFF_B|I_3|B 0 I2|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI2|_DFF_B|I_T|B I2|_DFF_B|T1 I2|_DFF_B|I_T|MID  2e-12
II2|_DFF_B|I_T|B 0 I2|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI2|_DFF_B|I_6|B I2|_DFF_B|Q1 I2|_DFF_B|I_6|MID  2e-12
II2|_DFF_B|I_6|B 0 I2|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI2|_DFF_B|1|1 I2|_DFF_B|A1 I2|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|1|P I2|_DFF_B|1|MID_SERIES 0  2e-13
RI2|_DFF_B|1|B I2|_DFF_B|A1 I2|_DFF_B|1|MID_SHUNT  2.7439617672
LI2|_DFF_B|1|RB I2|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|23|1 I2|_DFF_B|A2 I2|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|23|B I2|_DFF_B|A2 I2|_DFF_B|23|MID_SHUNT  3.84154647408
LI2|_DFF_B|23|RB I2|_DFF_B|23|MID_SHUNT I2|_DFF_B|A3  2.1704737578552e-12
BI2|_DFF_B|3|1 I2|_DFF_B|A3 I2|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|3|P I2|_DFF_B|3|MID_SERIES 0  2e-13
RI2|_DFF_B|3|B I2|_DFF_B|A3 I2|_DFF_B|3|MID_SHUNT  2.7439617672
LI2|_DFF_B|3|RB I2|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|4|1 I2|_DFF_B|A4 I2|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|4|P I2|_DFF_B|4|MID_SERIES 0  2e-13
RI2|_DFF_B|4|B I2|_DFF_B|A4 I2|_DFF_B|4|MID_SHUNT  2.7439617672
LI2|_DFF_B|4|RB I2|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|T|1 I2|_DFF_B|T1 I2|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|T|P I2|_DFF_B|T|MID_SERIES 0  2e-13
RI2|_DFF_B|T|B I2|_DFF_B|T1 I2|_DFF_B|T|MID_SHUNT  2.7439617672
LI2|_DFF_B|T|RB I2|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI2|_DFF_B|45|1 I2|_DFF_B|T2 I2|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI2|_DFF_B|45|B I2|_DFF_B|T2 I2|_DFF_B|45|MID_SHUNT  3.84154647408
LI2|_DFF_B|45|RB I2|_DFF_B|45|MID_SHUNT I2|_DFF_B|A4  2.1704737578552e-12
BI2|_DFF_B|6|1 I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI2|_DFF_B|6|P I2|_DFF_B|6|MID_SERIES 0  2e-13
RI2|_DFF_B|6|B I2|_DFF_B|Q1 I2|_DFF_B|6|MID_SHUNT  2.7439617672
LI2|_DFF_B|6|RB I2|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI2|_XOR|I_A1|B I2|_XOR|A1 I2|_XOR|I_A1|MID  2e-12
II2|_XOR|I_A1|B 0 I2|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_A3|B I2|_XOR|A3 I2|_XOR|I_A3|MID  2e-12
II2|_XOR|I_A3|B 0 I2|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B1|B I2|_XOR|B1 I2|_XOR|I_B1|MID  2e-12
II2|_XOR|I_B1|B 0 I2|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_B3|B I2|_XOR|B3 I2|_XOR|I_B3|MID  2e-12
II2|_XOR|I_B3|B 0 I2|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI2|_XOR|I_Q1|B I2|_XOR|Q1 I2|_XOR|I_Q1|MID  2e-12
II2|_XOR|I_Q1|B 0 I2|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_XOR|A1|1 I2|_XOR|A1 I2|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A1|P I2|_XOR|A1|MID_SERIES 0  5e-13
RI2|_XOR|A1|B I2|_XOR|A1 I2|_XOR|A1|MID_SHUNT  2.7439617672
LI2|_XOR|A1|RB I2|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A2|1 I2|_XOR|A2 I2|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A2|P I2|_XOR|A2|MID_SERIES 0  5e-13
RI2|_XOR|A2|B I2|_XOR|A2 I2|_XOR|A2|MID_SHUNT  2.7439617672
LI2|_XOR|A2|RB I2|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|A3|1 I2|_XOR|A2 I2|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|A3|P I2|_XOR|A3|MID_SERIES I2|_XOR|A3  1.2e-12
RI2|_XOR|A3|B I2|_XOR|A2 I2|_XOR|A3|MID_SHUNT  2.7439617672
LI2|_XOR|A3|RB I2|_XOR|A3|MID_SHUNT I2|_XOR|A3  2.050338398468e-12
BI2|_XOR|B1|1 I2|_XOR|B1 I2|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B1|P I2|_XOR|B1|MID_SERIES 0  5e-13
RI2|_XOR|B1|B I2|_XOR|B1 I2|_XOR|B1|MID_SHUNT  2.7439617672
LI2|_XOR|B1|RB I2|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B2|1 I2|_XOR|B2 I2|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B2|P I2|_XOR|B2|MID_SERIES 0  5e-13
RI2|_XOR|B2|B I2|_XOR|B2 I2|_XOR|B2|MID_SHUNT  2.7439617672
LI2|_XOR|B2|RB I2|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|B3|1 I2|_XOR|B2 I2|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|B3|P I2|_XOR|B3|MID_SERIES I2|_XOR|B3  1.2e-12
RI2|_XOR|B3|B I2|_XOR|B2 I2|_XOR|B3|MID_SHUNT  2.7439617672
LI2|_XOR|B3|RB I2|_XOR|B3|MID_SHUNT I2|_XOR|B3  2.050338398468e-12
BI2|_XOR|T1|1 I2|_XOR|T1 I2|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|T1|P I2|_XOR|T1|MID_SERIES 0  5e-13
RI2|_XOR|T1|B I2|_XOR|T1 I2|_XOR|T1|MID_SHUNT  2.7439617672
LI2|_XOR|T1|RB I2|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|T2|1 I2|_XOR|T2 I2|_XOR|ABTQ JJMIT AREA=2.0
RI2|_XOR|T2|B I2|_XOR|T2 I2|_XOR|T2|MID_SHUNT  3.429952209
LI2|_XOR|T2|RB I2|_XOR|T2|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|AB|1 I2|_XOR|AB I2|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI2|_XOR|AB|P I2|_XOR|AB|MID_SERIES I2|_XOR|ABTQ  1.2e-12
RI2|_XOR|AB|B I2|_XOR|AB I2|_XOR|AB|MID_SHUNT  3.429952209
LI2|_XOR|AB|RB I2|_XOR|AB|MID_SHUNT I2|_XOR|ABTQ  2.437922998085e-12
BI2|_XOR|ABTQ|1 I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|ABTQ|P I2|_XOR|ABTQ|MID_SERIES 0  5e-13
RI2|_XOR|ABTQ|B I2|_XOR|ABTQ I2|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI2|_XOR|ABTQ|RB I2|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI2|_XOR|Q1|1 I2|_XOR|Q1 I2|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_XOR|Q1|P I2|_XOR|Q1|MID_SERIES 0  5e-13
RI2|_XOR|Q1|B I2|_XOR|Q1 I2|_XOR|Q1|MID_SHUNT  2.7439617672
LI2|_XOR|Q1|RB I2|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI2|_AND|I_A1|B I2|_AND|A1 I2|_AND|I_A1|MID  2e-12
II2|_AND|I_A1|B 0 I2|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_B1|B I2|_AND|B1 I2|_AND|I_B1|MID  2e-12
II2|_AND|I_B1|B 0 I2|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q3|B I2|_AND|Q3 I2|_AND|I_Q3|MID  2e-12
II2|_AND|I_Q3|B 0 I2|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI2|_AND|I_Q2|B I2|_AND|Q2 I2|_AND|I_Q2|MID  2e-12
II2|_AND|I_Q2|B 0 I2|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI2|_AND|I_Q1|B I2|_AND|Q1 I2|_AND|I_Q1|MID  2e-12
II2|_AND|I_Q1|B 0 I2|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI2|_AND|A1|1 I2|_AND|A1 I2|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A1|P I2|_AND|A1|MID_SERIES 0  2e-13
RI2|_AND|A1|B I2|_AND|A1 I2|_AND|A1|MID_SHUNT  2.7439617672
LI2|_AND|A1|RB I2|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A2|1 I2|_AND|A2 I2|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|A2|P I2|_AND|A2|MID_SERIES 0  2e-13
RI2|_AND|A2|B I2|_AND|A2 I2|_AND|A2|MID_SHUNT  2.7439617672
LI2|_AND|A2|RB I2|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|A12|1 I2|_AND|A2 I2|_AND|A3 JJMIT AREA=1.7857142857142858
RI2|_AND|A12|B I2|_AND|A2 I2|_AND|A12|MID_SHUNT  3.84154647408
LI2|_AND|A12|RB I2|_AND|A12|MID_SHUNT I2|_AND|A3  2.1704737578552e-12
BI2|_AND|B1|1 I2|_AND|B1 I2|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B1|P I2|_AND|B1|MID_SERIES 0  2e-13
RI2|_AND|B1|B I2|_AND|B1 I2|_AND|B1|MID_SHUNT  2.7439617672
LI2|_AND|B1|RB I2|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B2|1 I2|_AND|B2 I2|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|B2|P I2|_AND|B2|MID_SERIES 0  2e-13
RI2|_AND|B2|B I2|_AND|B2 I2|_AND|B2|MID_SHUNT  2.7439617672
LI2|_AND|B2|RB I2|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|B12|1 I2|_AND|B2 I2|_AND|B3 JJMIT AREA=1.7857142857142858
RI2|_AND|B12|B I2|_AND|B2 I2|_AND|B12|MID_SHUNT  3.84154647408
LI2|_AND|B12|RB I2|_AND|B12|MID_SHUNT I2|_AND|B3  2.1704737578552e-12
BI2|_AND|Q2|1 I2|_AND|Q2 I2|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q2|P I2|_AND|Q2|MID_SERIES 0  2e-13
RI2|_AND|Q2|B I2|_AND|Q2 I2|_AND|Q2|MID_SHUNT  2.7439617672
LI2|_AND|Q2|RB I2|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI2|_AND|Q1|1 I2|_AND|Q1 I2|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI2|_AND|Q1|P I2|_AND|Q1|MID_SERIES 0  2e-13
RI2|_AND|Q1|B I2|_AND|Q1 I2|_AND|Q1|MID_SHUNT  2.7439617672
LI2|_AND|Q1|RB I2|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_A|I_D1|B I3|_SPL_A|D1 I3|_SPL_A|I_D1|MID  2e-12
II3|_SPL_A|I_D1|B 0 I3|_SPL_A|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_D2|B I3|_SPL_A|D2 I3|_SPL_A|I_D2|MID  2e-12
II3|_SPL_A|I_D2|B 0 I3|_SPL_A|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_A|I_Q1|B I3|_SPL_A|QA1 I3|_SPL_A|I_Q1|MID  2e-12
II3|_SPL_A|I_Q1|B 0 I3|_SPL_A|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_A|I_Q2|B I3|_SPL_A|QB1 I3|_SPL_A|I_Q2|MID  2e-12
II3|_SPL_A|I_Q2|B 0 I3|_SPL_A|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_A|1|1 I3|_SPL_A|D1 I3|_SPL_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|1|P I3|_SPL_A|1|MID_SERIES 0  2e-13
RI3|_SPL_A|1|B I3|_SPL_A|D1 I3|_SPL_A|1|MID_SHUNT  2.7439617672
LI3|_SPL_A|1|RB I3|_SPL_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|2|1 I3|_SPL_A|D2 I3|_SPL_A|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|2|P I3|_SPL_A|2|MID_SERIES 0  2e-13
RI3|_SPL_A|2|B I3|_SPL_A|D2 I3|_SPL_A|2|MID_SHUNT  2.7439617672
LI3|_SPL_A|2|RB I3|_SPL_A|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|A|1 I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|A|P I3|_SPL_A|A|MID_SERIES 0  2e-13
RI3|_SPL_A|A|B I3|_SPL_A|QA1 I3|_SPL_A|A|MID_SHUNT  2.7439617672
LI3|_SPL_A|A|RB I3|_SPL_A|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_A|B|1 I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_A|B|P I3|_SPL_A|B|MID_SERIES 0  2e-13
RI3|_SPL_A|B|B I3|_SPL_A|QB1 I3|_SPL_A|B|MID_SHUNT  2.7439617672
LI3|_SPL_A|B|RB I3|_SPL_A|B|MID_SHUNT 0  1.550338398468e-12
LI3|_SPL_B|I_D1|B I3|_SPL_B|D1 I3|_SPL_B|I_D1|MID  2e-12
II3|_SPL_B|I_D1|B 0 I3|_SPL_B|I_D1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_D2|B I3|_SPL_B|D2 I3|_SPL_B|I_D2|MID  2e-12
II3|_SPL_B|I_D2|B 0 I3|_SPL_B|I_D2|MID  PWL(0 0 5e-12 0.0002205)
LI3|_SPL_B|I_Q1|B I3|_SPL_B|QA1 I3|_SPL_B|I_Q1|MID  2e-12
II3|_SPL_B|I_Q1|B 0 I3|_SPL_B|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
LI3|_SPL_B|I_Q2|B I3|_SPL_B|QB1 I3|_SPL_B|I_Q2|MID  2e-12
II3|_SPL_B|I_Q2|B 0 I3|_SPL_B|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
BI3|_SPL_B|1|1 I3|_SPL_B|D1 I3|_SPL_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|1|P I3|_SPL_B|1|MID_SERIES 0  2e-13
RI3|_SPL_B|1|B I3|_SPL_B|D1 I3|_SPL_B|1|MID_SHUNT  2.7439617672
LI3|_SPL_B|1|RB I3|_SPL_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|2|1 I3|_SPL_B|D2 I3|_SPL_B|2|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|2|P I3|_SPL_B|2|MID_SERIES 0  2e-13
RI3|_SPL_B|2|B I3|_SPL_B|D2 I3|_SPL_B|2|MID_SHUNT  2.7439617672
LI3|_SPL_B|2|RB I3|_SPL_B|2|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|A|1 I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|A|P I3|_SPL_B|A|MID_SERIES 0  2e-13
RI3|_SPL_B|A|B I3|_SPL_B|QA1 I3|_SPL_B|A|MID_SHUNT  2.7439617672
LI3|_SPL_B|A|RB I3|_SPL_B|A|MID_SHUNT 0  1.550338398468e-12
BI3|_SPL_B|B|1 I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SERIES JJMIT AREA=2.5
LI3|_SPL_B|B|P I3|_SPL_B|B|MID_SERIES 0  2e-13
RI3|_SPL_B|B|B I3|_SPL_B|QB1 I3|_SPL_B|B|MID_SHUNT  2.7439617672
LI3|_SPL_B|B|RB I3|_SPL_B|B|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_A|I_1|B I3|_DFF_A|A1 I3|_DFF_A|I_1|MID  2e-12
II3|_DFF_A|I_1|B 0 I3|_DFF_A|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_3|B I3|_DFF_A|A3 I3|_DFF_A|I_3|MID  2e-12
II3|_DFF_A|I_3|B 0 I3|_DFF_A|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_A|I_T|B I3|_DFF_A|T1 I3|_DFF_A|I_T|MID  2e-12
II3|_DFF_A|I_T|B 0 I3|_DFF_A|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_A|I_6|B I3|_DFF_A|Q1 I3|_DFF_A|I_6|MID  2e-12
II3|_DFF_A|I_6|B 0 I3|_DFF_A|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_A|1|1 I3|_DFF_A|A1 I3|_DFF_A|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|1|P I3|_DFF_A|1|MID_SERIES 0  2e-13
RI3|_DFF_A|1|B I3|_DFF_A|A1 I3|_DFF_A|1|MID_SHUNT  2.7439617672
LI3|_DFF_A|1|RB I3|_DFF_A|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|23|1 I3|_DFF_A|A2 I3|_DFF_A|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|23|B I3|_DFF_A|A2 I3|_DFF_A|23|MID_SHUNT  3.84154647408
LI3|_DFF_A|23|RB I3|_DFF_A|23|MID_SHUNT I3|_DFF_A|A3  2.1704737578552e-12
BI3|_DFF_A|3|1 I3|_DFF_A|A3 I3|_DFF_A|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|3|P I3|_DFF_A|3|MID_SERIES 0  2e-13
RI3|_DFF_A|3|B I3|_DFF_A|A3 I3|_DFF_A|3|MID_SHUNT  2.7439617672
LI3|_DFF_A|3|RB I3|_DFF_A|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|4|1 I3|_DFF_A|A4 I3|_DFF_A|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|4|P I3|_DFF_A|4|MID_SERIES 0  2e-13
RI3|_DFF_A|4|B I3|_DFF_A|A4 I3|_DFF_A|4|MID_SHUNT  2.7439617672
LI3|_DFF_A|4|RB I3|_DFF_A|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|T|1 I3|_DFF_A|T1 I3|_DFF_A|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|T|P I3|_DFF_A|T|MID_SERIES 0  2e-13
RI3|_DFF_A|T|B I3|_DFF_A|T1 I3|_DFF_A|T|MID_SHUNT  2.7439617672
LI3|_DFF_A|T|RB I3|_DFF_A|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_A|45|1 I3|_DFF_A|T2 I3|_DFF_A|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_A|45|B I3|_DFF_A|T2 I3|_DFF_A|45|MID_SHUNT  3.84154647408
LI3|_DFF_A|45|RB I3|_DFF_A|45|MID_SHUNT I3|_DFF_A|A4  2.1704737578552e-12
BI3|_DFF_A|6|1 I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_A|6|P I3|_DFF_A|6|MID_SERIES 0  2e-13
RI3|_DFF_A|6|B I3|_DFF_A|Q1 I3|_DFF_A|6|MID_SHUNT  2.7439617672
LI3|_DFF_A|6|RB I3|_DFF_A|6|MID_SHUNT 0  1.550338398468e-12
LI3|_DFF_B|I_1|B I3|_DFF_B|A1 I3|_DFF_B|I_1|MID  2e-12
II3|_DFF_B|I_1|B 0 I3|_DFF_B|I_1|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_3|B I3|_DFF_B|A3 I3|_DFF_B|I_3|MID  2e-12
II3|_DFF_B|I_3|B 0 I3|_DFF_B|I_3|MID  PWL(0 0 5e-12 0.00025)
LI3|_DFF_B|I_T|B I3|_DFF_B|T1 I3|_DFF_B|I_T|MID  2e-12
II3|_DFF_B|I_T|B 0 I3|_DFF_B|I_T|MID  PWL(0 0 5e-12 0.000175)
LI3|_DFF_B|I_6|B I3|_DFF_B|Q1 I3|_DFF_B|I_6|MID  2e-12
II3|_DFF_B|I_6|B 0 I3|_DFF_B|I_6|MID  PWL(0 0 5e-12 0.000175)
BI3|_DFF_B|1|1 I3|_DFF_B|A1 I3|_DFF_B|1|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|1|P I3|_DFF_B|1|MID_SERIES 0  2e-13
RI3|_DFF_B|1|B I3|_DFF_B|A1 I3|_DFF_B|1|MID_SHUNT  2.7439617672
LI3|_DFF_B|1|RB I3|_DFF_B|1|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|23|1 I3|_DFF_B|A2 I3|_DFF_B|A3 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|23|B I3|_DFF_B|A2 I3|_DFF_B|23|MID_SHUNT  3.84154647408
LI3|_DFF_B|23|RB I3|_DFF_B|23|MID_SHUNT I3|_DFF_B|A3  2.1704737578552e-12
BI3|_DFF_B|3|1 I3|_DFF_B|A3 I3|_DFF_B|3|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|3|P I3|_DFF_B|3|MID_SERIES 0  2e-13
RI3|_DFF_B|3|B I3|_DFF_B|A3 I3|_DFF_B|3|MID_SHUNT  2.7439617672
LI3|_DFF_B|3|RB I3|_DFF_B|3|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|4|1 I3|_DFF_B|A4 I3|_DFF_B|4|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|4|P I3|_DFF_B|4|MID_SERIES 0  2e-13
RI3|_DFF_B|4|B I3|_DFF_B|A4 I3|_DFF_B|4|MID_SHUNT  2.7439617672
LI3|_DFF_B|4|RB I3|_DFF_B|4|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|T|1 I3|_DFF_B|T1 I3|_DFF_B|T|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|T|P I3|_DFF_B|T|MID_SERIES 0  2e-13
RI3|_DFF_B|T|B I3|_DFF_B|T1 I3|_DFF_B|T|MID_SHUNT  2.7439617672
LI3|_DFF_B|T|RB I3|_DFF_B|T|MID_SHUNT 0  1.550338398468e-12
BI3|_DFF_B|45|1 I3|_DFF_B|T2 I3|_DFF_B|A4 JJMIT AREA=1.7857142857142858
RI3|_DFF_B|45|B I3|_DFF_B|T2 I3|_DFF_B|45|MID_SHUNT  3.84154647408
LI3|_DFF_B|45|RB I3|_DFF_B|45|MID_SHUNT I3|_DFF_B|A4  2.1704737578552e-12
BI3|_DFF_B|6|1 I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SERIES JJMIT AREA=2.5
LI3|_DFF_B|6|P I3|_DFF_B|6|MID_SERIES 0  2e-13
RI3|_DFF_B|6|B I3|_DFF_B|Q1 I3|_DFF_B|6|MID_SHUNT  2.7439617672
LI3|_DFF_B|6|RB I3|_DFF_B|6|MID_SHUNT 0  1.550338398468e-12
LI3|_XOR|I_A1|B I3|_XOR|A1 I3|_XOR|I_A1|MID  2e-12
II3|_XOR|I_A1|B 0 I3|_XOR|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_A3|B I3|_XOR|A3 I3|_XOR|I_A3|MID  2e-12
II3|_XOR|I_A3|B 0 I3|_XOR|I_A3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B1|B I3|_XOR|B1 I3|_XOR|I_B1|MID  2e-12
II3|_XOR|I_B1|B 0 I3|_XOR|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_B3|B I3|_XOR|B3 I3|_XOR|I_B3|MID  2e-12
II3|_XOR|I_B3|B 0 I3|_XOR|I_B3|MID  PWL(0 0 5e-12 0.000175)
LI3|_XOR|I_Q1|B I3|_XOR|Q1 I3|_XOR|I_Q1|MID  2e-12
II3|_XOR|I_Q1|B 0 I3|_XOR|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_XOR|A1|1 I3|_XOR|A1 I3|_XOR|A1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A1|P I3|_XOR|A1|MID_SERIES 0  5e-13
RI3|_XOR|A1|B I3|_XOR|A1 I3|_XOR|A1|MID_SHUNT  2.7439617672
LI3|_XOR|A1|RB I3|_XOR|A1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A2|1 I3|_XOR|A2 I3|_XOR|A2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A2|P I3|_XOR|A2|MID_SERIES 0  5e-13
RI3|_XOR|A2|B I3|_XOR|A2 I3|_XOR|A2|MID_SHUNT  2.7439617672
LI3|_XOR|A2|RB I3|_XOR|A2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|A3|1 I3|_XOR|A2 I3|_XOR|A3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|A3|P I3|_XOR|A3|MID_SERIES I3|_XOR|A3  1.2e-12
RI3|_XOR|A3|B I3|_XOR|A2 I3|_XOR|A3|MID_SHUNT  2.7439617672
LI3|_XOR|A3|RB I3|_XOR|A3|MID_SHUNT I3|_XOR|A3  2.050338398468e-12
BI3|_XOR|B1|1 I3|_XOR|B1 I3|_XOR|B1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B1|P I3|_XOR|B1|MID_SERIES 0  5e-13
RI3|_XOR|B1|B I3|_XOR|B1 I3|_XOR|B1|MID_SHUNT  2.7439617672
LI3|_XOR|B1|RB I3|_XOR|B1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B2|1 I3|_XOR|B2 I3|_XOR|B2|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B2|P I3|_XOR|B2|MID_SERIES 0  5e-13
RI3|_XOR|B2|B I3|_XOR|B2 I3|_XOR|B2|MID_SHUNT  2.7439617672
LI3|_XOR|B2|RB I3|_XOR|B2|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|B3|1 I3|_XOR|B2 I3|_XOR|B3|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|B3|P I3|_XOR|B3|MID_SERIES I3|_XOR|B3  1.2e-12
RI3|_XOR|B3|B I3|_XOR|B2 I3|_XOR|B3|MID_SHUNT  2.7439617672
LI3|_XOR|B3|RB I3|_XOR|B3|MID_SHUNT I3|_XOR|B3  2.050338398468e-12
BI3|_XOR|T1|1 I3|_XOR|T1 I3|_XOR|T1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|T1|P I3|_XOR|T1|MID_SERIES 0  5e-13
RI3|_XOR|T1|B I3|_XOR|T1 I3|_XOR|T1|MID_SHUNT  2.7439617672
LI3|_XOR|T1|RB I3|_XOR|T1|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|T2|1 I3|_XOR|T2 I3|_XOR|ABTQ JJMIT AREA=2.0
RI3|_XOR|T2|B I3|_XOR|T2 I3|_XOR|T2|MID_SHUNT  3.429952209
LI3|_XOR|T2|RB I3|_XOR|T2|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|AB|1 I3|_XOR|AB I3|_XOR|AB|MID_SERIES JJMIT AREA=2.0
LI3|_XOR|AB|P I3|_XOR|AB|MID_SERIES I3|_XOR|ABTQ  1.2e-12
RI3|_XOR|AB|B I3|_XOR|AB I3|_XOR|AB|MID_SHUNT  3.429952209
LI3|_XOR|AB|RB I3|_XOR|AB|MID_SHUNT I3|_XOR|ABTQ  2.437922998085e-12
BI3|_XOR|ABTQ|1 I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|ABTQ|P I3|_XOR|ABTQ|MID_SERIES 0  5e-13
RI3|_XOR|ABTQ|B I3|_XOR|ABTQ I3|_XOR|ABTQ|MID_SHUNT  2.7439617672
LI3|_XOR|ABTQ|RB I3|_XOR|ABTQ|MID_SHUNT 0  2.050338398468e-12
BI3|_XOR|Q1|1 I3|_XOR|Q1 I3|_XOR|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_XOR|Q1|P I3|_XOR|Q1|MID_SERIES 0  5e-13
RI3|_XOR|Q1|B I3|_XOR|Q1 I3|_XOR|Q1|MID_SHUNT  2.7439617672
LI3|_XOR|Q1|RB I3|_XOR|Q1|MID_SHUNT 0  2.050338398468e-12
LI3|_AND|I_A1|B I3|_AND|A1 I3|_AND|I_A1|MID  2e-12
II3|_AND|I_A1|B 0 I3|_AND|I_A1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_B1|B I3|_AND|B1 I3|_AND|I_B1|MID  2e-12
II3|_AND|I_B1|B 0 I3|_AND|I_B1|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q3|B I3|_AND|Q3 I3|_AND|I_Q3|MID  2e-12
II3|_AND|I_Q3|B 0 I3|_AND|I_Q3|MID  PWL(0 0 5e-12 5e-05)
LI3|_AND|I_Q2|B I3|_AND|Q2 I3|_AND|I_Q2|MID  2e-12
II3|_AND|I_Q2|B 0 I3|_AND|I_Q2|MID  PWL(0 0 5e-12 0.000175)
LI3|_AND|I_Q1|B I3|_AND|Q1 I3|_AND|I_Q1|MID  2e-12
II3|_AND|I_Q1|B 0 I3|_AND|I_Q1|MID  PWL(0 0 5e-12 0.000175)
BI3|_AND|A1|1 I3|_AND|A1 I3|_AND|A1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A1|P I3|_AND|A1|MID_SERIES 0  2e-13
RI3|_AND|A1|B I3|_AND|A1 I3|_AND|A1|MID_SHUNT  2.7439617672
LI3|_AND|A1|RB I3|_AND|A1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A2|1 I3|_AND|A2 I3|_AND|A2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|A2|P I3|_AND|A2|MID_SERIES 0  2e-13
RI3|_AND|A2|B I3|_AND|A2 I3|_AND|A2|MID_SHUNT  2.7439617672
LI3|_AND|A2|RB I3|_AND|A2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|A12|1 I3|_AND|A2 I3|_AND|A3 JJMIT AREA=1.7857142857142858
RI3|_AND|A12|B I3|_AND|A2 I3|_AND|A12|MID_SHUNT  3.84154647408
LI3|_AND|A12|RB I3|_AND|A12|MID_SHUNT I3|_AND|A3  2.1704737578552e-12
BI3|_AND|B1|1 I3|_AND|B1 I3|_AND|B1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B1|P I3|_AND|B1|MID_SERIES 0  2e-13
RI3|_AND|B1|B I3|_AND|B1 I3|_AND|B1|MID_SHUNT  2.7439617672
LI3|_AND|B1|RB I3|_AND|B1|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B2|1 I3|_AND|B2 I3|_AND|B2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|B2|P I3|_AND|B2|MID_SERIES 0  2e-13
RI3|_AND|B2|B I3|_AND|B2 I3|_AND|B2|MID_SHUNT  2.7439617672
LI3|_AND|B2|RB I3|_AND|B2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|B12|1 I3|_AND|B2 I3|_AND|B3 JJMIT AREA=1.7857142857142858
RI3|_AND|B12|B I3|_AND|B2 I3|_AND|B12|MID_SHUNT  3.84154647408
LI3|_AND|B12|RB I3|_AND|B12|MID_SHUNT I3|_AND|B3  2.1704737578552e-12
BI3|_AND|Q2|1 I3|_AND|Q2 I3|_AND|Q2|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q2|P I3|_AND|Q2|MID_SERIES 0  2e-13
RI3|_AND|Q2|B I3|_AND|Q2 I3|_AND|Q2|MID_SHUNT  2.7439617672
LI3|_AND|Q2|RB I3|_AND|Q2|MID_SHUNT 0  1.550338398468e-12
BI3|_AND|Q1|1 I3|_AND|Q1 I3|_AND|Q1|MID_SERIES JJMIT AREA=2.5
LI3|_AND|Q1|P I3|_AND|Q1|MID_SERIES 0  2e-13
RI3|_AND|Q1|B I3|_AND|Q1 I3|_AND|Q1|MID_SHUNT  2.7439617672
LI3|_AND|Q1|RB I3|_AND|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL1|I_D1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|I_D1|MID  2e-12
ISPL_IP2_0|SPL1|I_D1|B 0 SPL_IP2_0|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL1|I_D2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|I_D2|MID  2e-12
ISPL_IP2_0|SPL1|I_D2|B 0 SPL_IP2_0|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_IP2_0|SPL1|I_Q1|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|I_Q1|MID  2e-12
ISPL_IP2_0|SPL1|I_Q1|B 0 SPL_IP2_0|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL1|I_Q2|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|I_Q2|MID  2e-12
ISPL_IP2_0|SPL1|I_Q2|B 0 SPL_IP2_0|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_IP2_0|SPL1|1|1 SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|1|P SPL_IP2_0|SPL1|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|1|B SPL_IP2_0|SPL1|D1 SPL_IP2_0|SPL1|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|1|RB SPL_IP2_0|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|2|1 SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|2|P SPL_IP2_0|SPL1|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|2|B SPL_IP2_0|SPL1|D2 SPL_IP2_0|SPL1|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|2|RB SPL_IP2_0|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|A|1 SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|A|P SPL_IP2_0|SPL1|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|A|B SPL_IP2_0|SPL1|QA1 SPL_IP2_0|SPL1|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|A|RB SPL_IP2_0|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL1|B|1 SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL1|B|P SPL_IP2_0|SPL1|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL1|B|B SPL_IP2_0|SPL1|QB1 SPL_IP2_0|SPL1|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL1|B|RB SPL_IP2_0|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_IP2_0|SPL2|I_D1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|I_D1|MID  2e-12
ISPL_IP2_0|SPL2|I_D1|B 0 SPL_IP2_0|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL2|I_D2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|I_D2|MID  2e-12
ISPL_IP2_0|SPL2|I_D2|B 0 SPL_IP2_0|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_IP2_0|SPL2|I_Q1|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|I_Q1|MID  2e-12
ISPL_IP2_0|SPL2|I_Q1|B 0 SPL_IP2_0|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_IP2_0|SPL2|I_Q2|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|I_Q2|MID  2e-12
ISPL_IP2_0|SPL2|I_Q2|B 0 SPL_IP2_0|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_IP2_0|SPL2|1|1 SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|1|P SPL_IP2_0|SPL2|1|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|1|B SPL_IP2_0|SPL2|D1 SPL_IP2_0|SPL2|1|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|1|RB SPL_IP2_0|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|2|1 SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|2|P SPL_IP2_0|SPL2|2|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|2|B SPL_IP2_0|SPL2|D2 SPL_IP2_0|SPL2|2|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|2|RB SPL_IP2_0|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|A|1 SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|A|P SPL_IP2_0|SPL2|A|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|A|B SPL_IP2_0|SPL2|QA1 SPL_IP2_0|SPL2|A|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|A|RB SPL_IP2_0|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_IP2_0|SPL2|B|1 SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_IP2_0|SPL2|B|P SPL_IP2_0|SPL2|B|MID_SERIES 0  2e-13
RSPL_IP2_0|SPL2|B|B SPL_IP2_0|SPL2|QB1 SPL_IP2_0|SPL2|B|MID_SHUNT  2.7439617672
LSPL_IP2_0|SPL2|B|RB SPL_IP2_0|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|P|I_1|B _PG0_01|P|A1 _PG0_01|P|I_1|MID  2e-12
I_PG0_01|P|I_1|B 0 _PG0_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_3|B _PG0_01|P|A3 _PG0_01|P|I_3|MID  2e-12
I_PG0_01|P|I_3|B 0 _PG0_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|P|I_T|B _PG0_01|P|T1 _PG0_01|P|I_T|MID  2e-12
I_PG0_01|P|I_T|B 0 _PG0_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|P|I_6|B _PG0_01|P|Q1 _PG0_01|P|I_6|MID  2e-12
I_PG0_01|P|I_6|B 0 _PG0_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|P|1|1 _PG0_01|P|A1 _PG0_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|1|P _PG0_01|P|1|MID_SERIES 0  2e-13
R_PG0_01|P|1|B _PG0_01|P|A1 _PG0_01|P|1|MID_SHUNT  2.7439617672
L_PG0_01|P|1|RB _PG0_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|23|1 _PG0_01|P|A2 _PG0_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|P|23|B _PG0_01|P|A2 _PG0_01|P|23|MID_SHUNT  3.84154647408
L_PG0_01|P|23|RB _PG0_01|P|23|MID_SHUNT _PG0_01|P|A3  2.1704737578552e-12
B_PG0_01|P|3|1 _PG0_01|P|A3 _PG0_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|3|P _PG0_01|P|3|MID_SERIES 0  2e-13
R_PG0_01|P|3|B _PG0_01|P|A3 _PG0_01|P|3|MID_SHUNT  2.7439617672
L_PG0_01|P|3|RB _PG0_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|4|1 _PG0_01|P|A4 _PG0_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|4|P _PG0_01|P|4|MID_SERIES 0  2e-13
R_PG0_01|P|4|B _PG0_01|P|A4 _PG0_01|P|4|MID_SHUNT  2.7439617672
L_PG0_01|P|4|RB _PG0_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|T|1 _PG0_01|P|T1 _PG0_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|T|P _PG0_01|P|T|MID_SERIES 0  2e-13
R_PG0_01|P|T|B _PG0_01|P|T1 _PG0_01|P|T|MID_SHUNT  2.7439617672
L_PG0_01|P|T|RB _PG0_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|P|45|1 _PG0_01|P|T2 _PG0_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|P|45|B _PG0_01|P|T2 _PG0_01|P|45|MID_SHUNT  3.84154647408
L_PG0_01|P|45|RB _PG0_01|P|45|MID_SHUNT _PG0_01|P|A4  2.1704737578552e-12
B_PG0_01|P|6|1 _PG0_01|P|Q1 _PG0_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|P|6|P _PG0_01|P|6|MID_SERIES 0  2e-13
R_PG0_01|P|6|B _PG0_01|P|Q1 _PG0_01|P|6|MID_SHUNT  2.7439617672
L_PG0_01|P|6|RB _PG0_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_01|G|I_1|B _PG0_01|G|A1 _PG0_01|G|I_1|MID  2e-12
I_PG0_01|G|I_1|B 0 _PG0_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_3|B _PG0_01|G|A3 _PG0_01|G|I_3|MID  2e-12
I_PG0_01|G|I_3|B 0 _PG0_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_01|G|I_T|B _PG0_01|G|T1 _PG0_01|G|I_T|MID  2e-12
I_PG0_01|G|I_T|B 0 _PG0_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_01|G|I_6|B _PG0_01|G|Q1 _PG0_01|G|I_6|MID  2e-12
I_PG0_01|G|I_6|B 0 _PG0_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_01|G|1|1 _PG0_01|G|A1 _PG0_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|1|P _PG0_01|G|1|MID_SERIES 0  2e-13
R_PG0_01|G|1|B _PG0_01|G|A1 _PG0_01|G|1|MID_SHUNT  2.7439617672
L_PG0_01|G|1|RB _PG0_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|23|1 _PG0_01|G|A2 _PG0_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_01|G|23|B _PG0_01|G|A2 _PG0_01|G|23|MID_SHUNT  3.84154647408
L_PG0_01|G|23|RB _PG0_01|G|23|MID_SHUNT _PG0_01|G|A3  2.1704737578552e-12
B_PG0_01|G|3|1 _PG0_01|G|A3 _PG0_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|3|P _PG0_01|G|3|MID_SERIES 0  2e-13
R_PG0_01|G|3|B _PG0_01|G|A3 _PG0_01|G|3|MID_SHUNT  2.7439617672
L_PG0_01|G|3|RB _PG0_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|4|1 _PG0_01|G|A4 _PG0_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|4|P _PG0_01|G|4|MID_SERIES 0  2e-13
R_PG0_01|G|4|B _PG0_01|G|A4 _PG0_01|G|4|MID_SHUNT  2.7439617672
L_PG0_01|G|4|RB _PG0_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|T|1 _PG0_01|G|T1 _PG0_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|T|P _PG0_01|G|T|MID_SERIES 0  2e-13
R_PG0_01|G|T|B _PG0_01|G|T1 _PG0_01|G|T|MID_SHUNT  2.7439617672
L_PG0_01|G|T|RB _PG0_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_01|G|45|1 _PG0_01|G|T2 _PG0_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_01|G|45|B _PG0_01|G|T2 _PG0_01|G|45|MID_SHUNT  3.84154647408
L_PG0_01|G|45|RB _PG0_01|G|45|MID_SHUNT _PG0_01|G|A4  2.1704737578552e-12
B_PG0_01|G|6|1 _PG0_01|G|Q1 _PG0_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_01|G|6|P _PG0_01|G|6|MID_SERIES 0  2e-13
R_PG0_01|G|6|B _PG0_01|G|Q1 _PG0_01|G|6|MID_SHUNT  2.7439617672
L_PG0_01|G|6|RB _PG0_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_SPL_G1|I_D1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|I_D1|MID  2e-12
I_PG1_01|_SPL_G1|I_D1|B 0 _PG1_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_D2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|I_D2|MID  2e-12
I_PG1_01|_SPL_G1|I_D2|B 0 _PG1_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG1_01|_SPL_G1|I_Q1|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|I_Q1|MID  2e-12
I_PG1_01|_SPL_G1|I_Q1|B 0 _PG1_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG1_01|_SPL_G1|I_Q2|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|I_Q2|MID  2e-12
I_PG1_01|_SPL_G1|I_Q2|B 0 _PG1_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG1_01|_SPL_G1|1|1 _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|1|P _PG1_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|1|B _PG1_01|_SPL_G1|D1 _PG1_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|1|RB _PG1_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|2|1 _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|2|P _PG1_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|2|B _PG1_01|_SPL_G1|D2 _PG1_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|2|RB _PG1_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|A|1 _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|A|P _PG1_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|A|B _PG1_01|_SPL_G1|QA1 _PG1_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|A|RB _PG1_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_SPL_G1|B|1 _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_SPL_G1|B|P _PG1_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG1_01|_SPL_G1|B|B _PG1_01|_SPL_G1|QB1 _PG1_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG1_01|_SPL_G1|B|RB _PG1_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_PG|I_A1|B _PG1_01|_PG|A1 _PG1_01|_PG|I_A1|MID  2e-12
I_PG1_01|_PG|I_A1|B 0 _PG1_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_B1|B _PG1_01|_PG|B1 _PG1_01|_PG|I_B1|MID  2e-12
I_PG1_01|_PG|I_B1|B 0 _PG1_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q3|B _PG1_01|_PG|Q3 _PG1_01|_PG|I_Q3|MID  2e-12
I_PG1_01|_PG|I_Q3|B 0 _PG1_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_PG|I_Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|I_Q2|MID  2e-12
I_PG1_01|_PG|I_Q2|B 0 _PG1_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_PG|I_Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|I_Q1|MID  2e-12
I_PG1_01|_PG|I_Q1|B 0 _PG1_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_PG|A1|1 _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A1|P _PG1_01|_PG|A1|MID_SERIES 0  2e-13
R_PG1_01|_PG|A1|B _PG1_01|_PG|A1 _PG1_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A1|RB _PG1_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A2|1 _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|A2|P _PG1_01|_PG|A2|MID_SERIES 0  2e-13
R_PG1_01|_PG|A2|B _PG1_01|_PG|A2 _PG1_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|A2|RB _PG1_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|A12|1 _PG1_01|_PG|A2 _PG1_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|A12|B _PG1_01|_PG|A2 _PG1_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|A12|RB _PG1_01|_PG|A12|MID_SHUNT _PG1_01|_PG|A3  2.1704737578552e-12
B_PG1_01|_PG|B1|1 _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B1|P _PG1_01|_PG|B1|MID_SERIES 0  2e-13
R_PG1_01|_PG|B1|B _PG1_01|_PG|B1 _PG1_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B1|RB _PG1_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B2|1 _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|B2|P _PG1_01|_PG|B2|MID_SERIES 0  2e-13
R_PG1_01|_PG|B2|B _PG1_01|_PG|B2 _PG1_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|B2|RB _PG1_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|B12|1 _PG1_01|_PG|B2 _PG1_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_PG|B12|B _PG1_01|_PG|B2 _PG1_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_PG|B12|RB _PG1_01|_PG|B12|MID_SHUNT _PG1_01|_PG|B3  2.1704737578552e-12
B_PG1_01|_PG|Q2|1 _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q2|P _PG1_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q2|B _PG1_01|_PG|Q2 _PG1_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q2|RB _PG1_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_PG|Q1|1 _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_PG|Q1|P _PG1_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_PG|Q1|B _PG1_01|_PG|Q1 _PG1_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_PG|Q1|RB _PG1_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_GG|I_A1|B _PG1_01|_GG|A1 _PG1_01|_GG|I_A1|MID  2e-12
I_PG1_01|_GG|I_A1|B 0 _PG1_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_B1|B _PG1_01|_GG|B1 _PG1_01|_GG|I_B1|MID  2e-12
I_PG1_01|_GG|I_B1|B 0 _PG1_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q3|B _PG1_01|_GG|Q3 _PG1_01|_GG|I_Q3|MID  2e-12
I_PG1_01|_GG|I_Q3|B 0 _PG1_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_GG|I_Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|I_Q2|MID  2e-12
I_PG1_01|_GG|I_Q2|B 0 _PG1_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_GG|I_Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|I_Q1|MID  2e-12
I_PG1_01|_GG|I_Q1|B 0 _PG1_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_GG|A1|1 _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A1|P _PG1_01|_GG|A1|MID_SERIES 0  2e-13
R_PG1_01|_GG|A1|B _PG1_01|_GG|A1 _PG1_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A1|RB _PG1_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A2|1 _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|A2|P _PG1_01|_GG|A2|MID_SERIES 0  2e-13
R_PG1_01|_GG|A2|B _PG1_01|_GG|A2 _PG1_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|A2|RB _PG1_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|A12|1 _PG1_01|_GG|A2 _PG1_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|A12|B _PG1_01|_GG|A2 _PG1_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|A12|RB _PG1_01|_GG|A12|MID_SHUNT _PG1_01|_GG|A3  2.1704737578552e-12
B_PG1_01|_GG|B1|1 _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B1|P _PG1_01|_GG|B1|MID_SERIES 0  2e-13
R_PG1_01|_GG|B1|B _PG1_01|_GG|B1 _PG1_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B1|RB _PG1_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B2|1 _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|B2|P _PG1_01|_GG|B2|MID_SERIES 0  2e-13
R_PG1_01|_GG|B2|B _PG1_01|_GG|B2 _PG1_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|B2|RB _PG1_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|B12|1 _PG1_01|_GG|B2 _PG1_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_GG|B12|B _PG1_01|_GG|B2 _PG1_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG1_01|_GG|B12|RB _PG1_01|_GG|B12|MID_SHUNT _PG1_01|_GG|B3  2.1704737578552e-12
B_PG1_01|_GG|Q2|1 _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q2|P _PG1_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q2|B _PG1_01|_GG|Q2 _PG1_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q2|RB _PG1_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_GG|Q1|1 _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_GG|Q1|P _PG1_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG1_01|_GG|Q1|B _PG1_01|_GG|Q1 _PG1_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_GG|Q1|RB _PG1_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_PG|I_1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|I_1|MID  2e-12
I_PG1_01|_DFF_PG|I_1|B 0 _PG1_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|I_3|MID  2e-12
I_PG1_01|_DFF_PG|I_3|B 0 _PG1_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_PG|I_T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|I_T|MID  2e-12
I_PG1_01|_DFF_PG|I_T|B 0 _PG1_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_PG|I_6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|I_6|MID  2e-12
I_PG1_01|_DFF_PG|I_6|B 0 _PG1_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_PG|1|1 _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|1|P _PG1_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|1|B _PG1_01|_DFF_PG|A1 _PG1_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|1|RB _PG1_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|23|1 _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|23|B _PG1_01|_DFF_PG|A2 _PG1_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|23|RB _PG1_01|_DFF_PG|23|MID_SHUNT _PG1_01|_DFF_PG|A3  2.1704737578552e-12
B_PG1_01|_DFF_PG|3|1 _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|3|P _PG1_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|3|B _PG1_01|_DFF_PG|A3 _PG1_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|3|RB _PG1_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|4|1 _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|4|P _PG1_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|4|B _PG1_01|_DFF_PG|A4 _PG1_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|4|RB _PG1_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|T|1 _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|T|P _PG1_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|T|B _PG1_01|_DFF_PG|T1 _PG1_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|T|RB _PG1_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_PG|45|1 _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_PG|45|B _PG1_01|_DFF_PG|T2 _PG1_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_PG|45|RB _PG1_01|_DFF_PG|45|MID_SHUNT _PG1_01|_DFF_PG|A4  2.1704737578552e-12
B_PG1_01|_DFF_PG|6|1 _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_PG|6|P _PG1_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_PG|6|B _PG1_01|_DFF_PG|Q1 _PG1_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_PG|6|RB _PG1_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_DFF_GG|I_1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|I_1|MID  2e-12
I_PG1_01|_DFF_GG|I_1|B 0 _PG1_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|I_3|MID  2e-12
I_PG1_01|_DFF_GG|I_3|B 0 _PG1_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG1_01|_DFF_GG|I_T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|I_T|MID  2e-12
I_PG1_01|_DFF_GG|I_T|B 0 _PG1_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_DFF_GG|I_6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|I_6|MID  2e-12
I_PG1_01|_DFF_GG|I_6|B 0 _PG1_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_DFF_GG|1|1 _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|1|P _PG1_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|1|B _PG1_01|_DFF_GG|A1 _PG1_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|1|RB _PG1_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|23|1 _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|23|B _PG1_01|_DFF_GG|A2 _PG1_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|23|RB _PG1_01|_DFF_GG|23|MID_SHUNT _PG1_01|_DFF_GG|A3  2.1704737578552e-12
B_PG1_01|_DFF_GG|3|1 _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|3|P _PG1_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|3|B _PG1_01|_DFF_GG|A3 _PG1_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|3|RB _PG1_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|4|1 _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|4|P _PG1_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|4|B _PG1_01|_DFF_GG|A4 _PG1_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|4|RB _PG1_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|T|1 _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|T|P _PG1_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|T|B _PG1_01|_DFF_GG|T1 _PG1_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|T|RB _PG1_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_DFF_GG|45|1 _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG1_01|_DFF_GG|45|B _PG1_01|_DFF_GG|T2 _PG1_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG1_01|_DFF_GG|45|RB _PG1_01|_DFF_GG|45|MID_SHUNT _PG1_01|_DFF_GG|A4  2.1704737578552e-12
B_PG1_01|_DFF_GG|6|1 _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_DFF_GG|6|P _PG1_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG1_01|_DFF_GG|6|B _PG1_01|_DFF_GG|Q1 _PG1_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG1_01|_DFF_GG|6|RB _PG1_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG1_01|_AND_G|I_A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|I_A1|MID  2e-12
I_PG1_01|_AND_G|I_A1|B 0 _PG1_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|I_B1|MID  2e-12
I_PG1_01|_AND_G|I_B1|B 0 _PG1_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q3|B _PG1_01|_AND_G|Q3 _PG1_01|_AND_G|I_Q3|MID  2e-12
I_PG1_01|_AND_G|I_Q3|B 0 _PG1_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG1_01|_AND_G|I_Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|I_Q2|MID  2e-12
I_PG1_01|_AND_G|I_Q2|B 0 _PG1_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG1_01|_AND_G|I_Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|I_Q1|MID  2e-12
I_PG1_01|_AND_G|I_Q1|B 0 _PG1_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG1_01|_AND_G|A1|1 _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A1|P _PG1_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A1|B _PG1_01|_AND_G|A1 _PG1_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A1|RB _PG1_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A2|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|A2|P _PG1_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|A2|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|A2|RB _PG1_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|A12|1 _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|A12|B _PG1_01|_AND_G|A2 _PG1_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|A12|RB _PG1_01|_AND_G|A12|MID_SHUNT _PG1_01|_AND_G|A3  2.1704737578552e-12
B_PG1_01|_AND_G|B1|1 _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B1|P _PG1_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B1|B _PG1_01|_AND_G|B1 _PG1_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B1|RB _PG1_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B2|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|B2|P _PG1_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|B2|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|B2|RB _PG1_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|B12|1 _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG1_01|_AND_G|B12|B _PG1_01|_AND_G|B2 _PG1_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG1_01|_AND_G|B12|RB _PG1_01|_AND_G|B12|MID_SHUNT _PG1_01|_AND_G|B3  2.1704737578552e-12
B_PG1_01|_AND_G|Q2|1 _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q2|P _PG1_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q2|B _PG1_01|_AND_G|Q2 _PG1_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q2|RB _PG1_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG1_01|_AND_G|Q1|1 _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG1_01|_AND_G|Q1|P _PG1_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG1_01|_AND_G|Q1|B _PG1_01|_AND_G|Q1 _PG1_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG1_01|_AND_G|Q1|RB _PG1_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|P|I_1|B _PG2_01|P|A1 _PG2_01|P|I_1|MID  2e-12
I_PG2_01|P|I_1|B 0 _PG2_01|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_3|B _PG2_01|P|A3 _PG2_01|P|I_3|MID  2e-12
I_PG2_01|P|I_3|B 0 _PG2_01|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|P|I_T|B _PG2_01|P|T1 _PG2_01|P|I_T|MID  2e-12
I_PG2_01|P|I_T|B 0 _PG2_01|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|P|I_6|B _PG2_01|P|Q1 _PG2_01|P|I_6|MID  2e-12
I_PG2_01|P|I_6|B 0 _PG2_01|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|P|1|1 _PG2_01|P|A1 _PG2_01|P|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|1|P _PG2_01|P|1|MID_SERIES 0  2e-13
R_PG2_01|P|1|B _PG2_01|P|A1 _PG2_01|P|1|MID_SHUNT  2.7439617672
L_PG2_01|P|1|RB _PG2_01|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|23|1 _PG2_01|P|A2 _PG2_01|P|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|P|23|B _PG2_01|P|A2 _PG2_01|P|23|MID_SHUNT  3.84154647408
L_PG2_01|P|23|RB _PG2_01|P|23|MID_SHUNT _PG2_01|P|A3  2.1704737578552e-12
B_PG2_01|P|3|1 _PG2_01|P|A3 _PG2_01|P|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|3|P _PG2_01|P|3|MID_SERIES 0  2e-13
R_PG2_01|P|3|B _PG2_01|P|A3 _PG2_01|P|3|MID_SHUNT  2.7439617672
L_PG2_01|P|3|RB _PG2_01|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|4|1 _PG2_01|P|A4 _PG2_01|P|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|4|P _PG2_01|P|4|MID_SERIES 0  2e-13
R_PG2_01|P|4|B _PG2_01|P|A4 _PG2_01|P|4|MID_SHUNT  2.7439617672
L_PG2_01|P|4|RB _PG2_01|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|T|1 _PG2_01|P|T1 _PG2_01|P|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|T|P _PG2_01|P|T|MID_SERIES 0  2e-13
R_PG2_01|P|T|B _PG2_01|P|T1 _PG2_01|P|T|MID_SHUNT  2.7439617672
L_PG2_01|P|T|RB _PG2_01|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|P|45|1 _PG2_01|P|T2 _PG2_01|P|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|P|45|B _PG2_01|P|T2 _PG2_01|P|45|MID_SHUNT  3.84154647408
L_PG2_01|P|45|RB _PG2_01|P|45|MID_SHUNT _PG2_01|P|A4  2.1704737578552e-12
B_PG2_01|P|6|1 _PG2_01|P|Q1 _PG2_01|P|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|P|6|P _PG2_01|P|6|MID_SERIES 0  2e-13
R_PG2_01|P|6|B _PG2_01|P|Q1 _PG2_01|P|6|MID_SHUNT  2.7439617672
L_PG2_01|P|6|RB _PG2_01|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_01|G|I_1|B _PG2_01|G|A1 _PG2_01|G|I_1|MID  2e-12
I_PG2_01|G|I_1|B 0 _PG2_01|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_3|B _PG2_01|G|A3 _PG2_01|G|I_3|MID  2e-12
I_PG2_01|G|I_3|B 0 _PG2_01|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_01|G|I_T|B _PG2_01|G|T1 _PG2_01|G|I_T|MID  2e-12
I_PG2_01|G|I_T|B 0 _PG2_01|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_01|G|I_6|B _PG2_01|G|Q1 _PG2_01|G|I_6|MID  2e-12
I_PG2_01|G|I_6|B 0 _PG2_01|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_01|G|1|1 _PG2_01|G|A1 _PG2_01|G|1|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|1|P _PG2_01|G|1|MID_SERIES 0  2e-13
R_PG2_01|G|1|B _PG2_01|G|A1 _PG2_01|G|1|MID_SHUNT  2.7439617672
L_PG2_01|G|1|RB _PG2_01|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|23|1 _PG2_01|G|A2 _PG2_01|G|A3 JJMIT AREA=1.7857142857142858
R_PG2_01|G|23|B _PG2_01|G|A2 _PG2_01|G|23|MID_SHUNT  3.84154647408
L_PG2_01|G|23|RB _PG2_01|G|23|MID_SHUNT _PG2_01|G|A3  2.1704737578552e-12
B_PG2_01|G|3|1 _PG2_01|G|A3 _PG2_01|G|3|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|3|P _PG2_01|G|3|MID_SERIES 0  2e-13
R_PG2_01|G|3|B _PG2_01|G|A3 _PG2_01|G|3|MID_SHUNT  2.7439617672
L_PG2_01|G|3|RB _PG2_01|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|4|1 _PG2_01|G|A4 _PG2_01|G|4|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|4|P _PG2_01|G|4|MID_SERIES 0  2e-13
R_PG2_01|G|4|B _PG2_01|G|A4 _PG2_01|G|4|MID_SHUNT  2.7439617672
L_PG2_01|G|4|RB _PG2_01|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|T|1 _PG2_01|G|T1 _PG2_01|G|T|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|T|P _PG2_01|G|T|MID_SERIES 0  2e-13
R_PG2_01|G|T|B _PG2_01|G|T1 _PG2_01|G|T|MID_SHUNT  2.7439617672
L_PG2_01|G|T|RB _PG2_01|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_01|G|45|1 _PG2_01|G|T2 _PG2_01|G|A4 JJMIT AREA=1.7857142857142858
R_PG2_01|G|45|B _PG2_01|G|T2 _PG2_01|G|45|MID_SHUNT  3.84154647408
L_PG2_01|G|45|RB _PG2_01|G|45|MID_SHUNT _PG2_01|G|A4  2.1704737578552e-12
B_PG2_01|G|6|1 _PG2_01|G|Q1 _PG2_01|G|6|MID_SERIES JJMIT AREA=2.5
L_PG2_01|G|6|P _PG2_01|G|6|MID_SERIES 0  2e-13
R_PG2_01|G|6|B _PG2_01|G|Q1 _PG2_01|G|6|MID_SHUNT  2.7439617672
L_PG2_01|G|6|RB _PG2_01|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_G1|I_D1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|I_D1|MID  2e-12
I_PG3_01|_SPL_G1|I_D1|B 0 _PG3_01|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_D2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|I_D2|MID  2e-12
I_PG3_01|_SPL_G1|I_D2|B 0 _PG3_01|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_G1|I_Q1|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|I_Q1|MID  2e-12
I_PG3_01|_SPL_G1|I_Q1|B 0 _PG3_01|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_G1|I_Q2|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|I_Q2|MID  2e-12
I_PG3_01|_SPL_G1|I_Q2|B 0 _PG3_01|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_G1|1|1 _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|1|P _PG3_01|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|1|B _PG3_01|_SPL_G1|D1 _PG3_01|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|1|RB _PG3_01|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|2|1 _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|2|P _PG3_01|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|2|B _PG3_01|_SPL_G1|D2 _PG3_01|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|2|RB _PG3_01|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|A|1 _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|A|P _PG3_01|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|A|B _PG3_01|_SPL_G1|QA1 _PG3_01|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|A|RB _PG3_01|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_G1|B|1 _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_G1|B|P _PG3_01|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_G1|B|B _PG3_01|_SPL_G1|QB1 _PG3_01|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_G1|B|RB _PG3_01|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_SPL_P1|I_D1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|I_D1|MID  2e-12
I_PG3_01|_SPL_P1|I_D1|B 0 _PG3_01|_SPL_P1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_D2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|I_D2|MID  2e-12
I_PG3_01|_SPL_P1|I_D2|B 0 _PG3_01|_SPL_P1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_01|_SPL_P1|I_Q1|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|I_Q1|MID  2e-12
I_PG3_01|_SPL_P1|I_Q1|B 0 _PG3_01|_SPL_P1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_01|_SPL_P1|I_Q2|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|I_Q2|MID  2e-12
I_PG3_01|_SPL_P1|I_Q2|B 0 _PG3_01|_SPL_P1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_01|_SPL_P1|1|1 _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|1|P _PG3_01|_SPL_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|1|B _PG3_01|_SPL_P1|D1 _PG3_01|_SPL_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|1|RB _PG3_01|_SPL_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|2|1 _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|2|P _PG3_01|_SPL_P1|2|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|2|B _PG3_01|_SPL_P1|D2 _PG3_01|_SPL_P1|2|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|2|RB _PG3_01|_SPL_P1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|A|1 _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|A|P _PG3_01|_SPL_P1|A|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|A|B _PG3_01|_SPL_P1|QA1 _PG3_01|_SPL_P1|A|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|A|RB _PG3_01|_SPL_P1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_SPL_P1|B|1 _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_SPL_P1|B|P _PG3_01|_SPL_P1|B|MID_SERIES 0  2e-13
R_PG3_01|_SPL_P1|B|B _PG3_01|_SPL_P1|QB1 _PG3_01|_SPL_P1|B|MID_SHUNT  2.7439617672
L_PG3_01|_SPL_P1|B|RB _PG3_01|_SPL_P1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_PG|I_A1|B _PG3_01|_PG|A1 _PG3_01|_PG|I_A1|MID  2e-12
I_PG3_01|_PG|I_A1|B 0 _PG3_01|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_B1|B _PG3_01|_PG|B1 _PG3_01|_PG|I_B1|MID  2e-12
I_PG3_01|_PG|I_B1|B 0 _PG3_01|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q3|B _PG3_01|_PG|Q3 _PG3_01|_PG|I_Q3|MID  2e-12
I_PG3_01|_PG|I_Q3|B 0 _PG3_01|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_PG|I_Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|I_Q2|MID  2e-12
I_PG3_01|_PG|I_Q2|B 0 _PG3_01|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_PG|I_Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|I_Q1|MID  2e-12
I_PG3_01|_PG|I_Q1|B 0 _PG3_01|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_PG|A1|1 _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A1|P _PG3_01|_PG|A1|MID_SERIES 0  2e-13
R_PG3_01|_PG|A1|B _PG3_01|_PG|A1 _PG3_01|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A1|RB _PG3_01|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A2|1 _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|A2|P _PG3_01|_PG|A2|MID_SERIES 0  2e-13
R_PG3_01|_PG|A2|B _PG3_01|_PG|A2 _PG3_01|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|A2|RB _PG3_01|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|A12|1 _PG3_01|_PG|A2 _PG3_01|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|A12|B _PG3_01|_PG|A2 _PG3_01|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|A12|RB _PG3_01|_PG|A12|MID_SHUNT _PG3_01|_PG|A3  2.1704737578552e-12
B_PG3_01|_PG|B1|1 _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B1|P _PG3_01|_PG|B1|MID_SERIES 0  2e-13
R_PG3_01|_PG|B1|B _PG3_01|_PG|B1 _PG3_01|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B1|RB _PG3_01|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B2|1 _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|B2|P _PG3_01|_PG|B2|MID_SERIES 0  2e-13
R_PG3_01|_PG|B2|B _PG3_01|_PG|B2 _PG3_01|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|B2|RB _PG3_01|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|B12|1 _PG3_01|_PG|B2 _PG3_01|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_PG|B12|B _PG3_01|_PG|B2 _PG3_01|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_PG|B12|RB _PG3_01|_PG|B12|MID_SHUNT _PG3_01|_PG|B3  2.1704737578552e-12
B_PG3_01|_PG|Q2|1 _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q2|P _PG3_01|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q2|B _PG3_01|_PG|Q2 _PG3_01|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q2|RB _PG3_01|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_PG|Q1|1 _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_PG|Q1|P _PG3_01|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_PG|Q1|B _PG3_01|_PG|Q1 _PG3_01|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_PG|Q1|RB _PG3_01|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_GG|I_A1|B _PG3_01|_GG|A1 _PG3_01|_GG|I_A1|MID  2e-12
I_PG3_01|_GG|I_A1|B 0 _PG3_01|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_B1|B _PG3_01|_GG|B1 _PG3_01|_GG|I_B1|MID  2e-12
I_PG3_01|_GG|I_B1|B 0 _PG3_01|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q3|B _PG3_01|_GG|Q3 _PG3_01|_GG|I_Q3|MID  2e-12
I_PG3_01|_GG|I_Q3|B 0 _PG3_01|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_GG|I_Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|I_Q2|MID  2e-12
I_PG3_01|_GG|I_Q2|B 0 _PG3_01|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_GG|I_Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|I_Q1|MID  2e-12
I_PG3_01|_GG|I_Q1|B 0 _PG3_01|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_GG|A1|1 _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A1|P _PG3_01|_GG|A1|MID_SERIES 0  2e-13
R_PG3_01|_GG|A1|B _PG3_01|_GG|A1 _PG3_01|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A1|RB _PG3_01|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A2|1 _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|A2|P _PG3_01|_GG|A2|MID_SERIES 0  2e-13
R_PG3_01|_GG|A2|B _PG3_01|_GG|A2 _PG3_01|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|A2|RB _PG3_01|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|A12|1 _PG3_01|_GG|A2 _PG3_01|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|A12|B _PG3_01|_GG|A2 _PG3_01|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|A12|RB _PG3_01|_GG|A12|MID_SHUNT _PG3_01|_GG|A3  2.1704737578552e-12
B_PG3_01|_GG|B1|1 _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B1|P _PG3_01|_GG|B1|MID_SERIES 0  2e-13
R_PG3_01|_GG|B1|B _PG3_01|_GG|B1 _PG3_01|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B1|RB _PG3_01|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B2|1 _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|B2|P _PG3_01|_GG|B2|MID_SERIES 0  2e-13
R_PG3_01|_GG|B2|B _PG3_01|_GG|B2 _PG3_01|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|B2|RB _PG3_01|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|B12|1 _PG3_01|_GG|B2 _PG3_01|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_GG|B12|B _PG3_01|_GG|B2 _PG3_01|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_01|_GG|B12|RB _PG3_01|_GG|B12|MID_SHUNT _PG3_01|_GG|B3  2.1704737578552e-12
B_PG3_01|_GG|Q2|1 _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q2|P _PG3_01|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q2|B _PG3_01|_GG|Q2 _PG3_01|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q2|RB _PG3_01|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_GG|Q1|1 _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_GG|Q1|P _PG3_01|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_01|_GG|Q1|B _PG3_01|_GG|Q1 _PG3_01|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_GG|Q1|RB _PG3_01|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P0|I_1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|I_1|MID  2e-12
I_PG3_01|_DFF_P0|I_1|B 0 _PG3_01|_DFF_P0|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|I_3|MID  2e-12
I_PG3_01|_DFF_P0|I_3|B 0 _PG3_01|_DFF_P0|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P0|I_T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|I_T|MID  2e-12
I_PG3_01|_DFF_P0|I_T|B 0 _PG3_01|_DFF_P0|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P0|I_6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|I_6|MID  2e-12
I_PG3_01|_DFF_P0|I_6|B 0 _PG3_01|_DFF_P0|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P0|1|1 _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|1|P _PG3_01|_DFF_P0|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|1|B _PG3_01|_DFF_P0|A1 _PG3_01|_DFF_P0|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|1|RB _PG3_01|_DFF_P0|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|23|1 _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|23|B _PG3_01|_DFF_P0|A2 _PG3_01|_DFF_P0|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|23|RB _PG3_01|_DFF_P0|23|MID_SHUNT _PG3_01|_DFF_P0|A3  2.1704737578552e-12
B_PG3_01|_DFF_P0|3|1 _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|3|P _PG3_01|_DFF_P0|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|3|B _PG3_01|_DFF_P0|A3 _PG3_01|_DFF_P0|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|3|RB _PG3_01|_DFF_P0|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|4|1 _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|4|P _PG3_01|_DFF_P0|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|4|B _PG3_01|_DFF_P0|A4 _PG3_01|_DFF_P0|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|4|RB _PG3_01|_DFF_P0|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|T|1 _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|T|P _PG3_01|_DFF_P0|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|T|B _PG3_01|_DFF_P0|T1 _PG3_01|_DFF_P0|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|T|RB _PG3_01|_DFF_P0|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P0|45|1 _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P0|45|B _PG3_01|_DFF_P0|T2 _PG3_01|_DFF_P0|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P0|45|RB _PG3_01|_DFF_P0|45|MID_SHUNT _PG3_01|_DFF_P0|A4  2.1704737578552e-12
B_PG3_01|_DFF_P0|6|1 _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P0|6|P _PG3_01|_DFF_P0|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P0|6|B _PG3_01|_DFF_P0|Q1 _PG3_01|_DFF_P0|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P0|6|RB _PG3_01|_DFF_P0|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_P1|I_1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|I_1|MID  2e-12
I_PG3_01|_DFF_P1|I_1|B 0 _PG3_01|_DFF_P1|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|I_3|MID  2e-12
I_PG3_01|_DFF_P1|I_3|B 0 _PG3_01|_DFF_P1|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_P1|I_T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|I_T|MID  2e-12
I_PG3_01|_DFF_P1|I_T|B 0 _PG3_01|_DFF_P1|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_P1|I_6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|I_6|MID  2e-12
I_PG3_01|_DFF_P1|I_6|B 0 _PG3_01|_DFF_P1|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_P1|1|1 _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|1|P _PG3_01|_DFF_P1|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|1|B _PG3_01|_DFF_P1|A1 _PG3_01|_DFF_P1|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|1|RB _PG3_01|_DFF_P1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|23|1 _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|23|B _PG3_01|_DFF_P1|A2 _PG3_01|_DFF_P1|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|23|RB _PG3_01|_DFF_P1|23|MID_SHUNT _PG3_01|_DFF_P1|A3  2.1704737578552e-12
B_PG3_01|_DFF_P1|3|1 _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|3|P _PG3_01|_DFF_P1|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|3|B _PG3_01|_DFF_P1|A3 _PG3_01|_DFF_P1|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|3|RB _PG3_01|_DFF_P1|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|4|1 _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|4|P _PG3_01|_DFF_P1|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|4|B _PG3_01|_DFF_P1|A4 _PG3_01|_DFF_P1|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|4|RB _PG3_01|_DFF_P1|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|T|1 _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|T|P _PG3_01|_DFF_P1|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|T|B _PG3_01|_DFF_P1|T1 _PG3_01|_DFF_P1|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|T|RB _PG3_01|_DFF_P1|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_P1|45|1 _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_P1|45|B _PG3_01|_DFF_P1|T2 _PG3_01|_DFF_P1|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_P1|45|RB _PG3_01|_DFF_P1|45|MID_SHUNT _PG3_01|_DFF_P1|A4  2.1704737578552e-12
B_PG3_01|_DFF_P1|6|1 _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_P1|6|P _PG3_01|_DFF_P1|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_P1|6|B _PG3_01|_DFF_P1|Q1 _PG3_01|_DFF_P1|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_P1|6|RB _PG3_01|_DFF_P1|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_PG|I_1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|I_1|MID  2e-12
I_PG3_01|_DFF_PG|I_1|B 0 _PG3_01|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|I_3|MID  2e-12
I_PG3_01|_DFF_PG|I_3|B 0 _PG3_01|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_PG|I_T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|I_T|MID  2e-12
I_PG3_01|_DFF_PG|I_T|B 0 _PG3_01|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_PG|I_6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|I_6|MID  2e-12
I_PG3_01|_DFF_PG|I_6|B 0 _PG3_01|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_PG|1|1 _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|1|P _PG3_01|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|1|B _PG3_01|_DFF_PG|A1 _PG3_01|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|1|RB _PG3_01|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|23|1 _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|23|B _PG3_01|_DFF_PG|A2 _PG3_01|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|23|RB _PG3_01|_DFF_PG|23|MID_SHUNT _PG3_01|_DFF_PG|A3  2.1704737578552e-12
B_PG3_01|_DFF_PG|3|1 _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|3|P _PG3_01|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|3|B _PG3_01|_DFF_PG|A3 _PG3_01|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|3|RB _PG3_01|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|4|1 _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|4|P _PG3_01|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|4|B _PG3_01|_DFF_PG|A4 _PG3_01|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|4|RB _PG3_01|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|T|1 _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|T|P _PG3_01|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|T|B _PG3_01|_DFF_PG|T1 _PG3_01|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|T|RB _PG3_01|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_PG|45|1 _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_PG|45|B _PG3_01|_DFF_PG|T2 _PG3_01|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_PG|45|RB _PG3_01|_DFF_PG|45|MID_SHUNT _PG3_01|_DFF_PG|A4  2.1704737578552e-12
B_PG3_01|_DFF_PG|6|1 _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_PG|6|P _PG3_01|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_PG|6|B _PG3_01|_DFF_PG|Q1 _PG3_01|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_PG|6|RB _PG3_01|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_DFF_GG|I_1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|I_1|MID  2e-12
I_PG3_01|_DFF_GG|I_1|B 0 _PG3_01|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|I_3|MID  2e-12
I_PG3_01|_DFF_GG|I_3|B 0 _PG3_01|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_01|_DFF_GG|I_T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|I_T|MID  2e-12
I_PG3_01|_DFF_GG|I_T|B 0 _PG3_01|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_DFF_GG|I_6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|I_6|MID  2e-12
I_PG3_01|_DFF_GG|I_6|B 0 _PG3_01|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_DFF_GG|1|1 _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|1|P _PG3_01|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|1|B _PG3_01|_DFF_GG|A1 _PG3_01|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|1|RB _PG3_01|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|23|1 _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|23|B _PG3_01|_DFF_GG|A2 _PG3_01|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|23|RB _PG3_01|_DFF_GG|23|MID_SHUNT _PG3_01|_DFF_GG|A3  2.1704737578552e-12
B_PG3_01|_DFF_GG|3|1 _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|3|P _PG3_01|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|3|B _PG3_01|_DFF_GG|A3 _PG3_01|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|3|RB _PG3_01|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|4|1 _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|4|P _PG3_01|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|4|B _PG3_01|_DFF_GG|A4 _PG3_01|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|4|RB _PG3_01|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|T|1 _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|T|P _PG3_01|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|T|B _PG3_01|_DFF_GG|T1 _PG3_01|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|T|RB _PG3_01|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_DFF_GG|45|1 _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_01|_DFF_GG|45|B _PG3_01|_DFF_GG|T2 _PG3_01|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_01|_DFF_GG|45|RB _PG3_01|_DFF_GG|45|MID_SHUNT _PG3_01|_DFF_GG|A4  2.1704737578552e-12
B_PG3_01|_DFF_GG|6|1 _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_DFF_GG|6|P _PG3_01|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_01|_DFF_GG|6|B _PG3_01|_DFF_GG|Q1 _PG3_01|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_01|_DFF_GG|6|RB _PG3_01|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_G|I_A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|I_A1|MID  2e-12
I_PG3_01|_AND_G|I_A1|B 0 _PG3_01|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|I_B1|MID  2e-12
I_PG3_01|_AND_G|I_B1|B 0 _PG3_01|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q3|B _PG3_01|_AND_G|Q3 _PG3_01|_AND_G|I_Q3|MID  2e-12
I_PG3_01|_AND_G|I_Q3|B 0 _PG3_01|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_G|I_Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|I_Q2|MID  2e-12
I_PG3_01|_AND_G|I_Q2|B 0 _PG3_01|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_G|I_Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|I_Q1|MID  2e-12
I_PG3_01|_AND_G|I_Q1|B 0 _PG3_01|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_G|A1|1 _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A1|P _PG3_01|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A1|B _PG3_01|_AND_G|A1 _PG3_01|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A1|RB _PG3_01|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A2|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|A2|P _PG3_01|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|A2|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|A2|RB _PG3_01|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|A12|1 _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|A12|B _PG3_01|_AND_G|A2 _PG3_01|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|A12|RB _PG3_01|_AND_G|A12|MID_SHUNT _PG3_01|_AND_G|A3  2.1704737578552e-12
B_PG3_01|_AND_G|B1|1 _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B1|P _PG3_01|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B1|B _PG3_01|_AND_G|B1 _PG3_01|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B1|RB _PG3_01|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B2|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|B2|P _PG3_01|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|B2|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|B2|RB _PG3_01|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|B12|1 _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_G|B12|B _PG3_01|_AND_G|B2 _PG3_01|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_G|B12|RB _PG3_01|_AND_G|B12|MID_SHUNT _PG3_01|_AND_G|B3  2.1704737578552e-12
B_PG3_01|_AND_G|Q2|1 _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q2|P _PG3_01|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q2|B _PG3_01|_AND_G|Q2 _PG3_01|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q2|RB _PG3_01|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_G|Q1|1 _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_G|Q1|P _PG3_01|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_G|Q1|B _PG3_01|_AND_G|Q1 _PG3_01|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_G|Q1|RB _PG3_01|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_01|_AND_P|I_A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|I_A1|MID  2e-12
I_PG3_01|_AND_P|I_A1|B 0 _PG3_01|_AND_P|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|I_B1|MID  2e-12
I_PG3_01|_AND_P|I_B1|B 0 _PG3_01|_AND_P|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q3|B _PG3_01|_AND_P|Q3 _PG3_01|_AND_P|I_Q3|MID  2e-12
I_PG3_01|_AND_P|I_Q3|B 0 _PG3_01|_AND_P|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_01|_AND_P|I_Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|I_Q2|MID  2e-12
I_PG3_01|_AND_P|I_Q2|B 0 _PG3_01|_AND_P|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_01|_AND_P|I_Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|I_Q1|MID  2e-12
I_PG3_01|_AND_P|I_Q1|B 0 _PG3_01|_AND_P|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_01|_AND_P|A1|1 _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A1|P _PG3_01|_AND_P|A1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A1|B _PG3_01|_AND_P|A1 _PG3_01|_AND_P|A1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A1|RB _PG3_01|_AND_P|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A2|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|A2|P _PG3_01|_AND_P|A2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|A2|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|A2|RB _PG3_01|_AND_P|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|A12|1 _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|A12|B _PG3_01|_AND_P|A2 _PG3_01|_AND_P|A12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|A12|RB _PG3_01|_AND_P|A12|MID_SHUNT _PG3_01|_AND_P|A3  2.1704737578552e-12
B_PG3_01|_AND_P|B1|1 _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B1|P _PG3_01|_AND_P|B1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B1|B _PG3_01|_AND_P|B1 _PG3_01|_AND_P|B1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B1|RB _PG3_01|_AND_P|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B2|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|B2|P _PG3_01|_AND_P|B2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|B2|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|B2|RB _PG3_01|_AND_P|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|B12|1 _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B3 JJMIT AREA=1.7857142857142858
R_PG3_01|_AND_P|B12|B _PG3_01|_AND_P|B2 _PG3_01|_AND_P|B12|MID_SHUNT  3.84154647408
L_PG3_01|_AND_P|B12|RB _PG3_01|_AND_P|B12|MID_SHUNT _PG3_01|_AND_P|B3  2.1704737578552e-12
B_PG3_01|_AND_P|Q2|1 _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q2|P _PG3_01|_AND_P|Q2|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q2|B _PG3_01|_AND_P|Q2 _PG3_01|_AND_P|Q2|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q2|RB _PG3_01|_AND_P|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_01|_AND_P|Q1|1 _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_01|_AND_P|Q1|P _PG3_01|_AND_P|Q1|MID_SERIES 0  2e-13
R_PG3_01|_AND_P|Q1|B _PG3_01|_AND_P|Q1 _PG3_01|_AND_P|Q1|MID_SHUNT  2.7439617672
L_PG3_01|_AND_P|Q1|RB _PG3_01|_AND_P|Q1|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL1|I_D1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|I_D1|MID  2e-12
ISPL_G1_1|SPL1|I_D1|B 0 SPL_G1_1|SPL1|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_D2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|I_D2|MID  2e-12
ISPL_G1_1|SPL1|I_D2|B 0 SPL_G1_1|SPL1|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL1|I_Q1|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|I_Q1|MID  2e-12
ISPL_G1_1|SPL1|I_Q1|B 0 SPL_G1_1|SPL1|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL1|I_Q2|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|I_Q2|MID  2e-12
ISPL_G1_1|SPL1|I_Q2|B 0 SPL_G1_1|SPL1|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL1|1|1 SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|1|P SPL_G1_1|SPL1|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|1|B SPL_G1_1|SPL1|D1 SPL_G1_1|SPL1|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|1|RB SPL_G1_1|SPL1|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|2|1 SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|2|P SPL_G1_1|SPL1|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|2|B SPL_G1_1|SPL1|D2 SPL_G1_1|SPL1|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|2|RB SPL_G1_1|SPL1|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|A|1 SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|A|P SPL_G1_1|SPL1|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|A|B SPL_G1_1|SPL1|QA1 SPL_G1_1|SPL1|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|A|RB SPL_G1_1|SPL1|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL1|B|1 SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL1|B|P SPL_G1_1|SPL1|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL1|B|B SPL_G1_1|SPL1|QB1 SPL_G1_1|SPL1|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL1|B|RB SPL_G1_1|SPL1|B|MID_SHUNT 0  1.550338398468e-12
LSPL_G1_1|SPL2|I_D1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|I_D1|MID  2e-12
ISPL_G1_1|SPL2|I_D1|B 0 SPL_G1_1|SPL2|I_D1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_D2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|I_D2|MID  2e-12
ISPL_G1_1|SPL2|I_D2|B 0 SPL_G1_1|SPL2|I_D2|MID  PWL(0 0 5e-12 0.000196)
LSPL_G1_1|SPL2|I_Q1|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|I_Q1|MID  2e-12
ISPL_G1_1|SPL2|I_Q1|B 0 SPL_G1_1|SPL2|I_Q1|MID  PWL(0 0 5e-12 0.00014)
LSPL_G1_1|SPL2|I_Q2|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|I_Q2|MID  2e-12
ISPL_G1_1|SPL2|I_Q2|B 0 SPL_G1_1|SPL2|I_Q2|MID  PWL(0 0 5e-12 0.00014)
BSPL_G1_1|SPL2|1|1 SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|1|P SPL_G1_1|SPL2|1|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|1|B SPL_G1_1|SPL2|D1 SPL_G1_1|SPL2|1|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|1|RB SPL_G1_1|SPL2|1|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|2|1 SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|2|P SPL_G1_1|SPL2|2|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|2|B SPL_G1_1|SPL2|D2 SPL_G1_1|SPL2|2|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|2|RB SPL_G1_1|SPL2|2|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|A|1 SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|A|P SPL_G1_1|SPL2|A|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|A|B SPL_G1_1|SPL2|QA1 SPL_G1_1|SPL2|A|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|A|RB SPL_G1_1|SPL2|A|MID_SHUNT 0  1.550338398468e-12
BSPL_G1_1|SPL2|B|1 SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SERIES JJMIT AREA=2.5
LSPL_G1_1|SPL2|B|P SPL_G1_1|SPL2|B|MID_SERIES 0  2e-13
RSPL_G1_1|SPL2|B|B SPL_G1_1|SPL2|QB1 SPL_G1_1|SPL2|B|MID_SHUNT  2.7439617672
LSPL_G1_1|SPL2|B|RB SPL_G1_1|SPL2|B|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|P|I_1|B _PG0_12|P|A1 _PG0_12|P|I_1|MID  2e-12
I_PG0_12|P|I_1|B 0 _PG0_12|P|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_3|B _PG0_12|P|A3 _PG0_12|P|I_3|MID  2e-12
I_PG0_12|P|I_3|B 0 _PG0_12|P|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|P|I_T|B _PG0_12|P|T1 _PG0_12|P|I_T|MID  2e-12
I_PG0_12|P|I_T|B 0 _PG0_12|P|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|P|I_6|B _PG0_12|P|Q1 _PG0_12|P|I_6|MID  2e-12
I_PG0_12|P|I_6|B 0 _PG0_12|P|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|P|1|1 _PG0_12|P|A1 _PG0_12|P|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|1|P _PG0_12|P|1|MID_SERIES 0  2e-13
R_PG0_12|P|1|B _PG0_12|P|A1 _PG0_12|P|1|MID_SHUNT  2.7439617672
L_PG0_12|P|1|RB _PG0_12|P|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|23|1 _PG0_12|P|A2 _PG0_12|P|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|P|23|B _PG0_12|P|A2 _PG0_12|P|23|MID_SHUNT  3.84154647408
L_PG0_12|P|23|RB _PG0_12|P|23|MID_SHUNT _PG0_12|P|A3  2.1704737578552e-12
B_PG0_12|P|3|1 _PG0_12|P|A3 _PG0_12|P|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|3|P _PG0_12|P|3|MID_SERIES 0  2e-13
R_PG0_12|P|3|B _PG0_12|P|A3 _PG0_12|P|3|MID_SHUNT  2.7439617672
L_PG0_12|P|3|RB _PG0_12|P|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|4|1 _PG0_12|P|A4 _PG0_12|P|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|4|P _PG0_12|P|4|MID_SERIES 0  2e-13
R_PG0_12|P|4|B _PG0_12|P|A4 _PG0_12|P|4|MID_SHUNT  2.7439617672
L_PG0_12|P|4|RB _PG0_12|P|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|T|1 _PG0_12|P|T1 _PG0_12|P|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|T|P _PG0_12|P|T|MID_SERIES 0  2e-13
R_PG0_12|P|T|B _PG0_12|P|T1 _PG0_12|P|T|MID_SHUNT  2.7439617672
L_PG0_12|P|T|RB _PG0_12|P|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|P|45|1 _PG0_12|P|T2 _PG0_12|P|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|P|45|B _PG0_12|P|T2 _PG0_12|P|45|MID_SHUNT  3.84154647408
L_PG0_12|P|45|RB _PG0_12|P|45|MID_SHUNT _PG0_12|P|A4  2.1704737578552e-12
B_PG0_12|P|6|1 _PG0_12|P|Q1 _PG0_12|P|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|P|6|P _PG0_12|P|6|MID_SERIES 0  2e-13
R_PG0_12|P|6|B _PG0_12|P|Q1 _PG0_12|P|6|MID_SHUNT  2.7439617672
L_PG0_12|P|6|RB _PG0_12|P|6|MID_SHUNT 0  1.550338398468e-12
L_PG0_12|G|I_1|B _PG0_12|G|A1 _PG0_12|G|I_1|MID  2e-12
I_PG0_12|G|I_1|B 0 _PG0_12|G|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_3|B _PG0_12|G|A3 _PG0_12|G|I_3|MID  2e-12
I_PG0_12|G|I_3|B 0 _PG0_12|G|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG0_12|G|I_T|B _PG0_12|G|T1 _PG0_12|G|I_T|MID  2e-12
I_PG0_12|G|I_T|B 0 _PG0_12|G|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG0_12|G|I_6|B _PG0_12|G|Q1 _PG0_12|G|I_6|MID  2e-12
I_PG0_12|G|I_6|B 0 _PG0_12|G|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG0_12|G|1|1 _PG0_12|G|A1 _PG0_12|G|1|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|1|P _PG0_12|G|1|MID_SERIES 0  2e-13
R_PG0_12|G|1|B _PG0_12|G|A1 _PG0_12|G|1|MID_SHUNT  2.7439617672
L_PG0_12|G|1|RB _PG0_12|G|1|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|23|1 _PG0_12|G|A2 _PG0_12|G|A3 JJMIT AREA=1.7857142857142858
R_PG0_12|G|23|B _PG0_12|G|A2 _PG0_12|G|23|MID_SHUNT  3.84154647408
L_PG0_12|G|23|RB _PG0_12|G|23|MID_SHUNT _PG0_12|G|A3  2.1704737578552e-12
B_PG0_12|G|3|1 _PG0_12|G|A3 _PG0_12|G|3|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|3|P _PG0_12|G|3|MID_SERIES 0  2e-13
R_PG0_12|G|3|B _PG0_12|G|A3 _PG0_12|G|3|MID_SHUNT  2.7439617672
L_PG0_12|G|3|RB _PG0_12|G|3|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|4|1 _PG0_12|G|A4 _PG0_12|G|4|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|4|P _PG0_12|G|4|MID_SERIES 0  2e-13
R_PG0_12|G|4|B _PG0_12|G|A4 _PG0_12|G|4|MID_SHUNT  2.7439617672
L_PG0_12|G|4|RB _PG0_12|G|4|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|T|1 _PG0_12|G|T1 _PG0_12|G|T|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|T|P _PG0_12|G|T|MID_SERIES 0  2e-13
R_PG0_12|G|T|B _PG0_12|G|T1 _PG0_12|G|T|MID_SHUNT  2.7439617672
L_PG0_12|G|T|RB _PG0_12|G|T|MID_SHUNT 0  1.550338398468e-12
B_PG0_12|G|45|1 _PG0_12|G|T2 _PG0_12|G|A4 JJMIT AREA=1.7857142857142858
R_PG0_12|G|45|B _PG0_12|G|T2 _PG0_12|G|45|MID_SHUNT  3.84154647408
L_PG0_12|G|45|RB _PG0_12|G|45|MID_SHUNT _PG0_12|G|A4  2.1704737578552e-12
B_PG0_12|G|6|1 _PG0_12|G|Q1 _PG0_12|G|6|MID_SERIES JJMIT AREA=2.5
L_PG0_12|G|6|P _PG0_12|G|6|MID_SERIES 0  2e-13
R_PG0_12|G|6|B _PG0_12|G|Q1 _PG0_12|G|6|MID_SHUNT  2.7439617672
L_PG0_12|G|6|RB _PG0_12|G|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_SPL_G1|I_D1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|I_D1|MID  2e-12
I_PG2_12|_SPL_G1|I_D1|B 0 _PG2_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_D2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|I_D2|MID  2e-12
I_PG2_12|_SPL_G1|I_D2|B 0 _PG2_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG2_12|_SPL_G1|I_Q1|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|I_Q1|MID  2e-12
I_PG2_12|_SPL_G1|I_Q1|B 0 _PG2_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG2_12|_SPL_G1|I_Q2|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|I_Q2|MID  2e-12
I_PG2_12|_SPL_G1|I_Q2|B 0 _PG2_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG2_12|_SPL_G1|1|1 _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|1|P _PG2_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|1|B _PG2_12|_SPL_G1|D1 _PG2_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|1|RB _PG2_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|2|1 _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|2|P _PG2_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|2|B _PG2_12|_SPL_G1|D2 _PG2_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|2|RB _PG2_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|A|1 _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|A|P _PG2_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|A|B _PG2_12|_SPL_G1|QA1 _PG2_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|A|RB _PG2_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_SPL_G1|B|1 _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_SPL_G1|B|P _PG2_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG2_12|_SPL_G1|B|B _PG2_12|_SPL_G1|QB1 _PG2_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG2_12|_SPL_G1|B|RB _PG2_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_PG|I_A1|B _PG2_12|_PG|A1 _PG2_12|_PG|I_A1|MID  2e-12
I_PG2_12|_PG|I_A1|B 0 _PG2_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_B1|B _PG2_12|_PG|B1 _PG2_12|_PG|I_B1|MID  2e-12
I_PG2_12|_PG|I_B1|B 0 _PG2_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q3|B _PG2_12|_PG|Q3 _PG2_12|_PG|I_Q3|MID  2e-12
I_PG2_12|_PG|I_Q3|B 0 _PG2_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_PG|I_Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|I_Q2|MID  2e-12
I_PG2_12|_PG|I_Q2|B 0 _PG2_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_PG|I_Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|I_Q1|MID  2e-12
I_PG2_12|_PG|I_Q1|B 0 _PG2_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_PG|A1|1 _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A1|P _PG2_12|_PG|A1|MID_SERIES 0  2e-13
R_PG2_12|_PG|A1|B _PG2_12|_PG|A1 _PG2_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A1|RB _PG2_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A2|1 _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|A2|P _PG2_12|_PG|A2|MID_SERIES 0  2e-13
R_PG2_12|_PG|A2|B _PG2_12|_PG|A2 _PG2_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|A2|RB _PG2_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|A12|1 _PG2_12|_PG|A2 _PG2_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|A12|B _PG2_12|_PG|A2 _PG2_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|A12|RB _PG2_12|_PG|A12|MID_SHUNT _PG2_12|_PG|A3  2.1704737578552e-12
B_PG2_12|_PG|B1|1 _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B1|P _PG2_12|_PG|B1|MID_SERIES 0  2e-13
R_PG2_12|_PG|B1|B _PG2_12|_PG|B1 _PG2_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B1|RB _PG2_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B2|1 _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|B2|P _PG2_12|_PG|B2|MID_SERIES 0  2e-13
R_PG2_12|_PG|B2|B _PG2_12|_PG|B2 _PG2_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|B2|RB _PG2_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|B12|1 _PG2_12|_PG|B2 _PG2_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_PG|B12|B _PG2_12|_PG|B2 _PG2_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_PG|B12|RB _PG2_12|_PG|B12|MID_SHUNT _PG2_12|_PG|B3  2.1704737578552e-12
B_PG2_12|_PG|Q2|1 _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q2|P _PG2_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q2|B _PG2_12|_PG|Q2 _PG2_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q2|RB _PG2_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_PG|Q1|1 _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_PG|Q1|P _PG2_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_PG|Q1|B _PG2_12|_PG|Q1 _PG2_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_PG|Q1|RB _PG2_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_GG|I_A1|B _PG2_12|_GG|A1 _PG2_12|_GG|I_A1|MID  2e-12
I_PG2_12|_GG|I_A1|B 0 _PG2_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_B1|B _PG2_12|_GG|B1 _PG2_12|_GG|I_B1|MID  2e-12
I_PG2_12|_GG|I_B1|B 0 _PG2_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q3|B _PG2_12|_GG|Q3 _PG2_12|_GG|I_Q3|MID  2e-12
I_PG2_12|_GG|I_Q3|B 0 _PG2_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_GG|I_Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|I_Q2|MID  2e-12
I_PG2_12|_GG|I_Q2|B 0 _PG2_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_GG|I_Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|I_Q1|MID  2e-12
I_PG2_12|_GG|I_Q1|B 0 _PG2_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_GG|A1|1 _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A1|P _PG2_12|_GG|A1|MID_SERIES 0  2e-13
R_PG2_12|_GG|A1|B _PG2_12|_GG|A1 _PG2_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A1|RB _PG2_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A2|1 _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|A2|P _PG2_12|_GG|A2|MID_SERIES 0  2e-13
R_PG2_12|_GG|A2|B _PG2_12|_GG|A2 _PG2_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|A2|RB _PG2_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|A12|1 _PG2_12|_GG|A2 _PG2_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|A12|B _PG2_12|_GG|A2 _PG2_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|A12|RB _PG2_12|_GG|A12|MID_SHUNT _PG2_12|_GG|A3  2.1704737578552e-12
B_PG2_12|_GG|B1|1 _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B1|P _PG2_12|_GG|B1|MID_SERIES 0  2e-13
R_PG2_12|_GG|B1|B _PG2_12|_GG|B1 _PG2_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B1|RB _PG2_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B2|1 _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|B2|P _PG2_12|_GG|B2|MID_SERIES 0  2e-13
R_PG2_12|_GG|B2|B _PG2_12|_GG|B2 _PG2_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|B2|RB _PG2_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|B12|1 _PG2_12|_GG|B2 _PG2_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_GG|B12|B _PG2_12|_GG|B2 _PG2_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG2_12|_GG|B12|RB _PG2_12|_GG|B12|MID_SHUNT _PG2_12|_GG|B3  2.1704737578552e-12
B_PG2_12|_GG|Q2|1 _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q2|P _PG2_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q2|B _PG2_12|_GG|Q2 _PG2_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q2|RB _PG2_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_GG|Q1|1 _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_GG|Q1|P _PG2_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG2_12|_GG|Q1|B _PG2_12|_GG|Q1 _PG2_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_GG|Q1|RB _PG2_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_PG|I_1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|I_1|MID  2e-12
I_PG2_12|_DFF_PG|I_1|B 0 _PG2_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|I_3|MID  2e-12
I_PG2_12|_DFF_PG|I_3|B 0 _PG2_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_PG|I_T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|I_T|MID  2e-12
I_PG2_12|_DFF_PG|I_T|B 0 _PG2_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_PG|I_6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|I_6|MID  2e-12
I_PG2_12|_DFF_PG|I_6|B 0 _PG2_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_PG|1|1 _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|1|P _PG2_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|1|B _PG2_12|_DFF_PG|A1 _PG2_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|1|RB _PG2_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|23|1 _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|23|B _PG2_12|_DFF_PG|A2 _PG2_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|23|RB _PG2_12|_DFF_PG|23|MID_SHUNT _PG2_12|_DFF_PG|A3  2.1704737578552e-12
B_PG2_12|_DFF_PG|3|1 _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|3|P _PG2_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|3|B _PG2_12|_DFF_PG|A3 _PG2_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|3|RB _PG2_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|4|1 _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|4|P _PG2_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|4|B _PG2_12|_DFF_PG|A4 _PG2_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|4|RB _PG2_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|T|1 _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|T|P _PG2_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|T|B _PG2_12|_DFF_PG|T1 _PG2_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|T|RB _PG2_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_PG|45|1 _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_PG|45|B _PG2_12|_DFF_PG|T2 _PG2_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_PG|45|RB _PG2_12|_DFF_PG|45|MID_SHUNT _PG2_12|_DFF_PG|A4  2.1704737578552e-12
B_PG2_12|_DFF_PG|6|1 _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_PG|6|P _PG2_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_PG|6|B _PG2_12|_DFF_PG|Q1 _PG2_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_PG|6|RB _PG2_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_DFF_GG|I_1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|I_1|MID  2e-12
I_PG2_12|_DFF_GG|I_1|B 0 _PG2_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|I_3|MID  2e-12
I_PG2_12|_DFF_GG|I_3|B 0 _PG2_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG2_12|_DFF_GG|I_T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|I_T|MID  2e-12
I_PG2_12|_DFF_GG|I_T|B 0 _PG2_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_DFF_GG|I_6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|I_6|MID  2e-12
I_PG2_12|_DFF_GG|I_6|B 0 _PG2_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_DFF_GG|1|1 _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|1|P _PG2_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|1|B _PG2_12|_DFF_GG|A1 _PG2_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|1|RB _PG2_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|23|1 _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|23|B _PG2_12|_DFF_GG|A2 _PG2_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|23|RB _PG2_12|_DFF_GG|23|MID_SHUNT _PG2_12|_DFF_GG|A3  2.1704737578552e-12
B_PG2_12|_DFF_GG|3|1 _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|3|P _PG2_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|3|B _PG2_12|_DFF_GG|A3 _PG2_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|3|RB _PG2_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|4|1 _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|4|P _PG2_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|4|B _PG2_12|_DFF_GG|A4 _PG2_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|4|RB _PG2_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|T|1 _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|T|P _PG2_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|T|B _PG2_12|_DFF_GG|T1 _PG2_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|T|RB _PG2_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_DFF_GG|45|1 _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG2_12|_DFF_GG|45|B _PG2_12|_DFF_GG|T2 _PG2_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG2_12|_DFF_GG|45|RB _PG2_12|_DFF_GG|45|MID_SHUNT _PG2_12|_DFF_GG|A4  2.1704737578552e-12
B_PG2_12|_DFF_GG|6|1 _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_DFF_GG|6|P _PG2_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG2_12|_DFF_GG|6|B _PG2_12|_DFF_GG|Q1 _PG2_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG2_12|_DFF_GG|6|RB _PG2_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG2_12|_AND_G|I_A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|I_A1|MID  2e-12
I_PG2_12|_AND_G|I_A1|B 0 _PG2_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|I_B1|MID  2e-12
I_PG2_12|_AND_G|I_B1|B 0 _PG2_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q3|B _PG2_12|_AND_G|Q3 _PG2_12|_AND_G|I_Q3|MID  2e-12
I_PG2_12|_AND_G|I_Q3|B 0 _PG2_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG2_12|_AND_G|I_Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|I_Q2|MID  2e-12
I_PG2_12|_AND_G|I_Q2|B 0 _PG2_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG2_12|_AND_G|I_Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|I_Q1|MID  2e-12
I_PG2_12|_AND_G|I_Q1|B 0 _PG2_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG2_12|_AND_G|A1|1 _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A1|P _PG2_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A1|B _PG2_12|_AND_G|A1 _PG2_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A1|RB _PG2_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A2|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|A2|P _PG2_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|A2|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|A2|RB _PG2_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|A12|1 _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|A12|B _PG2_12|_AND_G|A2 _PG2_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|A12|RB _PG2_12|_AND_G|A12|MID_SHUNT _PG2_12|_AND_G|A3  2.1704737578552e-12
B_PG2_12|_AND_G|B1|1 _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B1|P _PG2_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B1|B _PG2_12|_AND_G|B1 _PG2_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B1|RB _PG2_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B2|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|B2|P _PG2_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|B2|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|B2|RB _PG2_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|B12|1 _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG2_12|_AND_G|B12|B _PG2_12|_AND_G|B2 _PG2_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG2_12|_AND_G|B12|RB _PG2_12|_AND_G|B12|MID_SHUNT _PG2_12|_AND_G|B3  2.1704737578552e-12
B_PG2_12|_AND_G|Q2|1 _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q2|P _PG2_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q2|B _PG2_12|_AND_G|Q2 _PG2_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q2|RB _PG2_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG2_12|_AND_G|Q1|1 _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG2_12|_AND_G|Q1|P _PG2_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG2_12|_AND_G|Q1|B _PG2_12|_AND_G|Q1 _PG2_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG2_12|_AND_G|Q1|RB _PG2_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_SPL_G1|I_D1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|I_D1|MID  2e-12
I_PG3_12|_SPL_G1|I_D1|B 0 _PG3_12|_SPL_G1|I_D1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_D2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|I_D2|MID  2e-12
I_PG3_12|_SPL_G1|I_D2|B 0 _PG3_12|_SPL_G1|I_D2|MID  PWL(0 0 5e-12 0.0002205)
L_PG3_12|_SPL_G1|I_Q1|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|I_Q1|MID  2e-12
I_PG3_12|_SPL_G1|I_Q1|B 0 _PG3_12|_SPL_G1|I_Q1|MID  PWL(0 0 5e-12 0.0001575)
L_PG3_12|_SPL_G1|I_Q2|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|I_Q2|MID  2e-12
I_PG3_12|_SPL_G1|I_Q2|B 0 _PG3_12|_SPL_G1|I_Q2|MID  PWL(0 0 5e-12 0.0001575)
B_PG3_12|_SPL_G1|1|1 _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|1|P _PG3_12|_SPL_G1|1|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|1|B _PG3_12|_SPL_G1|D1 _PG3_12|_SPL_G1|1|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|1|RB _PG3_12|_SPL_G1|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|2|1 _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|2|P _PG3_12|_SPL_G1|2|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|2|B _PG3_12|_SPL_G1|D2 _PG3_12|_SPL_G1|2|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|2|RB _PG3_12|_SPL_G1|2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|A|1 _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|A|P _PG3_12|_SPL_G1|A|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|A|B _PG3_12|_SPL_G1|QA1 _PG3_12|_SPL_G1|A|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|A|RB _PG3_12|_SPL_G1|A|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_SPL_G1|B|1 _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_SPL_G1|B|P _PG3_12|_SPL_G1|B|MID_SERIES 0  2e-13
R_PG3_12|_SPL_G1|B|B _PG3_12|_SPL_G1|QB1 _PG3_12|_SPL_G1|B|MID_SHUNT  2.7439617672
L_PG3_12|_SPL_G1|B|RB _PG3_12|_SPL_G1|B|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_PG|I_A1|B _PG3_12|_PG|A1 _PG3_12|_PG|I_A1|MID  2e-12
I_PG3_12|_PG|I_A1|B 0 _PG3_12|_PG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_B1|B _PG3_12|_PG|B1 _PG3_12|_PG|I_B1|MID  2e-12
I_PG3_12|_PG|I_B1|B 0 _PG3_12|_PG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q3|B _PG3_12|_PG|Q3 _PG3_12|_PG|I_Q3|MID  2e-12
I_PG3_12|_PG|I_Q3|B 0 _PG3_12|_PG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_PG|I_Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|I_Q2|MID  2e-12
I_PG3_12|_PG|I_Q2|B 0 _PG3_12|_PG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_PG|I_Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|I_Q1|MID  2e-12
I_PG3_12|_PG|I_Q1|B 0 _PG3_12|_PG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_PG|A1|1 _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A1|P _PG3_12|_PG|A1|MID_SERIES 0  2e-13
R_PG3_12|_PG|A1|B _PG3_12|_PG|A1 _PG3_12|_PG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A1|RB _PG3_12|_PG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A2|1 _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|A2|P _PG3_12|_PG|A2|MID_SERIES 0  2e-13
R_PG3_12|_PG|A2|B _PG3_12|_PG|A2 _PG3_12|_PG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|A2|RB _PG3_12|_PG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|A12|1 _PG3_12|_PG|A2 _PG3_12|_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|A12|B _PG3_12|_PG|A2 _PG3_12|_PG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|A12|RB _PG3_12|_PG|A12|MID_SHUNT _PG3_12|_PG|A3  2.1704737578552e-12
B_PG3_12|_PG|B1|1 _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B1|P _PG3_12|_PG|B1|MID_SERIES 0  2e-13
R_PG3_12|_PG|B1|B _PG3_12|_PG|B1 _PG3_12|_PG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B1|RB _PG3_12|_PG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B2|1 _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|B2|P _PG3_12|_PG|B2|MID_SERIES 0  2e-13
R_PG3_12|_PG|B2|B _PG3_12|_PG|B2 _PG3_12|_PG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|B2|RB _PG3_12|_PG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|B12|1 _PG3_12|_PG|B2 _PG3_12|_PG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_PG|B12|B _PG3_12|_PG|B2 _PG3_12|_PG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_PG|B12|RB _PG3_12|_PG|B12|MID_SHUNT _PG3_12|_PG|B3  2.1704737578552e-12
B_PG3_12|_PG|Q2|1 _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q2|P _PG3_12|_PG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q2|B _PG3_12|_PG|Q2 _PG3_12|_PG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q2|RB _PG3_12|_PG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_PG|Q1|1 _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_PG|Q1|P _PG3_12|_PG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_PG|Q1|B _PG3_12|_PG|Q1 _PG3_12|_PG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_PG|Q1|RB _PG3_12|_PG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_GG|I_A1|B _PG3_12|_GG|A1 _PG3_12|_GG|I_A1|MID  2e-12
I_PG3_12|_GG|I_A1|B 0 _PG3_12|_GG|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_B1|B _PG3_12|_GG|B1 _PG3_12|_GG|I_B1|MID  2e-12
I_PG3_12|_GG|I_B1|B 0 _PG3_12|_GG|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q3|B _PG3_12|_GG|Q3 _PG3_12|_GG|I_Q3|MID  2e-12
I_PG3_12|_GG|I_Q3|B 0 _PG3_12|_GG|I_Q3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_GG|I_Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|I_Q2|MID  2e-12
I_PG3_12|_GG|I_Q2|B 0 _PG3_12|_GG|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_GG|I_Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|I_Q1|MID  2e-12
I_PG3_12|_GG|I_Q1|B 0 _PG3_12|_GG|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_GG|A1|1 _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A1|P _PG3_12|_GG|A1|MID_SERIES 0  2e-13
R_PG3_12|_GG|A1|B _PG3_12|_GG|A1 _PG3_12|_GG|A1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A1|RB _PG3_12|_GG|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A2|1 _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|A2|P _PG3_12|_GG|A2|MID_SERIES 0  2e-13
R_PG3_12|_GG|A2|B _PG3_12|_GG|A2 _PG3_12|_GG|A2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|A2|RB _PG3_12|_GG|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|A12|1 _PG3_12|_GG|A2 _PG3_12|_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|A12|B _PG3_12|_GG|A2 _PG3_12|_GG|A12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|A12|RB _PG3_12|_GG|A12|MID_SHUNT _PG3_12|_GG|A3  2.1704737578552e-12
B_PG3_12|_GG|B1|1 _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B1|P _PG3_12|_GG|B1|MID_SERIES 0  2e-13
R_PG3_12|_GG|B1|B _PG3_12|_GG|B1 _PG3_12|_GG|B1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B1|RB _PG3_12|_GG|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B2|1 _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|B2|P _PG3_12|_GG|B2|MID_SERIES 0  2e-13
R_PG3_12|_GG|B2|B _PG3_12|_GG|B2 _PG3_12|_GG|B2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|B2|RB _PG3_12|_GG|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|B12|1 _PG3_12|_GG|B2 _PG3_12|_GG|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_GG|B12|B _PG3_12|_GG|B2 _PG3_12|_GG|B12|MID_SHUNT  3.84154647408
L_PG3_12|_GG|B12|RB _PG3_12|_GG|B12|MID_SHUNT _PG3_12|_GG|B3  2.1704737578552e-12
B_PG3_12|_GG|Q2|1 _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q2|P _PG3_12|_GG|Q2|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q2|B _PG3_12|_GG|Q2 _PG3_12|_GG|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q2|RB _PG3_12|_GG|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_GG|Q1|1 _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_GG|Q1|P _PG3_12|_GG|Q1|MID_SERIES 0  2e-13
R_PG3_12|_GG|Q1|B _PG3_12|_GG|Q1 _PG3_12|_GG|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_GG|Q1|RB _PG3_12|_GG|Q1|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_PG|I_1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|I_1|MID  2e-12
I_PG3_12|_DFF_PG|I_1|B 0 _PG3_12|_DFF_PG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|I_3|MID  2e-12
I_PG3_12|_DFF_PG|I_3|B 0 _PG3_12|_DFF_PG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_PG|I_T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|I_T|MID  2e-12
I_PG3_12|_DFF_PG|I_T|B 0 _PG3_12|_DFF_PG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_PG|I_6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|I_6|MID  2e-12
I_PG3_12|_DFF_PG|I_6|B 0 _PG3_12|_DFF_PG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_PG|1|1 _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|1|P _PG3_12|_DFF_PG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|1|B _PG3_12|_DFF_PG|A1 _PG3_12|_DFF_PG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|1|RB _PG3_12|_DFF_PG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|23|1 _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|23|B _PG3_12|_DFF_PG|A2 _PG3_12|_DFF_PG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|23|RB _PG3_12|_DFF_PG|23|MID_SHUNT _PG3_12|_DFF_PG|A3  2.1704737578552e-12
B_PG3_12|_DFF_PG|3|1 _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|3|P _PG3_12|_DFF_PG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|3|B _PG3_12|_DFF_PG|A3 _PG3_12|_DFF_PG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|3|RB _PG3_12|_DFF_PG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|4|1 _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|4|P _PG3_12|_DFF_PG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|4|B _PG3_12|_DFF_PG|A4 _PG3_12|_DFF_PG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|4|RB _PG3_12|_DFF_PG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|T|1 _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|T|P _PG3_12|_DFF_PG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|T|B _PG3_12|_DFF_PG|T1 _PG3_12|_DFF_PG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|T|RB _PG3_12|_DFF_PG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_PG|45|1 _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_PG|45|B _PG3_12|_DFF_PG|T2 _PG3_12|_DFF_PG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_PG|45|RB _PG3_12|_DFF_PG|45|MID_SHUNT _PG3_12|_DFF_PG|A4  2.1704737578552e-12
B_PG3_12|_DFF_PG|6|1 _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_PG|6|P _PG3_12|_DFF_PG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_PG|6|B _PG3_12|_DFF_PG|Q1 _PG3_12|_DFF_PG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_PG|6|RB _PG3_12|_DFF_PG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_DFF_GG|I_1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|I_1|MID  2e-12
I_PG3_12|_DFF_GG|I_1|B 0 _PG3_12|_DFF_GG|I_1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|I_3|MID  2e-12
I_PG3_12|_DFF_GG|I_3|B 0 _PG3_12|_DFF_GG|I_3|MID  PWL(0 0 5e-12 0.00025)
L_PG3_12|_DFF_GG|I_T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|I_T|MID  2e-12
I_PG3_12|_DFF_GG|I_T|B 0 _PG3_12|_DFF_GG|I_T|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_DFF_GG|I_6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|I_6|MID  2e-12
I_PG3_12|_DFF_GG|I_6|B 0 _PG3_12|_DFF_GG|I_6|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_DFF_GG|1|1 _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|1|P _PG3_12|_DFF_GG|1|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|1|B _PG3_12|_DFF_GG|A1 _PG3_12|_DFF_GG|1|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|1|RB _PG3_12|_DFF_GG|1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|23|1 _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|23|B _PG3_12|_DFF_GG|A2 _PG3_12|_DFF_GG|23|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|23|RB _PG3_12|_DFF_GG|23|MID_SHUNT _PG3_12|_DFF_GG|A3  2.1704737578552e-12
B_PG3_12|_DFF_GG|3|1 _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|3|P _PG3_12|_DFF_GG|3|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|3|B _PG3_12|_DFF_GG|A3 _PG3_12|_DFF_GG|3|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|3|RB _PG3_12|_DFF_GG|3|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|4|1 _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|4|P _PG3_12|_DFF_GG|4|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|4|B _PG3_12|_DFF_GG|A4 _PG3_12|_DFF_GG|4|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|4|RB _PG3_12|_DFF_GG|4|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|T|1 _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|T|P _PG3_12|_DFF_GG|T|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|T|B _PG3_12|_DFF_GG|T1 _PG3_12|_DFF_GG|T|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|T|RB _PG3_12|_DFF_GG|T|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_DFF_GG|45|1 _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|A4 JJMIT AREA=1.7857142857142858
R_PG3_12|_DFF_GG|45|B _PG3_12|_DFF_GG|T2 _PG3_12|_DFF_GG|45|MID_SHUNT  3.84154647408
L_PG3_12|_DFF_GG|45|RB _PG3_12|_DFF_GG|45|MID_SHUNT _PG3_12|_DFF_GG|A4  2.1704737578552e-12
B_PG3_12|_DFF_GG|6|1 _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_DFF_GG|6|P _PG3_12|_DFF_GG|6|MID_SERIES 0  2e-13
R_PG3_12|_DFF_GG|6|B _PG3_12|_DFF_GG|Q1 _PG3_12|_DFF_GG|6|MID_SHUNT  2.7439617672
L_PG3_12|_DFF_GG|6|RB _PG3_12|_DFF_GG|6|MID_SHUNT 0  1.550338398468e-12
L_PG3_12|_AND_G|I_A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|I_A1|MID  2e-12
I_PG3_12|_AND_G|I_A1|B 0 _PG3_12|_AND_G|I_A1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|I_B1|MID  2e-12
I_PG3_12|_AND_G|I_B1|B 0 _PG3_12|_AND_G|I_B1|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q3|B _PG3_12|_AND_G|Q3 _PG3_12|_AND_G|I_Q3|MID  2e-12
I_PG3_12|_AND_G|I_Q3|B 0 _PG3_12|_AND_G|I_Q3|MID  PWL(0 0 5e-12 5e-05)
L_PG3_12|_AND_G|I_Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|I_Q2|MID  2e-12
I_PG3_12|_AND_G|I_Q2|B 0 _PG3_12|_AND_G|I_Q2|MID  PWL(0 0 5e-12 0.000175)
L_PG3_12|_AND_G|I_Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|I_Q1|MID  2e-12
I_PG3_12|_AND_G|I_Q1|B 0 _PG3_12|_AND_G|I_Q1|MID  PWL(0 0 5e-12 0.000175)
B_PG3_12|_AND_G|A1|1 _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A1|P _PG3_12|_AND_G|A1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A1|B _PG3_12|_AND_G|A1 _PG3_12|_AND_G|A1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A1|RB _PG3_12|_AND_G|A1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A2|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|A2|P _PG3_12|_AND_G|A2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|A2|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|A2|RB _PG3_12|_AND_G|A2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|A12|1 _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|A12|B _PG3_12|_AND_G|A2 _PG3_12|_AND_G|A12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|A12|RB _PG3_12|_AND_G|A12|MID_SHUNT _PG3_12|_AND_G|A3  2.1704737578552e-12
B_PG3_12|_AND_G|B1|1 _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B1|P _PG3_12|_AND_G|B1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B1|B _PG3_12|_AND_G|B1 _PG3_12|_AND_G|B1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B1|RB _PG3_12|_AND_G|B1|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B2|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|B2|P _PG3_12|_AND_G|B2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|B2|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|B2|RB _PG3_12|_AND_G|B2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|B12|1 _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B3 JJMIT AREA=1.7857142857142858
R_PG3_12|_AND_G|B12|B _PG3_12|_AND_G|B2 _PG3_12|_AND_G|B12|MID_SHUNT  3.84154647408
L_PG3_12|_AND_G|B12|RB _PG3_12|_AND_G|B12|MID_SHUNT _PG3_12|_AND_G|B3  2.1704737578552e-12
B_PG3_12|_AND_G|Q2|1 _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q2|P _PG3_12|_AND_G|Q2|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q2|B _PG3_12|_AND_G|Q2 _PG3_12|_AND_G|Q2|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q2|RB _PG3_12|_AND_G|Q2|MID_SHUNT 0  1.550338398468e-12
B_PG3_12|_AND_G|Q1|1 _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SERIES JJMIT AREA=2.5
L_PG3_12|_AND_G|Q1|P _PG3_12|_AND_G|Q1|MID_SERIES 0  2e-13
R_PG3_12|_AND_G|Q1|B _PG3_12|_AND_G|Q1 _PG3_12|_AND_G|Q1|MID_SHUNT  2.7439617672
L_PG3_12|_AND_G|Q1|RB _PG3_12|_AND_G|Q1|MID_SHUNT 0  1.550338398468e-12
.print DEVI R_S0
.print DEVI R_S1
.print DEVI R_S2
.print DEVI R_S3
.print DEVI R_S4
.print DEVI IA0|A
.print DEVI IB0|B
.print DEVI IA1|C
.print DEVI IB1|D
.print DEVI IA2|E
.print DEVI IB2|F
.print DEVI IA3|G
.print DEVI IB3|H
.print DEVI IT00|T
.print DEVI IT01|T
.print DEVI IT02|T
.print DEVI IT03|T
.print DEVI LSPL_IG0_0|1
.print DEVI LSPL_IG0_0|2
.print DEVI LSPL_IG0_0|3
.print DEVI LSPL_IG0_0|4
.print DEVI LSPL_IG0_0|5
.print DEVI LSPL_IG0_0|6
.print DEVI LSPL_IG0_0|7
.print DEVI LSPL_IP1_0|1
.print DEVI LSPL_IP1_0|2
.print DEVI LSPL_IP1_0|3
.print DEVI LSPL_IP1_0|4
.print DEVI LSPL_IP1_0|5
.print DEVI LSPL_IP1_0|6
.print DEVI LSPL_IP1_0|7
.print DEVI LSPL_IG2_0|1
.print DEVI LSPL_IG2_0|2
.print DEVI LSPL_IG2_0|3
.print DEVI LSPL_IG2_0|4
.print DEVI LSPL_IG2_0|5
.print DEVI LSPL_IG2_0|6
.print DEVI LSPL_IG2_0|7
.print DEVI LSPL_IP3_0|1
.print DEVI LSPL_IP3_0|2
.print DEVI LSPL_IP3_0|3
.print DEVI LSPL_IP3_0|4
.print DEVI LSPL_IP3_0|5
.print DEVI LSPL_IP3_0|6
.print DEVI LSPL_IP3_0|7
.print DEVI IT04|T
.print DEVI IT05|T
.print DEVI IT06|T
.print DEVI IT07|T
.print DEVI ID01|T
.print DEVI L_DFF_IP1_01|1
.print DEVI L_DFF_IP1_01|2
.print DEVI L_DFF_IP1_01|3
.print DEVI L_DFF_IP1_01|T
.print DEVI L_DFF_IP1_01|4
.print DEVI L_DFF_IP1_01|5
.print DEVI L_DFF_IP1_01|6
.print DEVI ID02|T
.print DEVI L_DFF_IP2_01|1
.print DEVI L_DFF_IP2_01|2
.print DEVI L_DFF_IP2_01|3
.print DEVI L_DFF_IP2_01|T
.print DEVI L_DFF_IP2_01|4
.print DEVI L_DFF_IP2_01|5
.print DEVI L_DFF_IP2_01|6
.print DEVI ID03|T
.print DEVI L_DFF_IP3_01|1
.print DEVI L_DFF_IP3_01|2
.print DEVI L_DFF_IP3_01|3
.print DEVI L_DFF_IP3_01|T
.print DEVI L_DFF_IP3_01|4
.print DEVI L_DFF_IP3_01|5
.print DEVI L_DFF_IP3_01|6
.print DEVI IT08|T
.print DEVI IT09|T
.print DEVI L_PG1_12|1
.print DEVI L_PG1_12|2
.print DEVI L_PG1_12|3
.print DEVI L_PG1_12|T
.print DEVI L_PG1_12|4
.print DEVI L_PG1_12|5
.print DEVI L_PG1_12|6
.print DEVI IT10|T
.print DEVI IT11|T
.print DEVI ID11|T
.print DEVI L_DFF_IP1_12|1
.print DEVI L_DFF_IP1_12|2
.print DEVI L_DFF_IP1_12|3
.print DEVI L_DFF_IP1_12|T
.print DEVI L_DFF_IP1_12|4
.print DEVI L_DFF_IP1_12|5
.print DEVI L_DFF_IP1_12|6
.print DEVI ID12|T
.print DEVI L_DFF_IP2_12|1
.print DEVI L_DFF_IP2_12|2
.print DEVI L_DFF_IP2_12|3
.print DEVI L_DFF_IP2_12|T
.print DEVI L_DFF_IP2_12|4
.print DEVI L_DFF_IP2_12|5
.print DEVI L_DFF_IP2_12|6
.print DEVI ID13|T
.print DEVI L_DFF_IP3_12|1
.print DEVI L_DFF_IP3_12|2
.print DEVI L_DFF_IP3_12|3
.print DEVI L_DFF_IP3_12|T
.print DEVI L_DFF_IP3_12|4
.print DEVI L_DFF_IP3_12|5
.print DEVI L_DFF_IP3_12|6
.print DEVI IT12|T
.print DEVI L_S0|1
.print DEVI L_S0|2
.print DEVI L_S0|3
.print DEVI L_S0|T
.print DEVI L_S0|4
.print DEVI L_S0|5
.print DEVI L_S0|6
.print DEVI IT13|T
.print DEVI BBUF_G0_2_TMP|1
.print DEVI BBUF_G0_2_TMP|2
.print DEVI BBUF_G0_2_TMP|3
.print DEVI BBUF_G0_2_TMP|4
.print DEVI IBUF_G0_2_TMP|B1
.print DEVI IBUF_G0_2_TMP|B2
.print DEVI IBUF_G0_2_TMP|B3
.print DEVI IBUF_G0_2_TMP|B4
.print DEVI LBUF_G0_2_TMP|1
.print DEVI LBUF_G0_2_TMP|2
.print DEVI LBUF_G0_2_TMP|3
.print DEVI LBUF_G0_2_TMP|4
.print DEVI LBUF_G0_2_TMP|5
.print DEVI LBUF_G0_2_TMP|P1
.print DEVI LBUF_G0_2_TMP|P2
.print DEVI LBUF_G0_2_TMP|P3
.print DEVI LBUF_G0_2_TMP|P4
.print DEVI LBUF_G0_2_TMP|B1
.print DEVI LBUF_G0_2_TMP|B2
.print DEVI LBUF_G0_2_TMP|B3
.print DEVI LBUF_G0_2_TMP|B4
.print DEVI RBUF_G0_2_TMP|B1
.print DEVI RBUF_G0_2_TMP|B2
.print DEVI RBUF_G0_2_TMP|B3
.print DEVI RBUF_G0_2_TMP|B4
.print DEVI LBUF_G0_2_TMP|RB1
.print DEVI LBUF_G0_2_TMP|RB2
.print DEVI LBUF_G0_2_TMP|RB3
.print DEVI LBUF_G0_2_TMP|RB4
.print DEVI LBUF_G0_2|1
.print DEVI LBUF_G0_2|2
.print DEVI LBUF_G0_2|3
.print DEVI LBUF_G0_2|4
.print DEVI BBUF_IP1_2_TMP|1
.print DEVI BBUF_IP1_2_TMP|2
.print DEVI BBUF_IP1_2_TMP|3
.print DEVI BBUF_IP1_2_TMP|4
.print DEVI IBUF_IP1_2_TMP|B1
.print DEVI IBUF_IP1_2_TMP|B2
.print DEVI IBUF_IP1_2_TMP|B3
.print DEVI IBUF_IP1_2_TMP|B4
.print DEVI LBUF_IP1_2_TMP|1
.print DEVI LBUF_IP1_2_TMP|2
.print DEVI LBUF_IP1_2_TMP|3
.print DEVI LBUF_IP1_2_TMP|4
.print DEVI LBUF_IP1_2_TMP|5
.print DEVI LBUF_IP1_2_TMP|P1
.print DEVI LBUF_IP1_2_TMP|P2
.print DEVI LBUF_IP1_2_TMP|P3
.print DEVI LBUF_IP1_2_TMP|P4
.print DEVI LBUF_IP1_2_TMP|B1
.print DEVI LBUF_IP1_2_TMP|B2
.print DEVI LBUF_IP1_2_TMP|B3
.print DEVI LBUF_IP1_2_TMP|B4
.print DEVI RBUF_IP1_2_TMP|B1
.print DEVI RBUF_IP1_2_TMP|B2
.print DEVI RBUF_IP1_2_TMP|B3
.print DEVI RBUF_IP1_2_TMP|B4
.print DEVI LBUF_IP1_2_TMP|RB1
.print DEVI LBUF_IP1_2_TMP|RB2
.print DEVI LBUF_IP1_2_TMP|RB3
.print DEVI LBUF_IP1_2_TMP|RB4
.print DEVI LBUF_IP1_2|1
.print DEVI LBUF_IP1_2|2
.print DEVI LBUF_IP1_2|3
.print DEVI LBUF_IP1_2|4
.print DEVI L_S1|A1
.print DEVI L_S1|A2
.print DEVI L_S1|A3
.print DEVI L_S1|B1
.print DEVI L_S1|B2
.print DEVI L_S1|B3
.print DEVI L_S1|T1
.print DEVI L_S1|T2
.print DEVI L_S1|Q2
.print DEVI L_S1|Q1
.print DEVI IT14|T
.print DEVI BBUF_G1_2_TMP|1
.print DEVI BBUF_G1_2_TMP|2
.print DEVI BBUF_G1_2_TMP|3
.print DEVI BBUF_G1_2_TMP|4
.print DEVI IBUF_G1_2_TMP|B1
.print DEVI IBUF_G1_2_TMP|B2
.print DEVI IBUF_G1_2_TMP|B3
.print DEVI IBUF_G1_2_TMP|B4
.print DEVI LBUF_G1_2_TMP|1
.print DEVI LBUF_G1_2_TMP|2
.print DEVI LBUF_G1_2_TMP|3
.print DEVI LBUF_G1_2_TMP|4
.print DEVI LBUF_G1_2_TMP|5
.print DEVI LBUF_G1_2_TMP|P1
.print DEVI LBUF_G1_2_TMP|P2
.print DEVI LBUF_G1_2_TMP|P3
.print DEVI LBUF_G1_2_TMP|P4
.print DEVI LBUF_G1_2_TMP|B1
.print DEVI LBUF_G1_2_TMP|B2
.print DEVI LBUF_G1_2_TMP|B3
.print DEVI LBUF_G1_2_TMP|B4
.print DEVI RBUF_G1_2_TMP|B1
.print DEVI RBUF_G1_2_TMP|B2
.print DEVI RBUF_G1_2_TMP|B3
.print DEVI RBUF_G1_2_TMP|B4
.print DEVI LBUF_G1_2_TMP|RB1
.print DEVI LBUF_G1_2_TMP|RB2
.print DEVI LBUF_G1_2_TMP|RB3
.print DEVI LBUF_G1_2_TMP|RB4
.print DEVI LBUF_G1_2|1
.print DEVI LBUF_G1_2|2
.print DEVI LBUF_G1_2|3
.print DEVI LBUF_G1_2|4
.print DEVI BBUF_IP2_2_TMP|1
.print DEVI BBUF_IP2_2_TMP|2
.print DEVI BBUF_IP2_2_TMP|3
.print DEVI BBUF_IP2_2_TMP|4
.print DEVI IBUF_IP2_2_TMP|B1
.print DEVI IBUF_IP2_2_TMP|B2
.print DEVI IBUF_IP2_2_TMP|B3
.print DEVI IBUF_IP2_2_TMP|B4
.print DEVI LBUF_IP2_2_TMP|1
.print DEVI LBUF_IP2_2_TMP|2
.print DEVI LBUF_IP2_2_TMP|3
.print DEVI LBUF_IP2_2_TMP|4
.print DEVI LBUF_IP2_2_TMP|5
.print DEVI LBUF_IP2_2_TMP|P1
.print DEVI LBUF_IP2_2_TMP|P2
.print DEVI LBUF_IP2_2_TMP|P3
.print DEVI LBUF_IP2_2_TMP|P4
.print DEVI LBUF_IP2_2_TMP|B1
.print DEVI LBUF_IP2_2_TMP|B2
.print DEVI LBUF_IP2_2_TMP|B3
.print DEVI LBUF_IP2_2_TMP|B4
.print DEVI RBUF_IP2_2_TMP|B1
.print DEVI RBUF_IP2_2_TMP|B2
.print DEVI RBUF_IP2_2_TMP|B3
.print DEVI RBUF_IP2_2_TMP|B4
.print DEVI LBUF_IP2_2_TMP|RB1
.print DEVI LBUF_IP2_2_TMP|RB2
.print DEVI LBUF_IP2_2_TMP|RB3
.print DEVI LBUF_IP2_2_TMP|RB4
.print DEVI LBUF_IP2_2|1
.print DEVI LBUF_IP2_2|2
.print DEVI LBUF_IP2_2|3
.print DEVI LBUF_IP2_2|4
.print DEVI L_S2|A1
.print DEVI L_S2|A2
.print DEVI L_S2|A3
.print DEVI L_S2|B1
.print DEVI L_S2|B2
.print DEVI L_S2|B3
.print DEVI L_S2|T1
.print DEVI L_S2|T2
.print DEVI L_S2|Q2
.print DEVI L_S2|Q1
.print DEVI IT15|T
.print DEVI BBUF_G2_2_TMP|1
.print DEVI BBUF_G2_2_TMP|2
.print DEVI BBUF_G2_2_TMP|3
.print DEVI BBUF_G2_2_TMP|4
.print DEVI IBUF_G2_2_TMP|B1
.print DEVI IBUF_G2_2_TMP|B2
.print DEVI IBUF_G2_2_TMP|B3
.print DEVI IBUF_G2_2_TMP|B4
.print DEVI LBUF_G2_2_TMP|1
.print DEVI LBUF_G2_2_TMP|2
.print DEVI LBUF_G2_2_TMP|3
.print DEVI LBUF_G2_2_TMP|4
.print DEVI LBUF_G2_2_TMP|5
.print DEVI LBUF_G2_2_TMP|P1
.print DEVI LBUF_G2_2_TMP|P2
.print DEVI LBUF_G2_2_TMP|P3
.print DEVI LBUF_G2_2_TMP|P4
.print DEVI LBUF_G2_2_TMP|B1
.print DEVI LBUF_G2_2_TMP|B2
.print DEVI LBUF_G2_2_TMP|B3
.print DEVI LBUF_G2_2_TMP|B4
.print DEVI RBUF_G2_2_TMP|B1
.print DEVI RBUF_G2_2_TMP|B2
.print DEVI RBUF_G2_2_TMP|B3
.print DEVI RBUF_G2_2_TMP|B4
.print DEVI LBUF_G2_2_TMP|RB1
.print DEVI LBUF_G2_2_TMP|RB2
.print DEVI LBUF_G2_2_TMP|RB3
.print DEVI LBUF_G2_2_TMP|RB4
.print DEVI LBUF_G2_2|1
.print DEVI LBUF_G2_2|2
.print DEVI LBUF_G2_2|3
.print DEVI LBUF_G2_2|4
.print DEVI L_S3|A1
.print DEVI L_S3|A2
.print DEVI L_S3|A3
.print DEVI L_S3|B1
.print DEVI L_S3|B2
.print DEVI L_S3|B3
.print DEVI L_S3|T1
.print DEVI L_S3|T2
.print DEVI L_S3|Q2
.print DEVI L_S3|Q1
.print DEVI IT16|T
.print DEVI L_S4|1
.print DEVI L_S4|2
.print DEVI L_S4|3
.print DEVI L_S4|T
.print DEVI L_S4|4
.print DEVI L_S4|5
.print DEVI L_S4|6
.print V IP1_2_TMP
.print V BUF_G0_2|1
.print V I3|B2
.print V BUF_G0_2_TMP|10
.print V _DFF_IP2_12|A2
.print V T14
.print V T08
.print V BUF_G0_2_TMP|11
.print V BUF_IP2_2_TMP|9
.print V BUF_IP2_2_TMP|101
.print V P2_1
.print V IG2_0_TO2
.print V BUF_G2_2_TMP|110
.print V _PG1_01|GG_SYNC
.print V BUF_G2_2_TMP|11
.print V _S4|A2
.print V _S0|A1
.print V _S0|A3
.print V G0_2_BUF
.print V _S0|Q1
.print V BUF_IP1_2_TMP|104
.print V _PG1_12|T1
.print V A1
.print V _S3|B1
.print V _S1|A3
.print V B3
.print V _DFF_IP2_01|A4
.print V _PG3_01|P1_COPY_2
.print V G1_2
.print V _S0|T1
.print V _DFF_IP1_01|Q1
.print V _S4|A1
.print V _S2|AB
.print V _PG2_12|PG
.print V _DFF_IP3_01|T1
.print V _PG1_12|Q1
.print V _S2|B2
.print V T06
.print V BUF_G0_2_TMP|9
.print V _DFF_IP2_12|T2
.print V G1_1_TO3
.print V BUF_IP2_2|6
.print V BUF_G0_2_TMP|2
.print V IP3_0_TO1
.print V BUF_G0_2_TMP|5
.print V BUF_G0_2_TMP|104
.print V BUF_IP2_2_TMP|107
.print V G2_2
.print V _S1|B2
.print V G0_2
.print V I1|B1
.print V BUF_G1_2_TMP|5
.print V _PG2_12|G1_COPY_1
.print V SPL_IP3_0|D2
.print V _S0|A2
.print V BUF_G1_2_TMP|7
.print V S3
.print V IP2_2_TMP
.print V BUF_G0_2_TMP|101
.print V BUF_IP1_2_TMP|110
.print V BUF_IP2_2_TMP|104
.print V SPL_IG2_0|JCT
.print V _S3|A1
.print V I1|A1_SYNC
.print V _S1|ABTQ
.print V _S3|B2
.print V BUF_G1_2_TMP|1
.print V T07
.print V BUF_G1_2_TMP|9
.print V _DFF_IP1_01|T2
.print V _S1|AB
.print V BUF_IP2_2_TMP|2
.print V I1|A1
.print V IG2_0_TO3
.print V BUF_G1_2_TMP|101
.print V _S2|B3
.print V SPL_IG0_0|QA1
.print V _PG1_12|A1
.print V BUF_G2_2|6
.print V I0|B2
.print V IP0_0
.print V _DFF_IP3_12|A1
.print V T13
.print V B2
.print V _DFF_IP3_12|A4
.print V _S2|A3
.print V _DFF_IP1_12|A1
.print V T12
.print V _DFF_IP3_01|A2
.print V _PG1_01|PG
.print V _S3|B3
.print V S4
.print V B0
.print V _PG1_12|A2
.print V T04
.print V _DFF_IP2_01|Q1
.print V BUF_G2_2_TMP|101
.print V SPL_IP3_0|QA1
.print V I2|A2
.print V BUF_IP2_2_TMP|3
.print V _S2|Q1
.print V T15
.print V _DFF_IP2_12|Q1
.print V BUF_G0_2_TMP|7
.print V SPL_IG2_0|QA1
.print V _PG3_12|GG
.print V _S1|T1
.print V T00
.print V BUF_G0_2_TMP|6
.print V IG0_0
.print V IP2_0_OUT
.print V BUF_IP1_2_TMP|12
.print V P3_1
.print V BUF_G2_2_TMP|2
.print V _PG3_01|G1_COPY_2
.print V BUF_G1_2_TMP|4
.print V SPL_IG0_0|D1
.print V G2_2_BUF
.print V _DFF_IP2_01|T1
.print V IP1_0_TO1
.print V _S2|B1
.print V G3_1
.print V BUF_IP2_2_TMP|5
.print V _DFF_IP3_12|A2
.print V BUF_IP2_2_TMP|1
.print V I3|A2
.print V _S4|Q1
.print V _DFF_IP3_12|A3
.print V _DFF_IP3_01|Q1
.print V _DFF_IP3_12|Q1
.print V IG1_0
.print V _PG3_01|PG
.print V _S3|A2
.print V BUF_G1_2_TMP|12
.print V BUF_G2_2_TMP|7
.print V BUF_IP1_2_TMP|8
.print V _DFF_IP1_01|A1
.print V I2|B1
.print V _DFF_IP1_12|A3
.print V _PG2_12|GG_SYNC
.print V P0_1
.print V BUF_IP2_2_TMP|11
.print V T11
.print V SPL_IP2_0|QTMP
.print V BUF_G1_2|4
.print V _DFF_IP3_01|A4
.print V _S0|T2
.print V _DFF_IP3_01|A1
.print V BUF_G0_2_TMP|1
.print V BUF_G2_2_TMP|3
.print V IP1_1_OUT
.print V BUF_G2_2_TMP|8
.print V BUF_IP1_2|1
.print V BUF_IP2_2|1
.print V SPL_IG2_0|D2
.print V T03
.print V _DFF_IP1_01|A4
.print V BUF_G2_2_TMP|1
.print V SPL_IG2_0|QB1
.print V BUF_IP1_2_TMP|3
.print V _PG3_12|G1_COPY_2
.print V BUF_IP1_2_TMP|11
.print V I2|B1_SYNC
.print V SPL_IG0_0|JCT
.print V G0_1
.print V _S3|A3
.print V G1_1_TO2
.print V _S4|T1
.print V IP1_0_OUT
.print V SPL_IP1_0|QB1
.print V BUF_IP1_2_TMP|101
.print V IG2_0
.print V I1|A2
.print V _PG3_01|G1_COPY_1
.print V BUF_G0_2_TMP|3
.print V A2
.print V _PG2_12|GG
.print V BUF_IP2_2_TMP|110
.print V SPL_IP1_0|D1
.print V BUF_G2_2_TMP|9
.print V SPL_IP3_0|JCT
.print V D12
.print V SPL_IG2_0|D1
.print V _PG1_12|A4
.print V _S2|T2
.print V SPL_IP1_0|JCT
.print V _DFF_IP1_12|T2
.print V IP1_2_OUT
.print V _S2|A1
.print V BUF_G0_2_TMP|107
.print V _S3|ABTQ
.print V BUF_G0_2_TMP|4
.print V _PG1_01|PG_SYNC
.print V IP1_0
.print V _DFF_IP1_01|T1
.print V BUF_IP2_2_TMP|4
.print V BUF_G2_2|4
.print V IP3_2_OUT
.print V I0|A1_SYNC
.print V BUF_IP1_2_TMP|10
.print V T09
.print V BUF_IP1_2|4
.print V G1_2_TMP
.print V I0|B1
.print V _PG3_01|GG_SYNC
.print V _DFF_IP1_12|A2
.print V _PG1_12|T2
.print V SPL_IG0_0|D2
.print V D11
.print V I3|A1
.print V _DFF_IP1_01|A3
.print V S1
.print V BUF_G2_2_TMP|104
.print V SPL_G1_1|QTMP
.print V _S2|ABTQ
.print V _DFF_IP1_12|T1
.print V _DFF_IP3_12|T2
.print V _S1|B3
.print V _PG2_12|G1_COPY_2
.print V S0
.print V I0|B1_SYNC
.print V BUF_G1_2_TMP|110
.print V _S3|T2
.print V BUF_G1_2_TMP|8
.print V _PG1_01|G1_COPY_1
.print V _DFF_IP3_01|A3
.print V IP2_1_OUT
.print V T16
.print V BUF_IP1_2_TMP|107
.print V _DFF_IP2_12|A3
.print V BUF_G0_2|6
.print V _PG3_01|GG
.print V _S0|A4
.print V BUF_IP1_2|6
.print V _DFF_IP2_01|A1
.print V _DFF_IP2_12|A4
.print V _PG3_12|PG
.print V _DFF_IP2_01|A3
.print V _PG1_01|G1_COPY_2
.print V _PG1_12|A3
.print V _S1|Q1
.print V SPL_IP3_0|D1
.print V BUF_G1_2_TMP|2
.print V IG3_0
.print V T01
.print V BUF_IP2_2_TMP|6
.print V BUF_G2_2_TMP|6
.print V _DFF_IP1_12|A4
.print V I1|B2
.print V SPL_IP1_0|D2
.print V I2|B2
.print V _DFF_IP3_01|T2
.print V BUF_G0_2_TMP|110
.print V BUF_G2_2_TMP|107
.print V G0_2_TMP
.print V _DFF_IP1_01|A2
.print V BUF_G2_2_TMP|5
.print V BUF_G1_2_TMP|107
.print V BUF_G2_2|1
.print V IP3_1_OUT
.print V IP3_0
.print V BUF_IP1_2_TMP|7
.print V G3_2
.print V A0
.print V A3
.print V _S1|T2
.print V IG0_0_TO1
.print V _PG3_12|G1_COPY_1
.print V BUF_G1_2_TMP|104
.print V IP1_2_OUT_BUF
.print V I2|A1_SYNC
.print V P0_2
.print V _S4|T2
.print V D02
.print V BUF_G0_2|4
.print V B1
.print V BUF_G0_2_TMP|12
.print V _S4|A3
.print V I3|B1_SYNC
.print V _PG3_12|GG_SYNC
.print V BUF_IP1_2_TMP|5
.print V _S1|A1
.print V _DFF_IP3_12|T1
.print V _S4|A4
.print V G2_2_TMP
.print V BUF_IP2_2_TMP|10
.print V S2
.print V _PG2_12|PG_SYNC
.print V BUF_IP1_2_TMP|9
.print V _DFF_IP1_12|Q1
.print V _PG3_01|PG_SYNC
.print V G1_2_BUF
.print V D03
.print V _PG3_01|P1_COPY_1
.print V _PG3_01|P0_SYNC
.print V _S3|AB
.print V BUF_IP1_2_TMP|6
.print V _DFF_IP2_12|A1
.print V BUF_G1_2_TMP|10
.print V T05
.print V I0|A2
.print V BUF_G2_2_TMP|12
.print V _S1|B1
.print V _DFF_IP2_01|T2
.print V BUF_G1_2_TMP|3
.print V _DFF_IP2_01|A2
.print V T02
.print V I2|A1
.print V _PG3_01|P1_SYNC
.print V I0|A1
.print V SPL_IG0_0|QB1
.print V BUF_IP2_2_TMP|12
.print V SPL_IP1_0|QA1
.print V BUF_IP1_2_TMP|1
.print V BUF_IP2_2|4
.print V BUF_G1_2|1
.print V IP3_0_OUT
.print V IP2_2_OUT_BUF
.print V I3|A1_SYNC
.print V _S1|A2
.print V T10
.print V BUF_G1_2|6
.print V I3|B1
.print V BUF_G2_2_TMP|10
.print V BUF_IP1_2_TMP|2
.print V IG0_0_TO0
.print V BUF_G0_2_TMP|8
.print V BUF_IP2_2_TMP|8
.print V D13
.print V _S2|A2
.print V _S3|Q1
.print V I1|B1_SYNC
.print V _PG3_12|PG_SYNC
.print V BUF_IP1_2_TMP|4
.print V BUF_G1_2_TMP|6
.print V IP2_0_TO2
.print V _PG1_01|GG
.print V _S2|T1
.print V G1_1_TO1
.print V IP2_0
.print V _S3|T1
.print V G2_1
.print V BUF_G2_2_TMP|4
.print V G1_1
.print V IP2_0_TO3
.print V IP2_2_OUT
.print V _DFF_IP2_12|T1
.print V SPL_IP3_0|QB1
.print V BUF_IP2_2_TMP|7
.print V D01
.print V BUF_G1_2_TMP|11
.print DEVP BBUF_G0_2_TMP|1
.print DEVP BBUF_G0_2_TMP|2
.print DEVP BBUF_G0_2_TMP|3
.print DEVP BBUF_G0_2_TMP|4
.print DEVP BBUF_IP1_2_TMP|1
.print DEVP BBUF_IP1_2_TMP|2
.print DEVP BBUF_IP1_2_TMP|3
.print DEVP BBUF_IP1_2_TMP|4
.print DEVP BBUF_G1_2_TMP|1
.print DEVP BBUF_G1_2_TMP|2
.print DEVP BBUF_G1_2_TMP|3
.print DEVP BBUF_G1_2_TMP|4
.print DEVP BBUF_IP2_2_TMP|1
.print DEVP BBUF_IP2_2_TMP|2
.print DEVP BBUF_IP2_2_TMP|3
.print DEVP BBUF_IP2_2_TMP|4
.print DEVP BBUF_G2_2_TMP|1
.print DEVP BBUF_G2_2_TMP|2
.print DEVP BBUF_G2_2_TMP|3
.print DEVP BBUF_G2_2_TMP|4
