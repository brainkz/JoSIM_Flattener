*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM TCLOCK=1e-10
.PARAM GLOBAL_SCALE=1.1
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.5E-12 800E-12
ROUT N1001 0  1
IA|A 0 A_IN  PWL(0 0 1.17e-10 0 1.2e-10 0.0007 1.23e-10 0 3.17e-10 0 3.2e-10 0.0007 3.23e-10 0 5.17e-10 0 5.2e-10 0.0007 5.23e-10 0 7.17e-10 0 7.2e-10 0.0007 7.23e-10 0 9.17e-10 0 9.2e-10 0.0007 9.23e-10 0 1.117e-09 0 1.12e-09 0.0007 1.123e-09 0 1.317e-09 0 1.32e-09 0.0007 1.323e-09 0 1.517e-09 0 1.52e-09 0.0007 1.523e-09 0 1.717e-09 0 1.72e-09 0.0007 1.723e-09 0 1.917e-09 0 1.92e-09 0.0007 1.923e-09 0 2.117e-09 0 2.12e-09 0.0007 2.123e-09 0 2.317e-09 0 2.32e-09 0.0007 2.323e-09 0 2.517e-09 0 2.52e-09 0.0007 2.523e-09 0 2.717e-09 0 2.72e-09 0.0007 2.723e-09 0 2.917e-09 0 2.92e-09 0.0007 2.923e-09 0 3.117e-09 0 3.12e-09 0.0007 3.123e-09 0 3.317e-09 0 3.32e-09 0.0007 3.323e-09 0 3.517e-09 0 3.52e-09 0.0007 3.523e-09 0 3.717e-09 0 3.72e-09 0.0007 3.723e-09 0 3.917e-09 0 3.92e-09 0.0007 3.923e-09 0 4.117e-09 0 4.12e-09 0.0007 4.123e-09 0 4.317e-09 0 4.32e-09 0.0007 4.323e-09 0 4.517e-09 0 4.52e-09 0.0007 4.523e-09 0 4.717e-09 0 4.72e-09 0.0007 4.723e-09 0 4.917e-09 0 4.92e-09 0.0007 4.923e-09 0 5.117e-09 0 5.12e-09 0.0007 5.123e-09 0 5.317e-09 0 5.32e-09 0.0007 5.323e-09 0 5.517e-09 0 5.52e-09 0.0007 5.523e-09 0 5.717e-09 0 5.72e-09 0.0007 5.723e-09 0 5.917e-09 0 5.92e-09 0.0007 5.923e-09 0 6.117e-09 0 6.12e-09 0.0007 6.123e-09 0 6.317e-09 0 6.32e-09 0.0007 6.323e-09 0 6.517e-09 0 6.52e-09 0.0007 6.523e-09 0 6.717e-09 0 6.72e-09 0.0007 6.723e-09 0 6.917e-09 0 6.92e-09 0.0007 6.923e-09 0 7.117e-09 0 7.12e-09 0.0007 7.123e-09 0 7.317e-09 0 7.32e-09 0.0007 7.323e-09 0 7.517e-09 0 7.52e-09 0.0007 7.523e-09 0 7.717e-09 0 7.72e-09 0.0007 7.723e-09 0 7.917e-09 0 7.92e-09 0.0007 7.923e-09 0 8.117e-09 0 8.12e-09 0.0007 8.123e-09 0 8.317e-09 0 8.32e-09 0.0007 8.323e-09 0 8.517e-09 0 8.52e-09 0.0007 8.523e-09 0 8.717e-09 0 8.72e-09 0.0007 8.723e-09 0 8.917e-09 0 8.92e-09 0.0007 8.923e-09 0 9.117e-09 0 9.12e-09 0.0007 9.123e-09 0 9.317e-09 0 9.32e-09 0.0007 9.323e-09 0 9.517e-09 0 9.52e-09 0.0007 9.523e-09 0 9.717e-09 0 9.72e-09 0.0007 9.723e-09 0 9.917e-09 0 9.92e-09 0.0007 9.923e-09 0 1.0117e-08 0 1.012e-08 0.0007 1.0123e-08 0 1.0317e-08 0 1.032e-08 0.0007 1.0323e-08 0 1.0517e-08 0 1.052e-08 0.0007 1.0523e-08 0 1.0717e-08 0 1.072e-08 0.0007 1.0723e-08 0 1.0917e-08 0 1.092e-08 0.0007 1.0923e-08 0 1.1117e-08 0 1.112e-08 0.0007 1.1123e-08 0 1.1317e-08 0 1.132e-08 0.0007 1.1323e-08 0 1.1517e-08 0 1.152e-08 0.0007 1.1523e-08 0 1.1717e-08 0 1.172e-08 0.0007 1.1723e-08 0 1.1917e-08 0 1.192e-08 0.0007 1.1923e-08 0 1.2117e-08 0 1.212e-08 0.0007 1.2123e-08 0 1.2317e-08 0 1.232e-08 0.0007 1.2323e-08 0 1.2517e-08 0 1.252e-08 0.0007 1.2523e-08 0 1.2717e-08 0 1.272e-08 0.0007 1.2723e-08 0 1.2917e-08 0 1.292e-08 0.0007 1.2923e-08 0 1.3117e-08 0 1.312e-08 0.0007 1.3123e-08 0 1.3317e-08 0 1.332e-08 0.0007 1.3323e-08 0 1.3517e-08 0 1.352e-08 0.0007 1.3523e-08 0 1.3717e-08 0 1.372e-08 0.0007 1.3723e-08 0 1.3917e-08 0 1.392e-08 0.0007 1.3923e-08 0 1.4117e-08 0 1.412e-08 0.0007 1.4123e-08 0 1.4317e-08 0 1.432e-08 0.0007 1.4323e-08 0 1.4517e-08 0 1.452e-08 0.0007 1.4523e-08 0 1.4717e-08 0 1.472e-08 0.0007 1.4723e-08 0 1.4917e-08 0 1.492e-08 0.0007 1.4923e-08 0 1.5117e-08 0 1.512e-08 0.0007 1.5123e-08 0 1.5317e-08 0 1.532e-08 0.0007 1.5323e-08 0 1.5517e-08 0 1.552e-08 0.0007 1.5523e-08 0 1.5717e-08 0 1.572e-08 0.0007 1.5723e-08 0 1.5917e-08 0 1.592e-08 0.0007 1.5923e-08 0 1.6117e-08 0 1.612e-08 0.0007 1.6123e-08 0 1.6317e-08 0 1.632e-08 0.0007 1.6323e-08 0 1.6517e-08 0 1.652e-08 0.0007 1.6523e-08 0 1.6717e-08 0 1.672e-08 0.0007 1.6723e-08 0 1.6917e-08 0 1.692e-08 0.0007 1.6923e-08 0 1.7117e-08 0 1.712e-08 0.0007 1.7123e-08 0 1.7317e-08 0 1.732e-08 0.0007 1.7323e-08 0 1.7517e-08 0 1.752e-08 0.0007 1.7523e-08 0 1.7717e-08 0 1.772e-08 0.0007 1.7723e-08 0 1.7917e-08 0 1.792e-08 0.0007 1.7923e-08 0 1.8117e-08 0 1.812e-08 0.0007 1.8123e-08 0 1.8317e-08 0 1.832e-08 0.0007 1.8323e-08 0 1.8517e-08 0 1.852e-08 0.0007 1.8523e-08 0 1.8717e-08 0 1.872e-08 0.0007 1.8723e-08 0 1.8917e-08 0 1.892e-08 0.0007 1.8923e-08 0 1.9117e-08 0 1.912e-08 0.0007 1.9123e-08 0 1.9317e-08 0 1.932e-08 0.0007 1.9323e-08 0 1.9517e-08 0 1.952e-08 0.0007 1.9523e-08 0 1.9717e-08 0 1.972e-08 0.0007 1.9723e-08 0 1.9917e-08 0 1.992e-08 0.0007 1.9923e-08 0 2.0117e-08 0 2.012e-08 0.0007 2.0123e-08 0 2.0317e-08 0 2.032e-08 0.0007 2.0323e-08 0 2.0517e-08 0 2.052e-08 0.0007 2.0523e-08 0 2.0717e-08 0 2.072e-08 0.0007 2.0723e-08 0 2.0917e-08 0 2.092e-08 0.0007 2.0923e-08 0 2.1117e-08 0 2.112e-08 0.0007 2.1123e-08 0 2.1317e-08 0 2.132e-08 0.0007 2.1323e-08 0 2.1517e-08 0 2.152e-08 0.0007 2.1523e-08 0 2.1717e-08 0 2.172e-08 0.0007 2.1723e-08 0 2.1917e-08 0 2.192e-08 0.0007 2.1923e-08 0 2.2117e-08 0 2.212e-08 0.0007 2.2123e-08 0 2.2317e-08 0 2.232e-08 0.0007 2.2323e-08 0 2.2517e-08 0 2.252e-08 0.0007 2.2523e-08 0 2.2717e-08 0 2.272e-08 0.0007 2.2723e-08 0 2.2917e-08 0 2.292e-08 0.0007 2.2923e-08 0 2.3117e-08 0 2.312e-08 0.0007 2.3123e-08 0 2.3317e-08 0 2.332e-08 0.0007 2.3323e-08 0 2.3517e-08 0 2.352e-08 0.0007 2.3523e-08 0 2.3717e-08 0 2.372e-08 0.0007 2.3723e-08 0 2.3917e-08 0 2.392e-08 0.0007 2.3923e-08 0 2.4117e-08 0 2.412e-08 0.0007 2.4123e-08 0 2.4317e-08 0 2.432e-08 0.0007 2.4323e-08 0 2.4517e-08 0 2.452e-08 0.0007 2.4523e-08 0 2.4717e-08 0 2.472e-08 0.0007 2.4723e-08 0 2.4917e-08 0 2.492e-08 0.0007 2.4923e-08 0 2.5117e-08 0 2.512e-08 0.0007 2.5123e-08 0 2.5317e-08 0 2.532e-08 0.0007 2.5323e-08 0 2.5517e-08 0 2.552e-08 0.0007 2.5523e-08 0)
IB|B 0 B_IN  PWL(0 0 2.27e-10 0 2.3e-10 0.0007 2.33e-10 0 3.27e-10 0 3.3e-10 0.0007 3.33e-10 0 6.27e-10 0 6.3e-10 0.0007 6.33e-10 0 7.27e-10 0 7.3e-10 0.0007 7.33e-10 0 1.027e-09 0 1.03e-09 0.0007 1.033e-09 0 1.127e-09 0 1.13e-09 0.0007 1.133e-09 0 1.427e-09 0 1.43e-09 0.0007 1.433e-09 0 1.527e-09 0 1.53e-09 0.0007 1.533e-09 0 1.827e-09 0 1.83e-09 0.0007 1.833e-09 0 1.927e-09 0 1.93e-09 0.0007 1.933e-09 0 2.227e-09 0 2.23e-09 0.0007 2.233e-09 0 2.327e-09 0 2.33e-09 0.0007 2.333e-09 0 2.627e-09 0 2.63e-09 0.0007 2.633e-09 0 2.727e-09 0 2.73e-09 0.0007 2.733e-09 0 3.027e-09 0 3.03e-09 0.0007 3.033e-09 0 3.127e-09 0 3.13e-09 0.0007 3.133e-09 0 3.427e-09 0 3.43e-09 0.0007 3.433e-09 0 3.527e-09 0 3.53e-09 0.0007 3.533e-09 0 3.827e-09 0 3.83e-09 0.0007 3.833e-09 0 3.927e-09 0 3.93e-09 0.0007 3.933e-09 0 4.227e-09 0 4.23e-09 0.0007 4.233e-09 0 4.327e-09 0 4.33e-09 0.0007 4.333e-09 0 4.627e-09 0 4.63e-09 0.0007 4.633e-09 0 4.727e-09 0 4.73e-09 0.0007 4.733e-09 0 5.027e-09 0 5.03e-09 0.0007 5.033e-09 0 5.127e-09 0 5.13e-09 0.0007 5.133e-09 0 5.427e-09 0 5.43e-09 0.0007 5.433e-09 0 5.527e-09 0 5.53e-09 0.0007 5.533e-09 0 5.827e-09 0 5.83e-09 0.0007 5.833e-09 0 5.927e-09 0 5.93e-09 0.0007 5.933e-09 0 6.227e-09 0 6.23e-09 0.0007 6.233e-09 0 6.327e-09 0 6.33e-09 0.0007 6.333e-09 0 6.627e-09 0 6.63e-09 0.0007 6.633e-09 0 6.727e-09 0 6.73e-09 0.0007 6.733e-09 0 7.027e-09 0 7.03e-09 0.0007 7.033e-09 0 7.127e-09 0 7.13e-09 0.0007 7.133e-09 0 7.427e-09 0 7.43e-09 0.0007 7.433e-09 0 7.527e-09 0 7.53e-09 0.0007 7.533e-09 0 7.827e-09 0 7.83e-09 0.0007 7.833e-09 0 7.927e-09 0 7.93e-09 0.0007 7.933e-09 0 8.227e-09 0 8.23e-09 0.0007 8.233e-09 0 8.327e-09 0 8.33e-09 0.0007 8.333e-09 0 8.627e-09 0 8.63e-09 0.0007 8.633e-09 0 8.727e-09 0 8.73e-09 0.0007 8.733e-09 0 9.027e-09 0 9.03e-09 0.0007 9.033e-09 0 9.127e-09 0 9.13e-09 0.0007 9.133e-09 0 9.427e-09 0 9.43e-09 0.0007 9.433e-09 0 9.527e-09 0 9.53e-09 0.0007 9.533e-09 0 9.827e-09 0 9.83e-09 0.0007 9.833e-09 0 9.927e-09 0 9.93e-09 0.0007 9.933e-09 0 1.0227e-08 0 1.023e-08 0.0007 1.0233e-08 0 1.0327e-08 0 1.033e-08 0.0007 1.0333e-08 0 1.0627e-08 0 1.063e-08 0.0007 1.0633e-08 0 1.0727e-08 0 1.073e-08 0.0007 1.0733e-08 0 1.1027e-08 0 1.103e-08 0.0007 1.1033e-08 0 1.1127e-08 0 1.113e-08 0.0007 1.1133e-08 0 1.1427e-08 0 1.143e-08 0.0007 1.1433e-08 0 1.1527e-08 0 1.153e-08 0.0007 1.1533e-08 0 1.1827e-08 0 1.183e-08 0.0007 1.1833e-08 0 1.1927e-08 0 1.193e-08 0.0007 1.1933e-08 0 1.2227e-08 0 1.223e-08 0.0007 1.2233e-08 0 1.2327e-08 0 1.233e-08 0.0007 1.2333e-08 0 1.2627e-08 0 1.263e-08 0.0007 1.2633e-08 0 1.2727e-08 0 1.273e-08 0.0007 1.2733e-08 0 1.3027e-08 0 1.303e-08 0.0007 1.3033e-08 0 1.3127e-08 0 1.313e-08 0.0007 1.3133e-08 0 1.3427e-08 0 1.343e-08 0.0007 1.3433e-08 0 1.3527e-08 0 1.353e-08 0.0007 1.3533e-08 0 1.3827e-08 0 1.383e-08 0.0007 1.3833e-08 0 1.3927e-08 0 1.393e-08 0.0007 1.3933e-08 0 1.4227e-08 0 1.423e-08 0.0007 1.4233e-08 0 1.4327e-08 0 1.433e-08 0.0007 1.4333e-08 0 1.4627e-08 0 1.463e-08 0.0007 1.4633e-08 0 1.4727e-08 0 1.473e-08 0.0007 1.4733e-08 0 1.5027e-08 0 1.503e-08 0.0007 1.5033e-08 0 1.5127e-08 0 1.513e-08 0.0007 1.5133e-08 0 1.5427e-08 0 1.543e-08 0.0007 1.5433e-08 0 1.5527e-08 0 1.553e-08 0.0007 1.5533e-08 0 1.5827e-08 0 1.583e-08 0.0007 1.5833e-08 0 1.5927e-08 0 1.593e-08 0.0007 1.5933e-08 0 1.6227e-08 0 1.623e-08 0.0007 1.6233e-08 0 1.6327e-08 0 1.633e-08 0.0007 1.6333e-08 0 1.6627e-08 0 1.663e-08 0.0007 1.6633e-08 0 1.6727e-08 0 1.673e-08 0.0007 1.6733e-08 0 1.7027e-08 0 1.703e-08 0.0007 1.7033e-08 0 1.7127e-08 0 1.713e-08 0.0007 1.7133e-08 0 1.7427e-08 0 1.743e-08 0.0007 1.7433e-08 0 1.7527e-08 0 1.753e-08 0.0007 1.7533e-08 0 1.7827e-08 0 1.783e-08 0.0007 1.7833e-08 0 1.7927e-08 0 1.793e-08 0.0007 1.7933e-08 0 1.8227e-08 0 1.823e-08 0.0007 1.8233e-08 0 1.8327e-08 0 1.833e-08 0.0007 1.8333e-08 0 1.8627e-08 0 1.863e-08 0.0007 1.8633e-08 0 1.8727e-08 0 1.873e-08 0.0007 1.8733e-08 0 1.9027e-08 0 1.903e-08 0.0007 1.9033e-08 0 1.9127e-08 0 1.913e-08 0.0007 1.9133e-08 0 1.9427e-08 0 1.943e-08 0.0007 1.9433e-08 0 1.9527e-08 0 1.953e-08 0.0007 1.9533e-08 0 1.9827e-08 0 1.983e-08 0.0007 1.9833e-08 0 1.9927e-08 0 1.993e-08 0.0007 1.9933e-08 0 2.0227e-08 0 2.023e-08 0.0007 2.0233e-08 0 2.0327e-08 0 2.033e-08 0.0007 2.0333e-08 0 2.0627e-08 0 2.063e-08 0.0007 2.0633e-08 0 2.0727e-08 0 2.073e-08 0.0007 2.0733e-08 0 2.1027e-08 0 2.103e-08 0.0007 2.1033e-08 0 2.1127e-08 0 2.113e-08 0.0007 2.1133e-08 0 2.1427e-08 0 2.143e-08 0.0007 2.1433e-08 0 2.1527e-08 0 2.153e-08 0.0007 2.1533e-08 0 2.1827e-08 0 2.183e-08 0.0007 2.1833e-08 0 2.1927e-08 0 2.193e-08 0.0007 2.1933e-08 0 2.2227e-08 0 2.223e-08 0.0007 2.2233e-08 0 2.2327e-08 0 2.233e-08 0.0007 2.2333e-08 0 2.2627e-08 0 2.263e-08 0.0007 2.2633e-08 0 2.2727e-08 0 2.273e-08 0.0007 2.2733e-08 0 2.3027e-08 0 2.303e-08 0.0007 2.3033e-08 0 2.3127e-08 0 2.313e-08 0.0007 2.3133e-08 0 2.3427e-08 0 2.343e-08 0.0007 2.3433e-08 0 2.3527e-08 0 2.353e-08 0.0007 2.3533e-08 0 2.3827e-08 0 2.383e-08 0.0007 2.3833e-08 0 2.3927e-08 0 2.393e-08 0.0007 2.3933e-08 0 2.4227e-08 0 2.423e-08 0.0007 2.4233e-08 0 2.4327e-08 0 2.433e-08 0.0007 2.4333e-08 0 2.4627e-08 0 2.463e-08 0.0007 2.4633e-08 0 2.4727e-08 0 2.473e-08 0.0007 2.4733e-08 0 2.5027e-08 0 2.503e-08 0.0007 2.5033e-08 0 2.5127e-08 0 2.513e-08 0.0007 2.5133e-08 0 2.5427e-08 0 2.543e-08 0.0007 2.5433e-08 0 2.5527e-08 0 2.553e-08 0.0007 2.5533e-08 0)
IT1|T 0 CLK1  PWL(0 0 9.7e-11 0 1e-10 0.0007 1.03e-10 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 2.97e-10 0 3e-10 0.0007 3.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 4.97e-10 0 5e-10 0.0007 5.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 6.97e-10 0 7e-10 0.0007 7.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 8.97e-10 0 9e-10 0.0007 9.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.097e-09 0 1.1e-09 0.0007 1.103e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.297e-09 0 1.3e-09 0.0007 1.303e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.497e-09 0 1.5e-09 0.0007 1.503e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.697e-09 0 1.7e-09 0.0007 1.703e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.897e-09 0 1.9e-09 0.0007 1.903e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.097e-09 0 2.1e-09 0.0007 2.103e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.297e-09 0 2.3e-09 0.0007 2.303e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.497e-09 0 2.5e-09 0.0007 2.503e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.697e-09 0 2.7e-09 0.0007 2.703e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.897e-09 0 2.9e-09 0.0007 2.903e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.097e-09 0 3.1e-09 0.0007 3.103e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.297e-09 0 3.3e-09 0.0007 3.303e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.497e-09 0 3.5e-09 0.0007 3.503e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.697e-09 0 3.7e-09 0.0007 3.703e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.897e-09 0 3.9e-09 0.0007 3.903e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.097e-09 0 4.1e-09 0.0007 4.103e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.297e-09 0 4.3e-09 0.0007 4.303e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.497e-09 0 4.5e-09 0.0007 4.503e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.697e-09 0 4.7e-09 0.0007 4.703e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.897e-09 0 4.9e-09 0.0007 4.903e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.097e-09 0 5.1e-09 0.0007 5.103e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.297e-09 0 5.3e-09 0.0007 5.303e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.497e-09 0 5.5e-09 0.0007 5.503e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.697e-09 0 5.7e-09 0.0007 5.703e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.897e-09 0 5.9e-09 0.0007 5.903e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.097e-09 0 6.1e-09 0.0007 6.103e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.297e-09 0 6.3e-09 0.0007 6.303e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.497e-09 0 6.5e-09 0.0007 6.503e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.697e-09 0 6.7e-09 0.0007 6.703e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.897e-09 0 6.9e-09 0.0007 6.903e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.097e-09 0 7.1e-09 0.0007 7.103e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.297e-09 0 7.3e-09 0.0007 7.303e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.497e-09 0 7.5e-09 0.0007 7.503e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.697e-09 0 7.7e-09 0.0007 7.703e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.897e-09 0 7.9e-09 0.0007 7.903e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.097e-09 0 8.1e-09 0.0007 8.103e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.297e-09 0 8.3e-09 0.0007 8.303e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.497e-09 0 8.5e-09 0.0007 8.503e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.697e-09 0 8.7e-09 0.0007 8.703e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.897e-09 0 8.9e-09 0.0007 8.903e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.097e-09 0 9.1e-09 0.0007 9.103e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.297e-09 0 9.3e-09 0.0007 9.303e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.497e-09 0 9.5e-09 0.0007 9.503e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.697e-09 0 9.7e-09 0.0007 9.703e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.897e-09 0 9.9e-09 0.0007 9.903e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0097e-08 0 1.01e-08 0.0007 1.0103e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0297e-08 0 1.03e-08 0.0007 1.0303e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0497e-08 0 1.05e-08 0.0007 1.0503e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0697e-08 0 1.07e-08 0.0007 1.0703e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0897e-08 0 1.09e-08 0.0007 1.0903e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1097e-08 0 1.11e-08 0.0007 1.1103e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1297e-08 0 1.13e-08 0.0007 1.1303e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1497e-08 0 1.15e-08 0.0007 1.1503e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1697e-08 0 1.17e-08 0.0007 1.1703e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1897e-08 0 1.19e-08 0.0007 1.1903e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2097e-08 0 1.21e-08 0.0007 1.2103e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2297e-08 0 1.23e-08 0.0007 1.2303e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2497e-08 0 1.25e-08 0.0007 1.2503e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2697e-08 0 1.27e-08 0.0007 1.2703e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2897e-08 0 1.29e-08 0.0007 1.2903e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3097e-08 0 1.31e-08 0.0007 1.3103e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3297e-08 0 1.33e-08 0.0007 1.3303e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3497e-08 0 1.35e-08 0.0007 1.3503e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3697e-08 0 1.37e-08 0.0007 1.3703e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3897e-08 0 1.39e-08 0.0007 1.3903e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4097e-08 0 1.41e-08 0.0007 1.4103e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4297e-08 0 1.43e-08 0.0007 1.4303e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4497e-08 0 1.45e-08 0.0007 1.4503e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4697e-08 0 1.47e-08 0.0007 1.4703e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4897e-08 0 1.49e-08 0.0007 1.4903e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5097e-08 0 1.51e-08 0.0007 1.5103e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5297e-08 0 1.53e-08 0.0007 1.5303e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5497e-08 0 1.55e-08 0.0007 1.5503e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5697e-08 0 1.57e-08 0.0007 1.5703e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5897e-08 0 1.59e-08 0.0007 1.5903e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6097e-08 0 1.61e-08 0.0007 1.6103e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6297e-08 0 1.63e-08 0.0007 1.6303e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6497e-08 0 1.65e-08 0.0007 1.6503e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6697e-08 0 1.67e-08 0.0007 1.6703e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7097e-08 0 1.71e-08 0.0007 1.7103e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7297e-08 0 1.73e-08 0.0007 1.7303e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7497e-08 0 1.75e-08 0.0007 1.7503e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7697e-08 0 1.77e-08 0.0007 1.7703e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7897e-08 0 1.79e-08 0.0007 1.7903e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8097e-08 0 1.81e-08 0.0007 1.8103e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8297e-08 0 1.83e-08 0.0007 1.8303e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8497e-08 0 1.85e-08 0.0007 1.8503e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8697e-08 0 1.87e-08 0.0007 1.8703e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8897e-08 0 1.89e-08 0.0007 1.8903e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9097e-08 0 1.91e-08 0.0007 1.9103e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9297e-08 0 1.93e-08 0.0007 1.9303e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9497e-08 0 1.95e-08 0.0007 1.9503e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9697e-08 0 1.97e-08 0.0007 1.9703e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9897e-08 0 1.99e-08 0.0007 1.9903e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0097e-08 0 2.01e-08 0.0007 2.0103e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0297e-08 0 2.03e-08 0.0007 2.0303e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0497e-08 0 2.05e-08 0.0007 2.0503e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0697e-08 0 2.07e-08 0.0007 2.0703e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0897e-08 0 2.09e-08 0.0007 2.0903e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1097e-08 0 2.11e-08 0.0007 2.1103e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1297e-08 0 2.13e-08 0.0007 2.1303e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1497e-08 0 2.15e-08 0.0007 2.1503e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1697e-08 0 2.17e-08 0.0007 2.1703e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1897e-08 0 2.19e-08 0.0007 2.1903e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2097e-08 0 2.21e-08 0.0007 2.2103e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2297e-08 0 2.23e-08 0.0007 2.2303e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2497e-08 0 2.25e-08 0.0007 2.2503e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2697e-08 0 2.27e-08 0.0007 2.2703e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2897e-08 0 2.29e-08 0.0007 2.2903e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3097e-08 0 2.31e-08 0.0007 2.3103e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3297e-08 0 2.33e-08 0.0007 2.3303e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3497e-08 0 2.35e-08 0.0007 2.3503e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3697e-08 0 2.37e-08 0.0007 2.3703e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3897e-08 0 2.39e-08 0.0007 2.3903e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4097e-08 0 2.41e-08 0.0007 2.4103e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4297e-08 0 2.43e-08 0.0007 2.4303e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4497e-08 0 2.45e-08 0.0007 2.4503e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4697e-08 0 2.47e-08 0.0007 2.4703e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4897e-08 0 2.49e-08 0.0007 2.4903e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5097e-08 0 2.51e-08 0.0007 2.5103e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5297e-08 0 2.53e-08 0.0007 2.5303e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5497e-08 0 2.55e-08 0.0007 2.5503e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5697e-08 0 2.57e-08 0.0007 2.5703e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5897e-08 0 2.59e-08 0.0007 2.5903e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6097e-08 0 2.61e-08 0.0007 2.6103e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6297e-08 0 2.63e-08 0.0007 2.6303e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6497e-08 0 2.65e-08 0.0007 2.6503e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6697e-08 0 2.67e-08 0.0007 2.6703e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6897e-08 0 2.69e-08 0.0007 2.6903e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7097e-08 0 2.71e-08 0.0007 2.7103e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7297e-08 0 2.73e-08 0.0007 2.7303e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7497e-08 0 2.75e-08 0.0007 2.7503e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7697e-08 0 2.77e-08 0.0007 2.7703e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7897e-08 0 2.79e-08 0.0007 2.7903e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8097e-08 0 2.81e-08 0.0007 2.8103e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8297e-08 0 2.83e-08 0.0007 2.8303e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8497e-08 0 2.85e-08 0.0007 2.8503e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8697e-08 0 2.87e-08 0.0007 2.8703e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8897e-08 0 2.89e-08 0.0007 2.8903e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9097e-08 0 2.91e-08 0.0007 2.9103e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9297e-08 0 2.93e-08 0.0007 2.9303e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9497e-08 0 2.95e-08 0.0007 2.9503e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9697e-08 0 2.97e-08 0.0007 2.9703e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9897e-08 0 2.99e-08 0.0007 2.9903e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0097e-08 0 3.01e-08 0.0007 3.0103e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0297e-08 0 3.03e-08 0.0007 3.0303e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0497e-08 0 3.05e-08 0.0007 3.0503e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0697e-08 0 3.07e-08 0.0007 3.0703e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0897e-08 0 3.09e-08 0.0007 3.0903e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1097e-08 0 3.11e-08 0.0007 3.1103e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1297e-08 0 3.13e-08 0.0007 3.1303e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1497e-08 0 3.15e-08 0.0007 3.1503e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1697e-08 0 3.17e-08 0.0007 3.1703e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1897e-08 0 3.19e-08 0.0007 3.1903e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2097e-08 0 3.21e-08 0.0007 3.2103e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2297e-08 0 3.23e-08 0.0007 3.2303e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2497e-08 0 3.25e-08 0.0007 3.2503e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2697e-08 0 3.27e-08 0.0007 3.2703e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2897e-08 0 3.29e-08 0.0007 3.2903e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3097e-08 0 3.31e-08 0.0007 3.3103e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3297e-08 0 3.33e-08 0.0007 3.3303e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3497e-08 0 3.35e-08 0.0007 3.3503e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3697e-08 0 3.37e-08 0.0007 3.3703e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3897e-08 0 3.39e-08 0.0007 3.3903e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4097e-08 0 3.41e-08 0.0007 3.4103e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4297e-08 0 3.43e-08 0.0007 3.4303e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4497e-08 0 3.45e-08 0.0007 3.4503e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4697e-08 0 3.47e-08 0.0007 3.4703e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4897e-08 0 3.49e-08 0.0007 3.4903e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5097e-08 0 3.51e-08 0.0007 3.5103e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5297e-08 0 3.53e-08 0.0007 3.5303e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5497e-08 0 3.55e-08 0.0007 3.5503e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5697e-08 0 3.57e-08 0.0007 3.5703e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5897e-08 0 3.59e-08 0.0007 3.5903e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6097e-08 0 3.61e-08 0.0007 3.6103e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6297e-08 0 3.63e-08 0.0007 3.6303e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6497e-08 0 3.65e-08 0.0007 3.6503e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6697e-08 0 3.67e-08 0.0007 3.6703e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6897e-08 0 3.69e-08 0.0007 3.6903e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7097e-08 0 3.71e-08 0.0007 3.7103e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7297e-08 0 3.73e-08 0.0007 3.7303e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7497e-08 0 3.75e-08 0.0007 3.7503e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7697e-08 0 3.77e-08 0.0007 3.7703e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7897e-08 0 3.79e-08 0.0007 3.7903e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8097e-08 0 3.81e-08 0.0007 3.8103e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8297e-08 0 3.83e-08 0.0007 3.8303e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8497e-08 0 3.85e-08 0.0007 3.8503e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8697e-08 0 3.87e-08 0.0007 3.8703e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8897e-08 0 3.89e-08 0.0007 3.8903e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9097e-08 0 3.91e-08 0.0007 3.9103e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9297e-08 0 3.93e-08 0.0007 3.9303e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9497e-08 0 3.95e-08 0.0007 3.9503e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9697e-08 0 3.97e-08 0.0007 3.9703e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9897e-08 0 3.99e-08 0.0007 3.9903e-08 0)
IT2|T 0 CLK2  PWL(0 0 9.7e-11 0 1e-10 0.0007 1.03e-10 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 2.97e-10 0 3e-10 0.0007 3.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 4.97e-10 0 5e-10 0.0007 5.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 6.97e-10 0 7e-10 0.0007 7.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 8.97e-10 0 9e-10 0.0007 9.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.097e-09 0 1.1e-09 0.0007 1.103e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.297e-09 0 1.3e-09 0.0007 1.303e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.497e-09 0 1.5e-09 0.0007 1.503e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.697e-09 0 1.7e-09 0.0007 1.703e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.897e-09 0 1.9e-09 0.0007 1.903e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.097e-09 0 2.1e-09 0.0007 2.103e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.297e-09 0 2.3e-09 0.0007 2.303e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.497e-09 0 2.5e-09 0.0007 2.503e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.697e-09 0 2.7e-09 0.0007 2.703e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.897e-09 0 2.9e-09 0.0007 2.903e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.097e-09 0 3.1e-09 0.0007 3.103e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.297e-09 0 3.3e-09 0.0007 3.303e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.497e-09 0 3.5e-09 0.0007 3.503e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.697e-09 0 3.7e-09 0.0007 3.703e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.897e-09 0 3.9e-09 0.0007 3.903e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.097e-09 0 4.1e-09 0.0007 4.103e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.297e-09 0 4.3e-09 0.0007 4.303e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.497e-09 0 4.5e-09 0.0007 4.503e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.697e-09 0 4.7e-09 0.0007 4.703e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.897e-09 0 4.9e-09 0.0007 4.903e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.097e-09 0 5.1e-09 0.0007 5.103e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.297e-09 0 5.3e-09 0.0007 5.303e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.497e-09 0 5.5e-09 0.0007 5.503e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.697e-09 0 5.7e-09 0.0007 5.703e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.897e-09 0 5.9e-09 0.0007 5.903e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.097e-09 0 6.1e-09 0.0007 6.103e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.297e-09 0 6.3e-09 0.0007 6.303e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.497e-09 0 6.5e-09 0.0007 6.503e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.697e-09 0 6.7e-09 0.0007 6.703e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.897e-09 0 6.9e-09 0.0007 6.903e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.097e-09 0 7.1e-09 0.0007 7.103e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.297e-09 0 7.3e-09 0.0007 7.303e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.497e-09 0 7.5e-09 0.0007 7.503e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.697e-09 0 7.7e-09 0.0007 7.703e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.897e-09 0 7.9e-09 0.0007 7.903e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.097e-09 0 8.1e-09 0.0007 8.103e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.297e-09 0 8.3e-09 0.0007 8.303e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.497e-09 0 8.5e-09 0.0007 8.503e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.697e-09 0 8.7e-09 0.0007 8.703e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.897e-09 0 8.9e-09 0.0007 8.903e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.097e-09 0 9.1e-09 0.0007 9.103e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.297e-09 0 9.3e-09 0.0007 9.303e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.497e-09 0 9.5e-09 0.0007 9.503e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.697e-09 0 9.7e-09 0.0007 9.703e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.897e-09 0 9.9e-09 0.0007 9.903e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0097e-08 0 1.01e-08 0.0007 1.0103e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0297e-08 0 1.03e-08 0.0007 1.0303e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0497e-08 0 1.05e-08 0.0007 1.0503e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0697e-08 0 1.07e-08 0.0007 1.0703e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0897e-08 0 1.09e-08 0.0007 1.0903e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1097e-08 0 1.11e-08 0.0007 1.1103e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1297e-08 0 1.13e-08 0.0007 1.1303e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1497e-08 0 1.15e-08 0.0007 1.1503e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1697e-08 0 1.17e-08 0.0007 1.1703e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1897e-08 0 1.19e-08 0.0007 1.1903e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2097e-08 0 1.21e-08 0.0007 1.2103e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2297e-08 0 1.23e-08 0.0007 1.2303e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2497e-08 0 1.25e-08 0.0007 1.2503e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2697e-08 0 1.27e-08 0.0007 1.2703e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2897e-08 0 1.29e-08 0.0007 1.2903e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3097e-08 0 1.31e-08 0.0007 1.3103e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3297e-08 0 1.33e-08 0.0007 1.3303e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3497e-08 0 1.35e-08 0.0007 1.3503e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3697e-08 0 1.37e-08 0.0007 1.3703e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3897e-08 0 1.39e-08 0.0007 1.3903e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4097e-08 0 1.41e-08 0.0007 1.4103e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4297e-08 0 1.43e-08 0.0007 1.4303e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4497e-08 0 1.45e-08 0.0007 1.4503e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4697e-08 0 1.47e-08 0.0007 1.4703e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4897e-08 0 1.49e-08 0.0007 1.4903e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5097e-08 0 1.51e-08 0.0007 1.5103e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5297e-08 0 1.53e-08 0.0007 1.5303e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5497e-08 0 1.55e-08 0.0007 1.5503e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5697e-08 0 1.57e-08 0.0007 1.5703e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5897e-08 0 1.59e-08 0.0007 1.5903e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6097e-08 0 1.61e-08 0.0007 1.6103e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6297e-08 0 1.63e-08 0.0007 1.6303e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6497e-08 0 1.65e-08 0.0007 1.6503e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6697e-08 0 1.67e-08 0.0007 1.6703e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7097e-08 0 1.71e-08 0.0007 1.7103e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7297e-08 0 1.73e-08 0.0007 1.7303e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7497e-08 0 1.75e-08 0.0007 1.7503e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7697e-08 0 1.77e-08 0.0007 1.7703e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7897e-08 0 1.79e-08 0.0007 1.7903e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8097e-08 0 1.81e-08 0.0007 1.8103e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8297e-08 0 1.83e-08 0.0007 1.8303e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8497e-08 0 1.85e-08 0.0007 1.8503e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8697e-08 0 1.87e-08 0.0007 1.8703e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8897e-08 0 1.89e-08 0.0007 1.8903e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9097e-08 0 1.91e-08 0.0007 1.9103e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9297e-08 0 1.93e-08 0.0007 1.9303e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9497e-08 0 1.95e-08 0.0007 1.9503e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9697e-08 0 1.97e-08 0.0007 1.9703e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9897e-08 0 1.99e-08 0.0007 1.9903e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0097e-08 0 2.01e-08 0.0007 2.0103e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0297e-08 0 2.03e-08 0.0007 2.0303e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0497e-08 0 2.05e-08 0.0007 2.0503e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0697e-08 0 2.07e-08 0.0007 2.0703e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0897e-08 0 2.09e-08 0.0007 2.0903e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1097e-08 0 2.11e-08 0.0007 2.1103e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1297e-08 0 2.13e-08 0.0007 2.1303e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1497e-08 0 2.15e-08 0.0007 2.1503e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1697e-08 0 2.17e-08 0.0007 2.1703e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1897e-08 0 2.19e-08 0.0007 2.1903e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2097e-08 0 2.21e-08 0.0007 2.2103e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2297e-08 0 2.23e-08 0.0007 2.2303e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2497e-08 0 2.25e-08 0.0007 2.2503e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2697e-08 0 2.27e-08 0.0007 2.2703e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2897e-08 0 2.29e-08 0.0007 2.2903e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3097e-08 0 2.31e-08 0.0007 2.3103e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3297e-08 0 2.33e-08 0.0007 2.3303e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3497e-08 0 2.35e-08 0.0007 2.3503e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3697e-08 0 2.37e-08 0.0007 2.3703e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3897e-08 0 2.39e-08 0.0007 2.3903e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4097e-08 0 2.41e-08 0.0007 2.4103e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4297e-08 0 2.43e-08 0.0007 2.4303e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4497e-08 0 2.45e-08 0.0007 2.4503e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4697e-08 0 2.47e-08 0.0007 2.4703e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4897e-08 0 2.49e-08 0.0007 2.4903e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5097e-08 0 2.51e-08 0.0007 2.5103e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5297e-08 0 2.53e-08 0.0007 2.5303e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5497e-08 0 2.55e-08 0.0007 2.5503e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5697e-08 0 2.57e-08 0.0007 2.5703e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5897e-08 0 2.59e-08 0.0007 2.5903e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6097e-08 0 2.61e-08 0.0007 2.6103e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6297e-08 0 2.63e-08 0.0007 2.6303e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6497e-08 0 2.65e-08 0.0007 2.6503e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6697e-08 0 2.67e-08 0.0007 2.6703e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6897e-08 0 2.69e-08 0.0007 2.6903e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7097e-08 0 2.71e-08 0.0007 2.7103e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7297e-08 0 2.73e-08 0.0007 2.7303e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7497e-08 0 2.75e-08 0.0007 2.7503e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7697e-08 0 2.77e-08 0.0007 2.7703e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7897e-08 0 2.79e-08 0.0007 2.7903e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8097e-08 0 2.81e-08 0.0007 2.8103e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8297e-08 0 2.83e-08 0.0007 2.8303e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8497e-08 0 2.85e-08 0.0007 2.8503e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8697e-08 0 2.87e-08 0.0007 2.8703e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8897e-08 0 2.89e-08 0.0007 2.8903e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9097e-08 0 2.91e-08 0.0007 2.9103e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9297e-08 0 2.93e-08 0.0007 2.9303e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9497e-08 0 2.95e-08 0.0007 2.9503e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9697e-08 0 2.97e-08 0.0007 2.9703e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9897e-08 0 2.99e-08 0.0007 2.9903e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0097e-08 0 3.01e-08 0.0007 3.0103e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0297e-08 0 3.03e-08 0.0007 3.0303e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0497e-08 0 3.05e-08 0.0007 3.0503e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0697e-08 0 3.07e-08 0.0007 3.0703e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0897e-08 0 3.09e-08 0.0007 3.0903e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1097e-08 0 3.11e-08 0.0007 3.1103e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1297e-08 0 3.13e-08 0.0007 3.1303e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1497e-08 0 3.15e-08 0.0007 3.1503e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1697e-08 0 3.17e-08 0.0007 3.1703e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1897e-08 0 3.19e-08 0.0007 3.1903e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2097e-08 0 3.21e-08 0.0007 3.2103e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2297e-08 0 3.23e-08 0.0007 3.2303e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2497e-08 0 3.25e-08 0.0007 3.2503e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2697e-08 0 3.27e-08 0.0007 3.2703e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2897e-08 0 3.29e-08 0.0007 3.2903e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3097e-08 0 3.31e-08 0.0007 3.3103e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3297e-08 0 3.33e-08 0.0007 3.3303e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3497e-08 0 3.35e-08 0.0007 3.3503e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3697e-08 0 3.37e-08 0.0007 3.3703e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3897e-08 0 3.39e-08 0.0007 3.3903e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4097e-08 0 3.41e-08 0.0007 3.4103e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4297e-08 0 3.43e-08 0.0007 3.4303e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4497e-08 0 3.45e-08 0.0007 3.4503e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4697e-08 0 3.47e-08 0.0007 3.4703e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4897e-08 0 3.49e-08 0.0007 3.4903e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5097e-08 0 3.51e-08 0.0007 3.5103e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5297e-08 0 3.53e-08 0.0007 3.5303e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5497e-08 0 3.55e-08 0.0007 3.5503e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5697e-08 0 3.57e-08 0.0007 3.5703e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5897e-08 0 3.59e-08 0.0007 3.5903e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6097e-08 0 3.61e-08 0.0007 3.6103e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6297e-08 0 3.63e-08 0.0007 3.6303e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6497e-08 0 3.65e-08 0.0007 3.6503e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6697e-08 0 3.67e-08 0.0007 3.6703e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6897e-08 0 3.69e-08 0.0007 3.6903e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7097e-08 0 3.71e-08 0.0007 3.7103e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7297e-08 0 3.73e-08 0.0007 3.7303e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7497e-08 0 3.75e-08 0.0007 3.7503e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7697e-08 0 3.77e-08 0.0007 3.7703e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7897e-08 0 3.79e-08 0.0007 3.7903e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8097e-08 0 3.81e-08 0.0007 3.8103e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8297e-08 0 3.83e-08 0.0007 3.8303e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8497e-08 0 3.85e-08 0.0007 3.8503e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8697e-08 0 3.87e-08 0.0007 3.8703e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8897e-08 0 3.89e-08 0.0007 3.8903e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9097e-08 0 3.91e-08 0.0007 3.9103e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9297e-08 0 3.93e-08 0.0007 3.9303e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9497e-08 0 3.95e-08 0.0007 3.9503e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9697e-08 0 3.97e-08 0.0007 3.9703e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9897e-08 0 3.99e-08 0.0007 3.9903e-08 0)
IT3|T 0 CLK3  PWL(0 0 9.7e-11 0 1e-10 0.0007 1.03e-10 0 1.97e-10 0 2e-10 0.0007 2.03e-10 0 2.97e-10 0 3e-10 0.0007 3.03e-10 0 3.97e-10 0 4e-10 0.0007 4.03e-10 0 4.97e-10 0 5e-10 0.0007 5.03e-10 0 5.97e-10 0 6e-10 0.0007 6.03e-10 0 6.97e-10 0 7e-10 0.0007 7.03e-10 0 7.97e-10 0 8e-10 0.0007 8.03e-10 0 8.97e-10 0 9e-10 0.0007 9.03e-10 0 9.97e-10 0 1e-09 0.0007 1.003e-09 0 1.097e-09 0 1.1e-09 0.0007 1.103e-09 0 1.197e-09 0 1.2e-09 0.0007 1.203e-09 0 1.297e-09 0 1.3e-09 0.0007 1.303e-09 0 1.397e-09 0 1.4e-09 0.0007 1.403e-09 0 1.497e-09 0 1.5e-09 0.0007 1.503e-09 0 1.597e-09 0 1.6e-09 0.0007 1.603e-09 0 1.697e-09 0 1.7e-09 0.0007 1.703e-09 0 1.797e-09 0 1.8e-09 0.0007 1.803e-09 0 1.897e-09 0 1.9e-09 0.0007 1.903e-09 0 1.997e-09 0 2e-09 0.0007 2.003e-09 0 2.097e-09 0 2.1e-09 0.0007 2.103e-09 0 2.197e-09 0 2.2e-09 0.0007 2.203e-09 0 2.297e-09 0 2.3e-09 0.0007 2.303e-09 0 2.397e-09 0 2.4e-09 0.0007 2.403e-09 0 2.497e-09 0 2.5e-09 0.0007 2.503e-09 0 2.597e-09 0 2.6e-09 0.0007 2.603e-09 0 2.697e-09 0 2.7e-09 0.0007 2.703e-09 0 2.797e-09 0 2.8e-09 0.0007 2.803e-09 0 2.897e-09 0 2.9e-09 0.0007 2.903e-09 0 2.997e-09 0 3e-09 0.0007 3.003e-09 0 3.097e-09 0 3.1e-09 0.0007 3.103e-09 0 3.197e-09 0 3.2e-09 0.0007 3.203e-09 0 3.297e-09 0 3.3e-09 0.0007 3.303e-09 0 3.397e-09 0 3.4e-09 0.0007 3.403e-09 0 3.497e-09 0 3.5e-09 0.0007 3.503e-09 0 3.597e-09 0 3.6e-09 0.0007 3.603e-09 0 3.697e-09 0 3.7e-09 0.0007 3.703e-09 0 3.797e-09 0 3.8e-09 0.0007 3.803e-09 0 3.897e-09 0 3.9e-09 0.0007 3.903e-09 0 3.997e-09 0 4e-09 0.0007 4.003e-09 0 4.097e-09 0 4.1e-09 0.0007 4.103e-09 0 4.197e-09 0 4.2e-09 0.0007 4.203e-09 0 4.297e-09 0 4.3e-09 0.0007 4.303e-09 0 4.397e-09 0 4.4e-09 0.0007 4.403e-09 0 4.497e-09 0 4.5e-09 0.0007 4.503e-09 0 4.597e-09 0 4.6e-09 0.0007 4.603e-09 0 4.697e-09 0 4.7e-09 0.0007 4.703e-09 0 4.797e-09 0 4.8e-09 0.0007 4.803e-09 0 4.897e-09 0 4.9e-09 0.0007 4.903e-09 0 4.997e-09 0 5e-09 0.0007 5.003e-09 0 5.097e-09 0 5.1e-09 0.0007 5.103e-09 0 5.197e-09 0 5.2e-09 0.0007 5.203e-09 0 5.297e-09 0 5.3e-09 0.0007 5.303e-09 0 5.397e-09 0 5.4e-09 0.0007 5.403e-09 0 5.497e-09 0 5.5e-09 0.0007 5.503e-09 0 5.597e-09 0 5.6e-09 0.0007 5.603e-09 0 5.697e-09 0 5.7e-09 0.0007 5.703e-09 0 5.797e-09 0 5.8e-09 0.0007 5.803e-09 0 5.897e-09 0 5.9e-09 0.0007 5.903e-09 0 5.997e-09 0 6e-09 0.0007 6.003e-09 0 6.097e-09 0 6.1e-09 0.0007 6.103e-09 0 6.197e-09 0 6.2e-09 0.0007 6.203e-09 0 6.297e-09 0 6.3e-09 0.0007 6.303e-09 0 6.397e-09 0 6.4e-09 0.0007 6.403e-09 0 6.497e-09 0 6.5e-09 0.0007 6.503e-09 0 6.597e-09 0 6.6e-09 0.0007 6.603e-09 0 6.697e-09 0 6.7e-09 0.0007 6.703e-09 0 6.797e-09 0 6.8e-09 0.0007 6.803e-09 0 6.897e-09 0 6.9e-09 0.0007 6.903e-09 0 6.997e-09 0 7e-09 0.0007 7.003e-09 0 7.097e-09 0 7.1e-09 0.0007 7.103e-09 0 7.197e-09 0 7.2e-09 0.0007 7.203e-09 0 7.297e-09 0 7.3e-09 0.0007 7.303e-09 0 7.397e-09 0 7.4e-09 0.0007 7.403e-09 0 7.497e-09 0 7.5e-09 0.0007 7.503e-09 0 7.597e-09 0 7.6e-09 0.0007 7.603e-09 0 7.697e-09 0 7.7e-09 0.0007 7.703e-09 0 7.797e-09 0 7.8e-09 0.0007 7.803e-09 0 7.897e-09 0 7.9e-09 0.0007 7.903e-09 0 7.997e-09 0 8e-09 0.0007 8.003e-09 0 8.097e-09 0 8.1e-09 0.0007 8.103e-09 0 8.197e-09 0 8.2e-09 0.0007 8.203e-09 0 8.297e-09 0 8.3e-09 0.0007 8.303e-09 0 8.397e-09 0 8.4e-09 0.0007 8.403e-09 0 8.497e-09 0 8.5e-09 0.0007 8.503e-09 0 8.597e-09 0 8.6e-09 0.0007 8.603e-09 0 8.697e-09 0 8.7e-09 0.0007 8.703e-09 0 8.797e-09 0 8.8e-09 0.0007 8.803e-09 0 8.897e-09 0 8.9e-09 0.0007 8.903e-09 0 8.997e-09 0 9e-09 0.0007 9.003e-09 0 9.097e-09 0 9.1e-09 0.0007 9.103e-09 0 9.197e-09 0 9.2e-09 0.0007 9.203e-09 0 9.297e-09 0 9.3e-09 0.0007 9.303e-09 0 9.397e-09 0 9.4e-09 0.0007 9.403e-09 0 9.497e-09 0 9.5e-09 0.0007 9.503e-09 0 9.597e-09 0 9.6e-09 0.0007 9.603e-09 0 9.697e-09 0 9.7e-09 0.0007 9.703e-09 0 9.797e-09 0 9.8e-09 0.0007 9.803e-09 0 9.897e-09 0 9.9e-09 0.0007 9.903e-09 0 9.997e-09 0 1e-08 0.0007 1.0003e-08 0 1.0097e-08 0 1.01e-08 0.0007 1.0103e-08 0 1.0197e-08 0 1.02e-08 0.0007 1.0203e-08 0 1.0297e-08 0 1.03e-08 0.0007 1.0303e-08 0 1.0397e-08 0 1.04e-08 0.0007 1.0403e-08 0 1.0497e-08 0 1.05e-08 0.0007 1.0503e-08 0 1.0597e-08 0 1.06e-08 0.0007 1.0603e-08 0 1.0697e-08 0 1.07e-08 0.0007 1.0703e-08 0 1.0797e-08 0 1.08e-08 0.0007 1.0803e-08 0 1.0897e-08 0 1.09e-08 0.0007 1.0903e-08 0 1.0997e-08 0 1.1e-08 0.0007 1.1003e-08 0 1.1097e-08 0 1.11e-08 0.0007 1.1103e-08 0 1.1197e-08 0 1.12e-08 0.0007 1.1203e-08 0 1.1297e-08 0 1.13e-08 0.0007 1.1303e-08 0 1.1397e-08 0 1.14e-08 0.0007 1.1403e-08 0 1.1497e-08 0 1.15e-08 0.0007 1.1503e-08 0 1.1597e-08 0 1.16e-08 0.0007 1.1603e-08 0 1.1697e-08 0 1.17e-08 0.0007 1.1703e-08 0 1.1797e-08 0 1.18e-08 0.0007 1.1803e-08 0 1.1897e-08 0 1.19e-08 0.0007 1.1903e-08 0 1.1997e-08 0 1.2e-08 0.0007 1.2003e-08 0 1.2097e-08 0 1.21e-08 0.0007 1.2103e-08 0 1.2197e-08 0 1.22e-08 0.0007 1.2203e-08 0 1.2297e-08 0 1.23e-08 0.0007 1.2303e-08 0 1.2397e-08 0 1.24e-08 0.0007 1.2403e-08 0 1.2497e-08 0 1.25e-08 0.0007 1.2503e-08 0 1.2597e-08 0 1.26e-08 0.0007 1.2603e-08 0 1.2697e-08 0 1.27e-08 0.0007 1.2703e-08 0 1.2797e-08 0 1.28e-08 0.0007 1.2803e-08 0 1.2897e-08 0 1.29e-08 0.0007 1.2903e-08 0 1.2997e-08 0 1.3e-08 0.0007 1.3003e-08 0 1.3097e-08 0 1.31e-08 0.0007 1.3103e-08 0 1.3197e-08 0 1.32e-08 0.0007 1.3203e-08 0 1.3297e-08 0 1.33e-08 0.0007 1.3303e-08 0 1.3397e-08 0 1.34e-08 0.0007 1.3403e-08 0 1.3497e-08 0 1.35e-08 0.0007 1.3503e-08 0 1.3597e-08 0 1.36e-08 0.0007 1.3603e-08 0 1.3697e-08 0 1.37e-08 0.0007 1.3703e-08 0 1.3797e-08 0 1.38e-08 0.0007 1.3803e-08 0 1.3897e-08 0 1.39e-08 0.0007 1.3903e-08 0 1.3997e-08 0 1.4e-08 0.0007 1.4003e-08 0 1.4097e-08 0 1.41e-08 0.0007 1.4103e-08 0 1.4197e-08 0 1.42e-08 0.0007 1.4203e-08 0 1.4297e-08 0 1.43e-08 0.0007 1.4303e-08 0 1.4397e-08 0 1.44e-08 0.0007 1.4403e-08 0 1.4497e-08 0 1.45e-08 0.0007 1.4503e-08 0 1.4597e-08 0 1.46e-08 0.0007 1.4603e-08 0 1.4697e-08 0 1.47e-08 0.0007 1.4703e-08 0 1.4797e-08 0 1.48e-08 0.0007 1.4803e-08 0 1.4897e-08 0 1.49e-08 0.0007 1.4903e-08 0 1.4997e-08 0 1.5e-08 0.0007 1.5003e-08 0 1.5097e-08 0 1.51e-08 0.0007 1.5103e-08 0 1.5197e-08 0 1.52e-08 0.0007 1.5203e-08 0 1.5297e-08 0 1.53e-08 0.0007 1.5303e-08 0 1.5397e-08 0 1.54e-08 0.0007 1.5403e-08 0 1.5497e-08 0 1.55e-08 0.0007 1.5503e-08 0 1.5597e-08 0 1.56e-08 0.0007 1.5603e-08 0 1.5697e-08 0 1.57e-08 0.0007 1.5703e-08 0 1.5797e-08 0 1.58e-08 0.0007 1.5803e-08 0 1.5897e-08 0 1.59e-08 0.0007 1.5903e-08 0 1.5997e-08 0 1.6e-08 0.0007 1.6003e-08 0 1.6097e-08 0 1.61e-08 0.0007 1.6103e-08 0 1.6197e-08 0 1.62e-08 0.0007 1.6203e-08 0 1.6297e-08 0 1.63e-08 0.0007 1.6303e-08 0 1.6397e-08 0 1.64e-08 0.0007 1.6403e-08 0 1.6497e-08 0 1.65e-08 0.0007 1.6503e-08 0 1.6597e-08 0 1.66e-08 0.0007 1.6603e-08 0 1.6697e-08 0 1.67e-08 0.0007 1.6703e-08 0 1.6797e-08 0 1.68e-08 0.0007 1.6803e-08 0 1.6897e-08 0 1.69e-08 0.0007 1.6903e-08 0 1.6997e-08 0 1.7e-08 0.0007 1.7003e-08 0 1.7097e-08 0 1.71e-08 0.0007 1.7103e-08 0 1.7197e-08 0 1.72e-08 0.0007 1.7203e-08 0 1.7297e-08 0 1.73e-08 0.0007 1.7303e-08 0 1.7397e-08 0 1.74e-08 0.0007 1.7403e-08 0 1.7497e-08 0 1.75e-08 0.0007 1.7503e-08 0 1.7597e-08 0 1.76e-08 0.0007 1.7603e-08 0 1.7697e-08 0 1.77e-08 0.0007 1.7703e-08 0 1.7797e-08 0 1.78e-08 0.0007 1.7803e-08 0 1.7897e-08 0 1.79e-08 0.0007 1.7903e-08 0 1.7997e-08 0 1.8e-08 0.0007 1.8003e-08 0 1.8097e-08 0 1.81e-08 0.0007 1.8103e-08 0 1.8197e-08 0 1.82e-08 0.0007 1.8203e-08 0 1.8297e-08 0 1.83e-08 0.0007 1.8303e-08 0 1.8397e-08 0 1.84e-08 0.0007 1.8403e-08 0 1.8497e-08 0 1.85e-08 0.0007 1.8503e-08 0 1.8597e-08 0 1.86e-08 0.0007 1.8603e-08 0 1.8697e-08 0 1.87e-08 0.0007 1.8703e-08 0 1.8797e-08 0 1.88e-08 0.0007 1.8803e-08 0 1.8897e-08 0 1.89e-08 0.0007 1.8903e-08 0 1.8997e-08 0 1.9e-08 0.0007 1.9003e-08 0 1.9097e-08 0 1.91e-08 0.0007 1.9103e-08 0 1.9197e-08 0 1.92e-08 0.0007 1.9203e-08 0 1.9297e-08 0 1.93e-08 0.0007 1.9303e-08 0 1.9397e-08 0 1.94e-08 0.0007 1.9403e-08 0 1.9497e-08 0 1.95e-08 0.0007 1.9503e-08 0 1.9597e-08 0 1.96e-08 0.0007 1.9603e-08 0 1.9697e-08 0 1.97e-08 0.0007 1.9703e-08 0 1.9797e-08 0 1.98e-08 0.0007 1.9803e-08 0 1.9897e-08 0 1.99e-08 0.0007 1.9903e-08 0 1.9997e-08 0 2e-08 0.0007 2.0003e-08 0 2.0097e-08 0 2.01e-08 0.0007 2.0103e-08 0 2.0197e-08 0 2.02e-08 0.0007 2.0203e-08 0 2.0297e-08 0 2.03e-08 0.0007 2.0303e-08 0 2.0397e-08 0 2.04e-08 0.0007 2.0403e-08 0 2.0497e-08 0 2.05e-08 0.0007 2.0503e-08 0 2.0597e-08 0 2.06e-08 0.0007 2.0603e-08 0 2.0697e-08 0 2.07e-08 0.0007 2.0703e-08 0 2.0797e-08 0 2.08e-08 0.0007 2.0803e-08 0 2.0897e-08 0 2.09e-08 0.0007 2.0903e-08 0 2.0997e-08 0 2.1e-08 0.0007 2.1003e-08 0 2.1097e-08 0 2.11e-08 0.0007 2.1103e-08 0 2.1197e-08 0 2.12e-08 0.0007 2.1203e-08 0 2.1297e-08 0 2.13e-08 0.0007 2.1303e-08 0 2.1397e-08 0 2.14e-08 0.0007 2.1403e-08 0 2.1497e-08 0 2.15e-08 0.0007 2.1503e-08 0 2.1597e-08 0 2.16e-08 0.0007 2.1603e-08 0 2.1697e-08 0 2.17e-08 0.0007 2.1703e-08 0 2.1797e-08 0 2.18e-08 0.0007 2.1803e-08 0 2.1897e-08 0 2.19e-08 0.0007 2.1903e-08 0 2.1997e-08 0 2.2e-08 0.0007 2.2003e-08 0 2.2097e-08 0 2.21e-08 0.0007 2.2103e-08 0 2.2197e-08 0 2.22e-08 0.0007 2.2203e-08 0 2.2297e-08 0 2.23e-08 0.0007 2.2303e-08 0 2.2397e-08 0 2.24e-08 0.0007 2.2403e-08 0 2.2497e-08 0 2.25e-08 0.0007 2.2503e-08 0 2.2597e-08 0 2.26e-08 0.0007 2.2603e-08 0 2.2697e-08 0 2.27e-08 0.0007 2.2703e-08 0 2.2797e-08 0 2.28e-08 0.0007 2.2803e-08 0 2.2897e-08 0 2.29e-08 0.0007 2.2903e-08 0 2.2997e-08 0 2.3e-08 0.0007 2.3003e-08 0 2.3097e-08 0 2.31e-08 0.0007 2.3103e-08 0 2.3197e-08 0 2.32e-08 0.0007 2.3203e-08 0 2.3297e-08 0 2.33e-08 0.0007 2.3303e-08 0 2.3397e-08 0 2.34e-08 0.0007 2.3403e-08 0 2.3497e-08 0 2.35e-08 0.0007 2.3503e-08 0 2.3597e-08 0 2.36e-08 0.0007 2.3603e-08 0 2.3697e-08 0 2.37e-08 0.0007 2.3703e-08 0 2.3797e-08 0 2.38e-08 0.0007 2.3803e-08 0 2.3897e-08 0 2.39e-08 0.0007 2.3903e-08 0 2.3997e-08 0 2.4e-08 0.0007 2.4003e-08 0 2.4097e-08 0 2.41e-08 0.0007 2.4103e-08 0 2.4197e-08 0 2.42e-08 0.0007 2.4203e-08 0 2.4297e-08 0 2.43e-08 0.0007 2.4303e-08 0 2.4397e-08 0 2.44e-08 0.0007 2.4403e-08 0 2.4497e-08 0 2.45e-08 0.0007 2.4503e-08 0 2.4597e-08 0 2.46e-08 0.0007 2.4603e-08 0 2.4697e-08 0 2.47e-08 0.0007 2.4703e-08 0 2.4797e-08 0 2.48e-08 0.0007 2.4803e-08 0 2.4897e-08 0 2.49e-08 0.0007 2.4903e-08 0 2.4997e-08 0 2.5e-08 0.0007 2.5003e-08 0 2.5097e-08 0 2.51e-08 0.0007 2.5103e-08 0 2.5197e-08 0 2.52e-08 0.0007 2.5203e-08 0 2.5297e-08 0 2.53e-08 0.0007 2.5303e-08 0 2.5397e-08 0 2.54e-08 0.0007 2.5403e-08 0 2.5497e-08 0 2.55e-08 0.0007 2.5503e-08 0 2.5597e-08 0 2.56e-08 0.0007 2.5603e-08 0 2.5697e-08 0 2.57e-08 0.0007 2.5703e-08 0 2.5797e-08 0 2.58e-08 0.0007 2.5803e-08 0 2.5897e-08 0 2.59e-08 0.0007 2.5903e-08 0 2.5997e-08 0 2.6e-08 0.0007 2.6003e-08 0 2.6097e-08 0 2.61e-08 0.0007 2.6103e-08 0 2.6197e-08 0 2.62e-08 0.0007 2.6203e-08 0 2.6297e-08 0 2.63e-08 0.0007 2.6303e-08 0 2.6397e-08 0 2.64e-08 0.0007 2.6403e-08 0 2.6497e-08 0 2.65e-08 0.0007 2.6503e-08 0 2.6597e-08 0 2.66e-08 0.0007 2.6603e-08 0 2.6697e-08 0 2.67e-08 0.0007 2.6703e-08 0 2.6797e-08 0 2.68e-08 0.0007 2.6803e-08 0 2.6897e-08 0 2.69e-08 0.0007 2.6903e-08 0 2.6997e-08 0 2.7e-08 0.0007 2.7003e-08 0 2.7097e-08 0 2.71e-08 0.0007 2.7103e-08 0 2.7197e-08 0 2.72e-08 0.0007 2.7203e-08 0 2.7297e-08 0 2.73e-08 0.0007 2.7303e-08 0 2.7397e-08 0 2.74e-08 0.0007 2.7403e-08 0 2.7497e-08 0 2.75e-08 0.0007 2.7503e-08 0 2.7597e-08 0 2.76e-08 0.0007 2.7603e-08 0 2.7697e-08 0 2.77e-08 0.0007 2.7703e-08 0 2.7797e-08 0 2.78e-08 0.0007 2.7803e-08 0 2.7897e-08 0 2.79e-08 0.0007 2.7903e-08 0 2.7997e-08 0 2.8e-08 0.0007 2.8003e-08 0 2.8097e-08 0 2.81e-08 0.0007 2.8103e-08 0 2.8197e-08 0 2.82e-08 0.0007 2.8203e-08 0 2.8297e-08 0 2.83e-08 0.0007 2.8303e-08 0 2.8397e-08 0 2.84e-08 0.0007 2.8403e-08 0 2.8497e-08 0 2.85e-08 0.0007 2.8503e-08 0 2.8597e-08 0 2.86e-08 0.0007 2.8603e-08 0 2.8697e-08 0 2.87e-08 0.0007 2.8703e-08 0 2.8797e-08 0 2.88e-08 0.0007 2.8803e-08 0 2.8897e-08 0 2.89e-08 0.0007 2.8903e-08 0 2.8997e-08 0 2.9e-08 0.0007 2.9003e-08 0 2.9097e-08 0 2.91e-08 0.0007 2.9103e-08 0 2.9197e-08 0 2.92e-08 0.0007 2.9203e-08 0 2.9297e-08 0 2.93e-08 0.0007 2.9303e-08 0 2.9397e-08 0 2.94e-08 0.0007 2.9403e-08 0 2.9497e-08 0 2.95e-08 0.0007 2.9503e-08 0 2.9597e-08 0 2.96e-08 0.0007 2.9603e-08 0 2.9697e-08 0 2.97e-08 0.0007 2.9703e-08 0 2.9797e-08 0 2.98e-08 0.0007 2.9803e-08 0 2.9897e-08 0 2.99e-08 0.0007 2.9903e-08 0 2.9997e-08 0 3e-08 0.0007 3.0003e-08 0 3.0097e-08 0 3.01e-08 0.0007 3.0103e-08 0 3.0197e-08 0 3.02e-08 0.0007 3.0203e-08 0 3.0297e-08 0 3.03e-08 0.0007 3.0303e-08 0 3.0397e-08 0 3.04e-08 0.0007 3.0403e-08 0 3.0497e-08 0 3.05e-08 0.0007 3.0503e-08 0 3.0597e-08 0 3.06e-08 0.0007 3.0603e-08 0 3.0697e-08 0 3.07e-08 0.0007 3.0703e-08 0 3.0797e-08 0 3.08e-08 0.0007 3.0803e-08 0 3.0897e-08 0 3.09e-08 0.0007 3.0903e-08 0 3.0997e-08 0 3.1e-08 0.0007 3.1003e-08 0 3.1097e-08 0 3.11e-08 0.0007 3.1103e-08 0 3.1197e-08 0 3.12e-08 0.0007 3.1203e-08 0 3.1297e-08 0 3.13e-08 0.0007 3.1303e-08 0 3.1397e-08 0 3.14e-08 0.0007 3.1403e-08 0 3.1497e-08 0 3.15e-08 0.0007 3.1503e-08 0 3.1597e-08 0 3.16e-08 0.0007 3.1603e-08 0 3.1697e-08 0 3.17e-08 0.0007 3.1703e-08 0 3.1797e-08 0 3.18e-08 0.0007 3.1803e-08 0 3.1897e-08 0 3.19e-08 0.0007 3.1903e-08 0 3.1997e-08 0 3.2e-08 0.0007 3.2003e-08 0 3.2097e-08 0 3.21e-08 0.0007 3.2103e-08 0 3.2197e-08 0 3.22e-08 0.0007 3.2203e-08 0 3.2297e-08 0 3.23e-08 0.0007 3.2303e-08 0 3.2397e-08 0 3.24e-08 0.0007 3.2403e-08 0 3.2497e-08 0 3.25e-08 0.0007 3.2503e-08 0 3.2597e-08 0 3.26e-08 0.0007 3.2603e-08 0 3.2697e-08 0 3.27e-08 0.0007 3.2703e-08 0 3.2797e-08 0 3.28e-08 0.0007 3.2803e-08 0 3.2897e-08 0 3.29e-08 0.0007 3.2903e-08 0 3.2997e-08 0 3.3e-08 0.0007 3.3003e-08 0 3.3097e-08 0 3.31e-08 0.0007 3.3103e-08 0 3.3197e-08 0 3.32e-08 0.0007 3.3203e-08 0 3.3297e-08 0 3.33e-08 0.0007 3.3303e-08 0 3.3397e-08 0 3.34e-08 0.0007 3.3403e-08 0 3.3497e-08 0 3.35e-08 0.0007 3.3503e-08 0 3.3597e-08 0 3.36e-08 0.0007 3.3603e-08 0 3.3697e-08 0 3.37e-08 0.0007 3.3703e-08 0 3.3797e-08 0 3.38e-08 0.0007 3.3803e-08 0 3.3897e-08 0 3.39e-08 0.0007 3.3903e-08 0 3.3997e-08 0 3.4e-08 0.0007 3.4003e-08 0 3.4097e-08 0 3.41e-08 0.0007 3.4103e-08 0 3.4197e-08 0 3.42e-08 0.0007 3.4203e-08 0 3.4297e-08 0 3.43e-08 0.0007 3.4303e-08 0 3.4397e-08 0 3.44e-08 0.0007 3.4403e-08 0 3.4497e-08 0 3.45e-08 0.0007 3.4503e-08 0 3.4597e-08 0 3.46e-08 0.0007 3.4603e-08 0 3.4697e-08 0 3.47e-08 0.0007 3.4703e-08 0 3.4797e-08 0 3.48e-08 0.0007 3.4803e-08 0 3.4897e-08 0 3.49e-08 0.0007 3.4903e-08 0 3.4997e-08 0 3.5e-08 0.0007 3.5003e-08 0 3.5097e-08 0 3.51e-08 0.0007 3.5103e-08 0 3.5197e-08 0 3.52e-08 0.0007 3.5203e-08 0 3.5297e-08 0 3.53e-08 0.0007 3.5303e-08 0 3.5397e-08 0 3.54e-08 0.0007 3.5403e-08 0 3.5497e-08 0 3.55e-08 0.0007 3.5503e-08 0 3.5597e-08 0 3.56e-08 0.0007 3.5603e-08 0 3.5697e-08 0 3.57e-08 0.0007 3.5703e-08 0 3.5797e-08 0 3.58e-08 0.0007 3.5803e-08 0 3.5897e-08 0 3.59e-08 0.0007 3.5903e-08 0 3.5997e-08 0 3.6e-08 0.0007 3.6003e-08 0 3.6097e-08 0 3.61e-08 0.0007 3.6103e-08 0 3.6197e-08 0 3.62e-08 0.0007 3.6203e-08 0 3.6297e-08 0 3.63e-08 0.0007 3.6303e-08 0 3.6397e-08 0 3.64e-08 0.0007 3.6403e-08 0 3.6497e-08 0 3.65e-08 0.0007 3.6503e-08 0 3.6597e-08 0 3.66e-08 0.0007 3.6603e-08 0 3.6697e-08 0 3.67e-08 0.0007 3.6703e-08 0 3.6797e-08 0 3.68e-08 0.0007 3.6803e-08 0 3.6897e-08 0 3.69e-08 0.0007 3.6903e-08 0 3.6997e-08 0 3.7e-08 0.0007 3.7003e-08 0 3.7097e-08 0 3.71e-08 0.0007 3.7103e-08 0 3.7197e-08 0 3.72e-08 0.0007 3.7203e-08 0 3.7297e-08 0 3.73e-08 0.0007 3.7303e-08 0 3.7397e-08 0 3.74e-08 0.0007 3.7403e-08 0 3.7497e-08 0 3.75e-08 0.0007 3.7503e-08 0 3.7597e-08 0 3.76e-08 0.0007 3.7603e-08 0 3.7697e-08 0 3.77e-08 0.0007 3.7703e-08 0 3.7797e-08 0 3.78e-08 0.0007 3.7803e-08 0 3.7897e-08 0 3.79e-08 0.0007 3.7903e-08 0 3.7997e-08 0 3.8e-08 0.0007 3.8003e-08 0 3.8097e-08 0 3.81e-08 0.0007 3.8103e-08 0 3.8197e-08 0 3.82e-08 0.0007 3.8203e-08 0 3.8297e-08 0 3.83e-08 0.0007 3.8303e-08 0 3.8397e-08 0 3.84e-08 0.0007 3.8403e-08 0 3.8497e-08 0 3.85e-08 0.0007 3.8503e-08 0 3.8597e-08 0 3.86e-08 0.0007 3.8603e-08 0 3.8697e-08 0 3.87e-08 0.0007 3.8703e-08 0 3.8797e-08 0 3.88e-08 0.0007 3.8803e-08 0 3.8897e-08 0 3.89e-08 0.0007 3.8903e-08 0 3.8997e-08 0 3.9e-08 0.0007 3.9003e-08 0 3.9097e-08 0 3.91e-08 0.0007 3.9103e-08 0 3.9197e-08 0 3.92e-08 0.0007 3.9203e-08 0 3.9297e-08 0 3.93e-08 0.0007 3.9303e-08 0 3.9397e-08 0 3.94e-08 0.0007 3.9403e-08 0 3.9497e-08 0 3.95e-08 0.0007 3.9503e-08 0 3.9597e-08 0 3.96e-08 0.0007 3.9603e-08 0 3.9697e-08 0 3.97e-08 0.0007 3.9703e-08 0 3.9797e-08 0 3.98e-08 0.0007 3.9803e-08 0 3.9897e-08 0 3.99e-08 0.0007 3.9903e-08 0)
I_SPL_A|B1 0 _SPL_A|3  PWL(0 0 5e-12 0.000154)
I_SPL_A|B2 0 _SPL_A|6  PWL(0 0 5e-12 0.0002464)
I_SPL_A|B3 0 _SPL_A|10  PWL(0 0 5e-12 0.000154)
I_SPL_A|B4 0 _SPL_A|13  PWL(0 0 5e-12 0.000154)
L_SPL_A|B1 _SPL_A|3 _SPL_A|1  9.175e-13
L_SPL_A|B2 _SPL_A|6 _SPL_A|4  7.666e-13
L_SPL_A|B3 _SPL_A|10 _SPL_A|8  1.928e-12
L_SPL_A|B4 _SPL_A|13 _SPL_A|11  8.786e-13
B_SPL_A|1 _SPL_A|1 _SPL_A|2 JJMIT AREA=2.5
B_SPL_A|2 _SPL_A|4 _SPL_A|5 JJMIT AREA=3.0
B_SPL_A|3 _SPL_A|8 _SPL_A|9 JJMIT AREA=2.5
B_SPL_A|4 _SPL_A|11 _SPL_A|12 JJMIT AREA=2.5
L_SPL_A|1 A_IN _SPL_A|1  2.063e-12
L_SPL_A|2 _SPL_A|1 _SPL_A|4  3.637e-12
L_SPL_A|3 _SPL_A|4 _SPL_A|7  1.278e-12
L_SPL_A|4 _SPL_A|7 _SPL_A|8  1.305e-12
L_SPL_A|5 _SPL_A|8 A_D  2.05e-12
L_SPL_A|6 _SPL_A|7 _SPL_A|11  1.315e-12
L_SPL_A|7 _SPL_A|11 A_OR  2.06e-12
L_SPL_A|P1 _SPL_A|2 0  4.676e-13
L_SPL_A|P2 _SPL_A|5 0  4.498e-13
L_SPL_A|P3 _SPL_A|9 0  5.183e-13
L_SPL_A|P4 _SPL_A|12 0  4.639e-13
R_SPL_A|B1 _SPL_A|1 _SPL_A|101  2.7439617672
L_SPL_A|RB1 _SPL_A|101 0  1.550338398468e-12
R_SPL_A|B2 _SPL_A|4 _SPL_A|104  2.286634806
L_SPL_A|RB2 _SPL_A|104 0  1.29194866539e-12
R_SPL_A|B3 _SPL_A|8 _SPL_A|108  2.7439617672
L_SPL_A|RB3 _SPL_A|108 0  1.550338398468e-12
R_SPL_A|B4 _SPL_A|11 _SPL_A|111  2.7439617672
L_SPL_A|RB4 _SPL_A|111 0  1.550338398468e-12
I_SPL_B|B1 0 _SPL_B|3  PWL(0 0 5e-12 0.000154)
I_SPL_B|B2 0 _SPL_B|6  PWL(0 0 5e-12 0.0002464)
I_SPL_B|B3 0 _SPL_B|10  PWL(0 0 5e-12 0.000154)
I_SPL_B|B4 0 _SPL_B|13  PWL(0 0 5e-12 0.000154)
L_SPL_B|B1 _SPL_B|3 _SPL_B|1  9.175e-13
L_SPL_B|B2 _SPL_B|6 _SPL_B|4  7.666e-13
L_SPL_B|B3 _SPL_B|10 _SPL_B|8  1.928e-12
L_SPL_B|B4 _SPL_B|13 _SPL_B|11  8.786e-13
B_SPL_B|1 _SPL_B|1 _SPL_B|2 JJMIT AREA=2.5
B_SPL_B|2 _SPL_B|4 _SPL_B|5 JJMIT AREA=3.0
B_SPL_B|3 _SPL_B|8 _SPL_B|9 JJMIT AREA=2.5
B_SPL_B|4 _SPL_B|11 _SPL_B|12 JJMIT AREA=2.5
L_SPL_B|1 B_IN _SPL_B|1  2.063e-12
L_SPL_B|2 _SPL_B|1 _SPL_B|4  3.637e-12
L_SPL_B|3 _SPL_B|4 _SPL_B|7  1.278e-12
L_SPL_B|4 _SPL_B|7 _SPL_B|8  1.305e-12
L_SPL_B|5 _SPL_B|8 B_D  2.05e-12
L_SPL_B|6 _SPL_B|7 _SPL_B|11  1.315e-12
L_SPL_B|7 _SPL_B|11 B_OR  2.06e-12
L_SPL_B|P1 _SPL_B|2 0  4.676e-13
L_SPL_B|P2 _SPL_B|5 0  4.498e-13
L_SPL_B|P3 _SPL_B|9 0  5.183e-13
L_SPL_B|P4 _SPL_B|12 0  4.639e-13
R_SPL_B|B1 _SPL_B|1 _SPL_B|101  2.7439617672
L_SPL_B|RB1 _SPL_B|101 0  1.550338398468e-12
R_SPL_B|B2 _SPL_B|4 _SPL_B|104  2.286634806
L_SPL_B|RB2 _SPL_B|104 0  1.29194866539e-12
R_SPL_B|B3 _SPL_B|8 _SPL_B|108  2.7439617672
L_SPL_B|RB3 _SPL_B|108 0  1.550338398468e-12
R_SPL_B|B4 _SPL_B|11 _SPL_B|111  2.7439617672
L_SPL_B|RB4 _SPL_B|111 0  1.550338398468e-12
B_OR|1 _OR|1 _OR|2 JJMIT AREA=2.5
B_OR|2 _OR|4 _OR|5 JJMIT AREA=2.5
B_OR|3 _OR|4 _OR|6 JJMIT AREA=1.92
B_OR|4 _OR|8 _OR|9 JJMIT AREA=2.5
B_OR|5 _OR|11 _OR|12 JJMIT AREA=2.5
B_OR|6 _OR|11 _OR|13 JJMIT AREA=1.92
B_OR|7 _OR|15 _OR|16 JJMIT AREA=2.53
B_OR|8 _OR|18 _OR|19 JJMIT AREA=2.5
I_OR|B1 0 _OR|3  PWL(0 0 5e-12 0.0001925)
I_OR|B2 0 _OR|10  PWL(0 0 5e-12 0.0001925)
I_OR|B3 0 _OR|14  PWL(0 0 5e-12 0.0002794)
I_OR|B4 0 _OR|17  PWL(0 0 5e-12 0.0002112)
I_OR|B5 0 _OR|20  PWL(0 0 5e-12 0.0001925)
L_OR|1 A_OR _OR|1  2.117e-12
L_OR|2 _OR|1 _OR|4  3.17e-12
L_OR|3 _OR|6 _OR|7  1.234e-12
L_OR|4 B_OR _OR|8  2.082e-12
L_OR|5 _OR|8 _OR|11  3.165e-12
L_OR|6 _OR|13 _OR|7  1.224e-12
L_OR|7 _OR|7 _OR|15  5.299e-12
L_OR|8 _OR|15 _OR|18  4.489e-12
L_OR|9 _OR|18 A_OR_B  2.077e-12
L_OR|P1 _OR|2 0  4.652e-13
L_OR|P2 _OR|5 0  4.457e-13
L_OR|P4 _OR|9 0  5.293e-13
L_OR|P5 _OR|12 0  4.452e-13
L_OR|P7 _OR|16 0  5.039e-13
L_OR|P8 _OR|19 0  4.984e-13
L_OR|B1 _OR|1 _OR|3  2e-12
L_OR|B2 _OR|8 _OR|10  2e-12
L_OR|B3 _OR|7 _OR|14  2e-12
L_OR|B4 _OR|15 _OR|17  2e-12
L_OR|B5 _OR|18 _OR|20  2e-12
R_OR|B1 _OR|1 _OR|101  2.7439617672
L_OR|RB1 _OR|101 0  1.550338398468e-12
R_OR|B2 _OR|4 _OR|104  2.7439617672
L_OR|RB2 _OR|104 0  1.550338398468e-12
R_OR|B3 _OR|4 _OR|106  3.572866884375
L_OR|RB3 _OR|106 _OR|6  2.018669789671875e-12
R_OR|B4 _OR|8 _OR|108  2.7439617672
L_OR|RB4 _OR|108 0  1.550338398468e-12
R_OR|B5 _OR|11 _OR|111  2.7439617672
L_OR|RB5 _OR|111 0  1.550338398468e-12
R_OR|B6 _OR|11 _OR|113  3.572866884375
L_OR|RB6 _OR|113 _OR|13  2.018669789671875e-12
R_OR|B7 _OR|15 _OR|115  2.7114246711462453
L_OR|RB7 _OR|115 0  1.5319549391976286e-12
R_OR|B8 _OR|18 _OR|118  2.7439617672
L_OR|RB8 _OR|118 0  1.550338398468e-12
B_NOT|1 _NOT|1 _NOT|2 JJMIT AREA=2.5
B_NOT|2 _NOT|4 _NOT|5 JJMIT AREA=2.57
B_NOT|3 _NOT|7 _NOT|8 JJMIT AREA=1.07
B_NOT|4 _NOT|13 _NOT|14 JJMIT AREA=2.5
B_NOT|5 _NOT|17 _NOT|18 JJMIT AREA=1.34
B_NOT|6 _NOT|10 _NOT|11 JJMIT AREA=3.03
B_NOT|7 _NOT|20 _NOT|18 JJMIT AREA=1.38
B_NOT|8 _NOT|18 _NOT|19 JJMIT AREA=0.8
B_NOT|9 _NOT|21 _NOT|22 JJMIT AREA=2.5
I_NOT|B1 0 _NOT|3  PWL(0 0 5e-12 0.0001925)
I_NOT|B2 0 _NOT|6  PWL(0 0 5e-12 9.57e-05)
I_NOT|B3 0 _NOT|9  PWL(0 0 5e-12 0.0002827)
I_NOT|B4 0 _NOT|15  PWL(0 0 5e-12 0.0001925)
I_NOT|B5 0 _NOT|23  PWL(0 0 5e-12 0.0001925)
L_NOT|B1 _NOT|3 _NOT|1  2e-12
L_NOT|B2 _NOT|6 _NOT|4  2e-12
L_NOT|B3 _NOT|8 _NOT|9  2e-12
L_NOT|B4 _NOT|13 _NOT|15  2e-12
L_NOT|B5 _NOT|21 _NOT|23  2e-12
L_NOT|1 A_OR_B _NOT|1  2.062e-12
L_NOT|2 _NOT|1 _NOT|4  1.889e-12
L_NOT|3 _NOT|4 _NOT|7  2.72e-12
L_NOT|4 CLK1 _NOT|13  2.057e-12
L_NOT|5 _NOT|13 _NOT|16  1.029e-12
L_NOT|6 _NOT|16 _NOT|17  1.241e-12
L_NOT|7 _NOT|16 _NOT|12  1.973e-12
L_NOT|8 _NOT|10 _NOT|12  1.003e-12
L_NOT|9 _NOT|10 _NOT|8  7.524e-12
L_NOT|10 _NOT|8 _NOT|20  1.234e-12
L_NOT|11 _NOT|18 _NOT|21  2.607e-12
L_NOT|12 _NOT|21 N0001  2.062e-12
L_NOT|P1 _NOT|2 0  5.271e-13
L_NOT|P2 _NOT|5 0  5.237e-13
L_NOT|P4 _NOT|14 0  4.759e-13
L_NOT|P6 _NOT|11 0  5.021e-13
L_NOT|P8 _NOT|19 0  6.33e-13
L_NOT|P9 _NOT|22 0  4.749e-13
R_NOT|B1 _NOT|1 _NOT|101  2.7439617672
L_NOT|RB1 _NOT|101 0  1.550338398468e-12
R_NOT|B2 _NOT|4 _NOT|104  2.6692235089494165
L_NOT|RB2 _NOT|104 _NOT|5  1.5081112825564204e-12
R_NOT|B3 _NOT|7 _NOT|107  6.411125624299065
L_NOT|RB3 _NOT|107 _NOT|8  3.622285977728972e-12
R_NOT|B4 _NOT|13 _NOT|113  2.7439617672
L_NOT|RB4 _NOT|113 0  1.550338398468e-12
R_NOT|B5 _NOT|17 _NOT|117  5.11933165522388
L_NOT|RB5 _NOT|117 _NOT|18  2.8924223852014925e-12
R_NOT|B6 _NOT|10 _NOT|110  2.2639948574257427
L_NOT|RB6 _NOT|110 0  1.2791570944455447e-12
R_NOT|B7 _NOT|20 _NOT|120  4.970945230434783
L_NOT|RB7 _NOT|120 _NOT|18  2.8085840551956523e-12
R_NOT|B8 _NOT|18 _NOT|118  8.574880522499999
L_NOT|RB8 _NOT|118 0  4.8448074952125e-12
R_NOT|B9 _NOT|21 _NOT|121  2.7439617672
L_NOT|RB9 _NOT|121 0  1.550338398468e-12
L_NOT|RD _NOT|12 _NOT|112  2e-12
R_NOT|D _NOT|112 0  4
B_DFF_A|1 _DFF_A|1 _DFF_A|2 JJMIT AREA=2.5
B_DFF_A|2 _DFF_A|4 _DFF_A|5 JJMIT AREA=1.61
B_DFF_A|3 _DFF_A|5 _DFF_A|6 JJMIT AREA=1.54
B_DFF_A|4 _DFF_A|8 _DFF_A|9 JJMIT AREA=1.69
B_DFF_A|5 _DFF_A|10 _DFF_A|8 JJMIT AREA=1.38
B_DFF_A|6 _DFF_A|11 _DFF_A|12 JJMIT AREA=2.5
B_DFF_A|7 _DFF_A|14 _DFF_A|15 JJMIT AREA=2.5
I_DFF_A|B1 0 _DFF_A|3  PWL(0 0 5e-12 0.0001925)
I_DFF_A|B2 0 _DFF_A|7  PWL(0 0 5e-12 0.0001903)
I_DFF_A|B3 0 _DFF_A|13  PWL(0 0 5e-12 0.0001925)
I_DFF_A|B4 0 _DFF_A|16  PWL(0 0 5e-12 0.0001925)
L_DFF_A|B1 _DFF_A|3 _DFF_A|1  2e-12
L_DFF_A|B2 _DFF_A|7 _DFF_A|5  2e-12
L_DFF_A|B3 _DFF_A|11 _DFF_A|13  2e-12
L_DFF_A|B4 _DFF_A|16 _DFF_A|14  2e-12
L_DFF_A|1 A_D _DFF_A|1  2.059e-12
L_DFF_A|2 _DFF_A|1 _DFF_A|4  4.123e-12
L_DFF_A|3 _DFF_A|5 _DFF_A|8  6.873e-12
L_DFF_A|4 _DFF_A|10 _DFF_A|11  5.195e-12
L_DFF_A|5 CLK2 _DFF_A|11  2.071e-12
L_DFF_A|6 _DFF_A|8 _DFF_A|14  3.287e-12
L_DFF_A|7 _DFF_A|14 A_AND  2.066e-12
L_DFF_A|P1 _DFF_A|2 0  5.042e-13
L_DFF_A|P3 _DFF_A|6 0  5.799e-13
L_DFF_A|P4 _DFF_A|9 0  5.733e-13
L_DFF_A|P6 _DFF_A|12 0  4.605e-13
L_DFF_A|P7 _DFF_A|15 0  4.961e-13
R_DFF_A|B1 _DFF_A|1 _DFF_A|101  2.7439617672
L_DFF_A|RB1 _DFF_A|101 0  1.550338398468e-12
R_DFF_A|B2 _DFF_A|4 _DFF_A|104  4.260810197515528
L_DFF_A|RB2 _DFF_A|104 _DFF_A|5  2.407357761596273e-12
R_DFF_A|B3 _DFF_A|5 _DFF_A|105  4.454483388311688
L_DFF_A|RB3 _DFF_A|105 0  2.516783114396104e-12
R_DFF_A|B4 _DFF_A|8 _DFF_A|108  4.059115040236686
L_DFF_A|RB4 _DFF_A|108 0  2.2933999977337278e-12
R_DFF_A|B5 _DFF_A|10 _DFF_A|110  4.970945230434783
L_DFF_A|RB5 _DFF_A|110 _DFF_A|8  2.8085840551956523e-12
R_DFF_A|B6 _DFF_A|11 _DFF_A|111  2.7439617672
L_DFF_A|RB6 _DFF_A|111 0  1.550338398468e-12
R_DFF_A|B7 _DFF_A|14 _DFF_A|114  2.7439617672
L_DFF_A|RB7 _DFF_A|114 0  1.550338398468e-12
B_DFF_B|1 _DFF_B|1 _DFF_B|2 JJMIT AREA=2.5
B_DFF_B|2 _DFF_B|4 _DFF_B|5 JJMIT AREA=1.61
B_DFF_B|3 _DFF_B|5 _DFF_B|6 JJMIT AREA=1.54
B_DFF_B|4 _DFF_B|8 _DFF_B|9 JJMIT AREA=1.69
B_DFF_B|5 _DFF_B|10 _DFF_B|8 JJMIT AREA=1.38
B_DFF_B|6 _DFF_B|11 _DFF_B|12 JJMIT AREA=2.5
B_DFF_B|7 _DFF_B|14 _DFF_B|15 JJMIT AREA=2.5
I_DFF_B|B1 0 _DFF_B|3  PWL(0 0 5e-12 0.0001925)
I_DFF_B|B2 0 _DFF_B|7  PWL(0 0 5e-12 0.0001903)
I_DFF_B|B3 0 _DFF_B|13  PWL(0 0 5e-12 0.0001925)
I_DFF_B|B4 0 _DFF_B|16  PWL(0 0 5e-12 0.0001925)
L_DFF_B|B1 _DFF_B|3 _DFF_B|1  2e-12
L_DFF_B|B2 _DFF_B|7 _DFF_B|5  2e-12
L_DFF_B|B3 _DFF_B|11 _DFF_B|13  2e-12
L_DFF_B|B4 _DFF_B|16 _DFF_B|14  2e-12
L_DFF_B|1 B_D _DFF_B|1  2.059e-12
L_DFF_B|2 _DFF_B|1 _DFF_B|4  4.123e-12
L_DFF_B|3 _DFF_B|5 _DFF_B|8  6.873e-12
L_DFF_B|4 _DFF_B|10 _DFF_B|11  5.195e-12
L_DFF_B|5 CLK3 _DFF_B|11  2.071e-12
L_DFF_B|6 _DFF_B|8 _DFF_B|14  3.287e-12
L_DFF_B|7 _DFF_B|14 B_AND  2.066e-12
L_DFF_B|P1 _DFF_B|2 0  5.042e-13
L_DFF_B|P3 _DFF_B|6 0  5.799e-13
L_DFF_B|P4 _DFF_B|9 0  5.733e-13
L_DFF_B|P6 _DFF_B|12 0  4.605e-13
L_DFF_B|P7 _DFF_B|15 0  4.961e-13
R_DFF_B|B1 _DFF_B|1 _DFF_B|101  2.7439617672
L_DFF_B|RB1 _DFF_B|101 0  1.550338398468e-12
R_DFF_B|B2 _DFF_B|4 _DFF_B|104  4.260810197515528
L_DFF_B|RB2 _DFF_B|104 _DFF_B|5  2.407357761596273e-12
R_DFF_B|B3 _DFF_B|5 _DFF_B|105  4.454483388311688
L_DFF_B|RB3 _DFF_B|105 0  2.516783114396104e-12
R_DFF_B|B4 _DFF_B|8 _DFF_B|108  4.059115040236686
L_DFF_B|RB4 _DFF_B|108 0  2.2933999977337278e-12
R_DFF_B|B5 _DFF_B|10 _DFF_B|110  4.970945230434783
L_DFF_B|RB5 _DFF_B|110 _DFF_B|8  2.8085840551956523e-12
R_DFF_B|B6 _DFF_B|11 _DFF_B|111  2.7439617672
L_DFF_B|RB6 _DFF_B|111 0  1.550338398468e-12
R_DFF_B|B7 _DFF_B|14 _DFF_B|114  2.7439617672
L_DFF_B|RB7 _DFF_B|114 0  1.550338398468e-12
B_AND|1 _AND|1 _AND|2 JJMIT AREA=2.5
B_AND|2 _AND|4 _AND|5 JJMIT AREA=2.5
B_AND|3 _AND|4 _AND|6 JJMIT AREA=1.92
B_AND|4 _AND|8 _AND|9 JJMIT AREA=2.5
B_AND|5 _AND|11 _AND|12 JJMIT AREA=2.5
B_AND|6 _AND|11 _AND|13 JJMIT AREA=1.92
B_AND|7 _AND|15 _AND|16 JJMIT AREA=2.53
B_AND|8 _AND|18 _AND|19 JJMIT AREA=2.5
I_AND|B1 0 _AND|3  PWL(0 0 5e-12 0.0001925)
I_AND|B2 0 _AND|10  PWL(0 0 5e-12 0.0001925)
I_AND|B3 0 _AND|14  PWL(0 0 5e-12 5.588e-05)
I_AND|B4 0 _AND|17  PWL(0 0 5e-12 0.0002112)
I_AND|B5 0 _AND|20  PWL(0 0 5e-12 0.0001925)
L_AND|1 A_AND _AND|1  2.117e-12
L_AND|2 _AND|1 _AND|4  3.17e-12
L_AND|3 _AND|6 _AND|7  1.234e-12
L_AND|4 B_AND _AND|8  2.082e-12
L_AND|5 _AND|8 _AND|11  3.165e-12
L_AND|6 _AND|13 _AND|7  1.224e-12
L_AND|7 _AND|7 _AND|15  5.299e-12
L_AND|8 _AND|15 _AND|18  4.489e-12
L_AND|9 _AND|18 N1000  2.077e-12
L_AND|P1 _AND|2 0  4.652e-13
L_AND|P2 _AND|5 0  4.457e-13
L_AND|P4 _AND|9 0  5.293e-13
L_AND|P5 _AND|12 0  4.452e-13
L_AND|P7 _AND|16 0  5.039e-13
L_AND|P8 _AND|19 0  4.984e-13
L_AND|B1 _AND|1 _AND|3  2e-12
L_AND|B2 _AND|8 _AND|10  2e-12
L_AND|B3 _AND|7 _AND|14  2e-12
L_AND|B4 _AND|15 _AND|17  2e-12
L_AND|B5 _AND|18 _AND|20  2e-12
R_AND|B1 _AND|1 _AND|101  2.7439617672
L_AND|RB1 _AND|101 0  1.550338398468e-12
R_AND|B2 _AND|4 _AND|104  2.7439617672
L_AND|RB2 _AND|104 0  1.550338398468e-12
R_AND|B3 _AND|4 _AND|106  3.572866884375
L_AND|RB3 _AND|106 _AND|6  2.018669789671875e-12
R_AND|B4 _AND|8 _AND|108  2.7439617672
L_AND|RB4 _AND|108 0  1.550338398468e-12
R_AND|B5 _AND|11 _AND|111  2.7439617672
L_AND|RB5 _AND|111 0  1.550338398468e-12
R_AND|B6 _AND|11 _AND|113  3.572866884375
L_AND|RB6 _AND|113 _AND|13  2.018669789671875e-12
R_AND|B7 _AND|15 _AND|115  2.7114246711462453
L_AND|RB7 _AND|115 0  1.5319549391976286e-12
R_AND|B8 _AND|18 _AND|118  2.7439617672
L_AND|RB8 _AND|118 0  1.550338398468e-12
B_XNOR|1 _XNOR|1 _XNOR|2 JJMIT AREA=2.5
B_XNOR|2 _XNOR|4 _XNOR|5 JJMIT AREA=2.5
B_XNOR|3 _XNOR|4 _XNOR|6 JJMIT AREA=1.92
B_XNOR|4 _XNOR|8 _XNOR|9 JJMIT AREA=2.5
B_XNOR|5 _XNOR|11 _XNOR|12 JJMIT AREA=2.5
B_XNOR|6 _XNOR|11 _XNOR|13 JJMIT AREA=1.92
B_XNOR|7 _XNOR|15 _XNOR|16 JJMIT AREA=2.53
B_XNOR|8 _XNOR|18 _XNOR|19 JJMIT AREA=2.5
I_XNOR|B1 0 _XNOR|3  PWL(0 0 5e-12 0.0001925)
I_XNOR|B2 0 _XNOR|10  PWL(0 0 5e-12 0.0001925)
I_XNOR|B3 0 _XNOR|14  PWL(0 0 5e-12 0.0002794)
I_XNOR|B4 0 _XNOR|17  PWL(0 0 5e-12 0.0002112)
I_XNOR|B5 0 _XNOR|20  PWL(0 0 5e-12 0.0001925)
L_XNOR|1 N0001 _XNOR|1  2.117e-12
L_XNOR|2 _XNOR|1 _XNOR|4  3.17e-12
L_XNOR|3 _XNOR|6 _XNOR|7  1.234e-12
L_XNOR|4 N1000 _XNOR|8  2.082e-12
L_XNOR|5 _XNOR|8 _XNOR|11  3.165e-12
L_XNOR|6 _XNOR|13 _XNOR|7  1.224e-12
L_XNOR|7 _XNOR|7 _XNOR|15  5.299e-12
L_XNOR|8 _XNOR|15 _XNOR|18  4.489e-12
L_XNOR|9 _XNOR|18 N1001  2.077e-12
L_XNOR|P1 _XNOR|2 0  4.652e-13
L_XNOR|P2 _XNOR|5 0  4.457e-13
L_XNOR|P4 _XNOR|9 0  5.293e-13
L_XNOR|P5 _XNOR|12 0  4.452e-13
L_XNOR|P7 _XNOR|16 0  5.039e-13
L_XNOR|P8 _XNOR|19 0  4.984e-13
L_XNOR|B1 _XNOR|1 _XNOR|3  2e-12
L_XNOR|B2 _XNOR|8 _XNOR|10  2e-12
L_XNOR|B3 _XNOR|7 _XNOR|14  2e-12
L_XNOR|B4 _XNOR|15 _XNOR|17  2e-12
L_XNOR|B5 _XNOR|18 _XNOR|20  2e-12
R_XNOR|B1 _XNOR|1 _XNOR|101  2.7439617672
L_XNOR|RB1 _XNOR|101 0  1.550338398468e-12
R_XNOR|B2 _XNOR|4 _XNOR|104  2.7439617672
L_XNOR|RB2 _XNOR|104 0  1.550338398468e-12
R_XNOR|B3 _XNOR|4 _XNOR|106  3.572866884375
L_XNOR|RB3 _XNOR|106 _XNOR|6  2.018669789671875e-12
R_XNOR|B4 _XNOR|8 _XNOR|108  2.7439617672
L_XNOR|RB4 _XNOR|108 0  1.550338398468e-12
R_XNOR|B5 _XNOR|11 _XNOR|111  2.7439617672
L_XNOR|RB5 _XNOR|111 0  1.550338398468e-12
R_XNOR|B6 _XNOR|11 _XNOR|113  3.572866884375
L_XNOR|RB6 _XNOR|113 _XNOR|13  2.018669789671875e-12
R_XNOR|B7 _XNOR|15 _XNOR|115  2.7114246711462453
L_XNOR|RB7 _XNOR|115 0  1.5319549391976286e-12
R_XNOR|B8 _XNOR|18 _XNOR|118  2.7439617672
L_XNOR|RB8 _XNOR|118 0  1.550338398468e-12
.print DEVI ROUT
.print DEVI IA|A
.print DEVI IB|B
.print DEVI IT1|T
.print DEVI IT2|T
.print DEVI IT3|T
.print DEVI I_SPL_A|B1
.print DEVI I_SPL_A|B2
.print DEVI I_SPL_A|B3
.print DEVI I_SPL_A|B4
.print DEVI L_SPL_A|B1
.print DEVI L_SPL_A|B2
.print DEVI L_SPL_A|B3
.print DEVI L_SPL_A|B4
.print DEVI B_SPL_A|1
.print DEVI B_SPL_A|2
.print DEVI B_SPL_A|3
.print DEVI B_SPL_A|4
.print DEVI L_SPL_A|1
.print DEVI L_SPL_A|2
.print DEVI L_SPL_A|3
.print DEVI L_SPL_A|4
.print DEVI L_SPL_A|5
.print DEVI L_SPL_A|6
.print DEVI L_SPL_A|7
.print DEVI L_SPL_A|P1
.print DEVI L_SPL_A|P2
.print DEVI L_SPL_A|P3
.print DEVI L_SPL_A|P4
.print DEVI R_SPL_A|B1
.print DEVI L_SPL_A|RB1
.print DEVI R_SPL_A|B2
.print DEVI L_SPL_A|RB2
.print DEVI R_SPL_A|B3
.print DEVI L_SPL_A|RB3
.print DEVI R_SPL_A|B4
.print DEVI L_SPL_A|RB4
.print DEVI I_SPL_B|B1
.print DEVI I_SPL_B|B2
.print DEVI I_SPL_B|B3
.print DEVI I_SPL_B|B4
.print DEVI L_SPL_B|B1
.print DEVI L_SPL_B|B2
.print DEVI L_SPL_B|B3
.print DEVI L_SPL_B|B4
.print DEVI B_SPL_B|1
.print DEVI B_SPL_B|2
.print DEVI B_SPL_B|3
.print DEVI B_SPL_B|4
.print DEVI L_SPL_B|1
.print DEVI L_SPL_B|2
.print DEVI L_SPL_B|3
.print DEVI L_SPL_B|4
.print DEVI L_SPL_B|5
.print DEVI L_SPL_B|6
.print DEVI L_SPL_B|7
.print DEVI L_SPL_B|P1
.print DEVI L_SPL_B|P2
.print DEVI L_SPL_B|P3
.print DEVI L_SPL_B|P4
.print DEVI R_SPL_B|B1
.print DEVI L_SPL_B|RB1
.print DEVI R_SPL_B|B2
.print DEVI L_SPL_B|RB2
.print DEVI R_SPL_B|B3
.print DEVI L_SPL_B|RB3
.print DEVI R_SPL_B|B4
.print DEVI L_SPL_B|RB4
.print DEVI B_OR|1
.print DEVI B_OR|2
.print DEVI B_OR|3
.print DEVI B_OR|4
.print DEVI B_OR|5
.print DEVI B_OR|6
.print DEVI B_OR|7
.print DEVI B_OR|8
.print DEVI I_OR|B1
.print DEVI I_OR|B2
.print DEVI I_OR|B3
.print DEVI I_OR|B4
.print DEVI I_OR|B5
.print DEVI L_OR|1
.print DEVI L_OR|2
.print DEVI L_OR|3
.print DEVI L_OR|4
.print DEVI L_OR|5
.print DEVI L_OR|6
.print DEVI L_OR|7
.print DEVI L_OR|8
.print DEVI L_OR|9
.print DEVI L_OR|P1
.print DEVI L_OR|P2
.print DEVI L_OR|P4
.print DEVI L_OR|P5
.print DEVI L_OR|P7
.print DEVI L_OR|P8
.print DEVI L_OR|B1
.print DEVI L_OR|B2
.print DEVI L_OR|B3
.print DEVI L_OR|B4
.print DEVI L_OR|B5
.print DEVI R_OR|B1
.print DEVI L_OR|RB1
.print DEVI R_OR|B2
.print DEVI L_OR|RB2
.print DEVI R_OR|B3
.print DEVI L_OR|RB3
.print DEVI R_OR|B4
.print DEVI L_OR|RB4
.print DEVI R_OR|B5
.print DEVI L_OR|RB5
.print DEVI R_OR|B6
.print DEVI L_OR|RB6
.print DEVI R_OR|B7
.print DEVI L_OR|RB7
.print DEVI R_OR|B8
.print DEVI L_OR|RB8
.print DEVI B_NOT|1
.print DEVI B_NOT|2
.print DEVI B_NOT|3
.print DEVI B_NOT|4
.print DEVI B_NOT|5
.print DEVI B_NOT|6
.print DEVI B_NOT|7
.print DEVI B_NOT|8
.print DEVI B_NOT|9
.print DEVI I_NOT|B1
.print DEVI I_NOT|B2
.print DEVI I_NOT|B3
.print DEVI I_NOT|B4
.print DEVI I_NOT|B5
.print DEVI L_NOT|B1
.print DEVI L_NOT|B2
.print DEVI L_NOT|B3
.print DEVI L_NOT|B4
.print DEVI L_NOT|B5
.print DEVI L_NOT|1
.print DEVI L_NOT|2
.print DEVI L_NOT|3
.print DEVI L_NOT|4
.print DEVI L_NOT|5
.print DEVI L_NOT|6
.print DEVI L_NOT|7
.print DEVI L_NOT|8
.print DEVI L_NOT|9
.print DEVI L_NOT|10
.print DEVI L_NOT|11
.print DEVI L_NOT|12
.print DEVI L_NOT|P1
.print DEVI L_NOT|P2
.print DEVI L_NOT|P4
.print DEVI L_NOT|P6
.print DEVI L_NOT|P8
.print DEVI L_NOT|P9
.print DEVI R_NOT|B1
.print DEVI L_NOT|RB1
.print DEVI R_NOT|B2
.print DEVI L_NOT|RB2
.print DEVI R_NOT|B3
.print DEVI L_NOT|RB3
.print DEVI R_NOT|B4
.print DEVI L_NOT|RB4
.print DEVI R_NOT|B5
.print DEVI L_NOT|RB5
.print DEVI R_NOT|B6
.print DEVI L_NOT|RB6
.print DEVI R_NOT|B7
.print DEVI L_NOT|RB7
.print DEVI R_NOT|B8
.print DEVI L_NOT|RB8
.print DEVI R_NOT|B9
.print DEVI L_NOT|RB9
.print DEVI L_NOT|RD
.print DEVI R_NOT|D
.print DEVI B_DFF_A|1
.print DEVI B_DFF_A|2
.print DEVI B_DFF_A|3
.print DEVI B_DFF_A|4
.print DEVI B_DFF_A|5
.print DEVI B_DFF_A|6
.print DEVI B_DFF_A|7
.print DEVI I_DFF_A|B1
.print DEVI I_DFF_A|B2
.print DEVI I_DFF_A|B3
.print DEVI I_DFF_A|B4
.print DEVI L_DFF_A|B1
.print DEVI L_DFF_A|B2
.print DEVI L_DFF_A|B3
.print DEVI L_DFF_A|B4
.print DEVI L_DFF_A|1
.print DEVI L_DFF_A|2
.print DEVI L_DFF_A|3
.print DEVI L_DFF_A|4
.print DEVI L_DFF_A|5
.print DEVI L_DFF_A|6
.print DEVI L_DFF_A|7
.print DEVI L_DFF_A|P1
.print DEVI L_DFF_A|P3
.print DEVI L_DFF_A|P4
.print DEVI L_DFF_A|P6
.print DEVI L_DFF_A|P7
.print DEVI R_DFF_A|B1
.print DEVI L_DFF_A|RB1
.print DEVI R_DFF_A|B2
.print DEVI L_DFF_A|RB2
.print DEVI R_DFF_A|B3
.print DEVI L_DFF_A|RB3
.print DEVI R_DFF_A|B4
.print DEVI L_DFF_A|RB4
.print DEVI R_DFF_A|B5
.print DEVI L_DFF_A|RB5
.print DEVI R_DFF_A|B6
.print DEVI L_DFF_A|RB6
.print DEVI R_DFF_A|B7
.print DEVI L_DFF_A|RB7
.print DEVI B_DFF_B|1
.print DEVI B_DFF_B|2
.print DEVI B_DFF_B|3
.print DEVI B_DFF_B|4
.print DEVI B_DFF_B|5
.print DEVI B_DFF_B|6
.print DEVI B_DFF_B|7
.print DEVI I_DFF_B|B1
.print DEVI I_DFF_B|B2
.print DEVI I_DFF_B|B3
.print DEVI I_DFF_B|B4
.print DEVI L_DFF_B|B1
.print DEVI L_DFF_B|B2
.print DEVI L_DFF_B|B3
.print DEVI L_DFF_B|B4
.print DEVI L_DFF_B|1
.print DEVI L_DFF_B|2
.print DEVI L_DFF_B|3
.print DEVI L_DFF_B|4
.print DEVI L_DFF_B|5
.print DEVI L_DFF_B|6
.print DEVI L_DFF_B|7
.print DEVI L_DFF_B|P1
.print DEVI L_DFF_B|P3
.print DEVI L_DFF_B|P4
.print DEVI L_DFF_B|P6
.print DEVI L_DFF_B|P7
.print DEVI R_DFF_B|B1
.print DEVI L_DFF_B|RB1
.print DEVI R_DFF_B|B2
.print DEVI L_DFF_B|RB2
.print DEVI R_DFF_B|B3
.print DEVI L_DFF_B|RB3
.print DEVI R_DFF_B|B4
.print DEVI L_DFF_B|RB4
.print DEVI R_DFF_B|B5
.print DEVI L_DFF_B|RB5
.print DEVI R_DFF_B|B6
.print DEVI L_DFF_B|RB6
.print DEVI R_DFF_B|B7
.print DEVI L_DFF_B|RB7
.print DEVI B_AND|1
.print DEVI B_AND|2
.print DEVI B_AND|3
.print DEVI B_AND|4
.print DEVI B_AND|5
.print DEVI B_AND|6
.print DEVI B_AND|7
.print DEVI B_AND|8
.print DEVI I_AND|B1
.print DEVI I_AND|B2
.print DEVI I_AND|B3
.print DEVI I_AND|B4
.print DEVI I_AND|B5
.print DEVI L_AND|1
.print DEVI L_AND|2
.print DEVI L_AND|3
.print DEVI L_AND|4
.print DEVI L_AND|5
.print DEVI L_AND|6
.print DEVI L_AND|7
.print DEVI L_AND|8
.print DEVI L_AND|9
.print DEVI L_AND|P1
.print DEVI L_AND|P2
.print DEVI L_AND|P4
.print DEVI L_AND|P5
.print DEVI L_AND|P7
.print DEVI L_AND|P8
.print DEVI L_AND|B1
.print DEVI L_AND|B2
.print DEVI L_AND|B3
.print DEVI L_AND|B4
.print DEVI L_AND|B5
.print DEVI R_AND|B1
.print DEVI L_AND|RB1
.print DEVI R_AND|B2
.print DEVI L_AND|RB2
.print DEVI R_AND|B3
.print DEVI L_AND|RB3
.print DEVI R_AND|B4
.print DEVI L_AND|RB4
.print DEVI R_AND|B5
.print DEVI L_AND|RB5
.print DEVI R_AND|B6
.print DEVI L_AND|RB6
.print DEVI R_AND|B7
.print DEVI L_AND|RB7
.print DEVI R_AND|B8
.print DEVI L_AND|RB8
.print DEVI B_XNOR|1
.print DEVI B_XNOR|2
.print DEVI B_XNOR|3
.print DEVI B_XNOR|4
.print DEVI B_XNOR|5
.print DEVI B_XNOR|6
.print DEVI B_XNOR|7
.print DEVI B_XNOR|8
.print DEVI I_XNOR|B1
.print DEVI I_XNOR|B2
.print DEVI I_XNOR|B3
.print DEVI I_XNOR|B4
.print DEVI I_XNOR|B5
.print DEVI L_XNOR|1
.print DEVI L_XNOR|2
.print DEVI L_XNOR|3
.print DEVI L_XNOR|4
.print DEVI L_XNOR|5
.print DEVI L_XNOR|6
.print DEVI L_XNOR|7
.print DEVI L_XNOR|8
.print DEVI L_XNOR|9
.print DEVI L_XNOR|P1
.print DEVI L_XNOR|P2
.print DEVI L_XNOR|P4
.print DEVI L_XNOR|P5
.print DEVI L_XNOR|P7
.print DEVI L_XNOR|P8
.print DEVI L_XNOR|B1
.print DEVI L_XNOR|B2
.print DEVI L_XNOR|B3
.print DEVI L_XNOR|B4
.print DEVI L_XNOR|B5
.print DEVI R_XNOR|B1
.print DEVI L_XNOR|RB1
.print DEVI R_XNOR|B2
.print DEVI L_XNOR|RB2
.print DEVI R_XNOR|B3
.print DEVI L_XNOR|RB3
.print DEVI R_XNOR|B4
.print DEVI L_XNOR|RB4
.print DEVI R_XNOR|B5
.print DEVI L_XNOR|RB5
.print DEVI R_XNOR|B6
.print DEVI L_XNOR|RB6
.print DEVI R_XNOR|B7
.print DEVI L_XNOR|RB7
.print DEVI R_XNOR|B8
.print DEVI L_XNOR|RB8
.print V _OR|1
.print V CLK1
.print V _SPL_A|8
.print V _SPL_B|8
.print V _NOT|113
.print V _OR|12
.print V _XNOR|11
.print V _DFF_B|13
.print V _AND|4
.print V _OR|5
.print V _DFF_A|8
.print V _XNOR|115
.print V _OR|115
.print V _SPL_A|3
.print V _DFF_B|4
.print V _XNOR|6
.print V _OR|11
.print V _OR|4
.print V _SPL_B|9
.print V _OR|10
.print V _XNOR|113
.print V _SPL_A|10
.print V _SPL_B|12
.print V _AND|2
.print V _OR|8
.print V _SPL_A|13
.print V _SPL_B|10
.print V _NOT|110
.print V _NOT|10
.print V _OR|16
.print V _XNOR|3
.print V _OR|19
.print V _DFF_A|101
.print V _DFF_A|4
.print V _NOT|14
.print V _DFF_B|101
.print V _AND|108
.print V _AND|1
.print V _XNOR|7
.print V _DFF_A|13
.print V _DFF_B|110
.print V _DFF_B|7
.print V _SPL_B|3
.print V _DFF_A|11
.print V _XNOR|19
.print V _SPL_B|7
.print V _DFF_A|14
.print V _SPL_A|5
.print V _NOT|5
.print V _AND|18
.print V _NOT|23
.print V _DFF_B|3
.print V _SPL_B|6
.print V _DFF_A|7
.print V _DFF_A|12
.print V _OR|118
.print V _NOT|118
.print V _XNOR|104
.print V _NOT|9
.print V _OR|6
.print V _NOT|120
.print V _XNOR|101
.print V _SPL_A|108
.print V _NOT|21
.print V _DFF_B|114
.print V B_IN
.print V _OR|111
.print V _OR|13
.print V _NOT|104
.print V _AND|20
.print V _AND|111
.print V _XNOR|10
.print V _NOT|13
.print V _DFF_A|1
.print V _SPL_B|4
.print V _DFF_A|6
.print V _SPL_B|11
.print V _AND|115
.print V N1001
.print V _NOT|121
.print V _DFF_B|14
.print V _AND|8
.print V _AND|16
.print V _DFF_A|3
.print V _NOT|18
.print V _NOT|20
.print V _DFF_B|2
.print V _DFF_B|11
.print V B_D
.print V _NOT|4
.print V _DFF_A|114
.print V _NOT|15
.print V CLK2
.print V _SPL_A|9
.print V A_OR
.print V _OR|7
.print V _AND|3
.print V _NOT|3
.print V _DFF_A|5
.print V _NOT|7
.print V _XNOR|18
.print V _OR|2
.print V _OR|9
.print V A_D
.print V _NOT|117
.print V _XNOR|111
.print V _SPL_A|12
.print V _AND|12
.print V _DFF_B|111
.print V CLK3
.print V _OR|18
.print V _AND|6
.print V _DFF_B|9
.print V _AND|14
.print V _SPL_A|104
.print V _XNOR|5
.print V N1000
.print V _XNOR|20
.print V _OR|17
.print V _NOT|22
.print V _OR|113
.print V _XNOR|1
.print V _NOT|17
.print V _NOT|8
.print V _NOT|1
.print V _XNOR|13
.print V _XNOR|15
.print V _AND|11
.print V _DFF_A|10
.print V _DFF_B|15
.print V _DFF_B|104
.print V _XNOR|14
.print V _AND|7
.print V _DFF_A|104
.print V _SPL_A|1
.print V _DFF_A|9
.print V _XNOR|12
.print V _OR|106
.print V _SPL_B|104
.print V _AND|19
.print V _AND|13
.print V _NOT|6
.print V _AND|101
.print V B_OR
.print V _AND|104
.print V _SPL_A|6
.print V _NOT|11
.print V _AND|113
.print V _XNOR|106
.print V _XNOR|9
.print V _XNOR|4
.print V _XNOR|16
.print V _XNOR|108
.print V _SPL_B|108
.print V _DFF_A|105
.print V _AND|118
.print V _XNOR|118
.print V _OR|104
.print V _SPL_B|5
.print V _AND|5
.print V _NOT|107
.print V A_AND
.print V _SPL_B|1
.print V _DFF_B|10
.print V B_AND
.print V _NOT|16
.print V _AND|9
.print V _OR|3
.print V _XNOR|2
.print V A_IN
.print V _NOT|2
.print V _XNOR|8
.print V _DFF_A|15
.print V _SPL_A|101
.print V _NOT|112
.print V _DFF_A|2
.print V _SPL_A|111
.print V _DFF_A|16
.print V N0001
.print V _SPL_A|7
.print V _DFF_B|5
.print V _OR|108
.print V _SPL_A|4
.print V _DFF_A|111
.print V _DFF_B|105
.print V _AND|17
.print V _DFF_A|110
.print V _AND|10
.print V _OR|15
.print V _OR|20
.print V _OR|14
.print V _DFF_B|6
.print V _SPL_A|11
.print V _DFF_B|16
.print V _DFF_B|108
.print V _AND|15
.print V _AND|106
.print V _NOT|12
.print V _SPL_B|2
.print V _SPL_B|101
.print V _DFF_A|108
.print V _SPL_A|2
.print V _OR|101
.print V _NOT|101
.print V _SPL_B|111
.print V _XNOR|17
.print V _DFF_B|1
.print V _DFF_B|12
.print V A_OR_B
.print V _DFF_B|8
.print V _SPL_B|13
.print V _NOT|19
.print DEVP B_SPL_A|1
.print DEVP B_SPL_A|2
.print DEVP B_SPL_A|3
.print DEVP B_SPL_A|4
.print DEVP B_SPL_B|1
.print DEVP B_SPL_B|2
.print DEVP B_SPL_B|3
.print DEVP B_SPL_B|4
.print DEVP B_OR|1
.print DEVP B_OR|2
.print DEVP B_OR|3
.print DEVP B_OR|4
.print DEVP B_OR|5
.print DEVP B_OR|6
.print DEVP B_OR|7
.print DEVP B_OR|8
.print DEVP B_NOT|1
.print DEVP B_NOT|2
.print DEVP B_NOT|3
.print DEVP B_NOT|4
.print DEVP B_NOT|5
.print DEVP B_NOT|6
.print DEVP B_NOT|7
.print DEVP B_NOT|8
.print DEVP B_NOT|9
.print DEVP B_DFF_A|1
.print DEVP B_DFF_A|2
.print DEVP B_DFF_A|3
.print DEVP B_DFF_A|4
.print DEVP B_DFF_A|5
.print DEVP B_DFF_A|6
.print DEVP B_DFF_A|7
.print DEVP B_DFF_B|1
.print DEVP B_DFF_B|2
.print DEVP B_DFF_B|3
.print DEVP B_DFF_B|4
.print DEVP B_DFF_B|5
.print DEVP B_DFF_B|6
.print DEVP B_DFF_B|7
.print DEVP B_AND|1
.print DEVP B_AND|2
.print DEVP B_AND|3
.print DEVP B_AND|4
.print DEVP B_AND|5
.print DEVP B_AND|6
.print DEVP B_AND|7
.print DEVP B_AND|8
.print DEVP B_XNOR|1
.print DEVP B_XNOR|2
.print DEVP B_XNOR|3
.print DEVP B_XNOR|4
.print DEVP B_XNOR|5
.print DEVP B_XNOR|6
.print DEVP B_XNOR|7
.print DEVP B_XNOR|8
