*
.PARAM PHI0=2.067833848e-15
.PARAM B0=1
.PARAM IC0=0.0001
.PARAM ICRS=0.0006859904418
.PARAM B0RS=6.859904418
.PARAM RSHEET=2
.PARAM LSHEET=1.13e-12
.PARAM LP=2e-13
.PARAM LPTL=2e-12
.PARAM IC=2.5
.PARAM LB=2e-12
.PARAM BIASCOEF=0.7
.PARAM OFFSET1=0.0
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.TRAN 0.5E-12 6E-09
ROUT ABXCD 0  1
IT1|T 0 T1  PWL(0 0 2.97e-10 0 3e-10 0.002 3.03e-10 0 5.97e-10 0 6e-10 0.002 6.03e-10 0 8.97e-10 0 9e-10 0.002 9.03e-10 0 1.197e-09 0 1.2e-09 0.002 1.203e-09 0 1.497e-09 0 1.5e-09 0.002 1.503e-09 0 1.797e-09 0 1.8e-09 0.002 1.803e-09 0 2.097e-09 0 2.1e-09 0.002 2.103e-09 0 2.397e-09 0 2.4e-09 0.002 2.403e-09 0 2.697e-09 0 2.7e-09 0.002 2.703e-09 0 2.997e-09 0 3e-09 0.002 3.003e-09 0 3.297e-09 0 3.3e-09 0.002 3.303e-09 0 3.597e-09 0 3.6e-09 0.002 3.603e-09 0 3.897e-09 0 3.9e-09 0.002 3.903e-09 0 4.197e-09 0 4.2e-09 0.002 4.203e-09 0 4.497e-09 0 4.5e-09 0.002 4.503e-09 0 4.797e-09 0 4.8e-09 0.002 4.803e-09 0 5.097e-09 0 5.1e-09 0.002 5.103e-09 0 5.397e-09 0 5.4e-09 0.002 5.403e-09 0 5.697e-09 0 5.7e-09 0.002 5.703e-09 0 5.997e-09 0 6e-09 0.002 6.003e-09 0 6.297e-09 0 6.3e-09 0.002 6.303e-09 0 6.597e-09 0 6.6e-09 0.002 6.603e-09 0 6.897e-09 0 6.9e-09 0.002 6.903e-09 0 7.197e-09 0 7.2e-09 0.002 7.203e-09 0 7.497e-09 0 7.5e-09 0.002 7.503e-09 0 7.797e-09 0 7.8e-09 0.002 7.803e-09 0 8.097e-09 0 8.1e-09 0.002 8.103e-09 0 8.397e-09 0 8.4e-09 0.002 8.403e-09 0 8.697e-09 0 8.7e-09 0.002 8.703e-09 0 8.997e-09 0 9e-09 0.002 9.003e-09 0 9.297e-09 0 9.3e-09 0.002 9.303e-09 0 9.597e-09 0 9.6e-09 0.002 9.603e-09 0 9.897e-09 0 9.9e-09 0.002 9.903e-09 0 1.0197e-08 0 1.02e-08 0.002 1.0203e-08 0 1.0497e-08 0 1.05e-08 0.002 1.0503e-08 0 1.0797e-08 0 1.08e-08 0.002 1.0803e-08 0 1.1097e-08 0 1.11e-08 0.002 1.1103e-08 0 1.1397e-08 0 1.14e-08 0.002 1.1403e-08 0 1.1697e-08 0 1.17e-08 0.002 1.1703e-08 0)
IDATA_A|A 0 A  PWL(0 0 6.57e-10 0 6.6e-10 0.0005 6.63e-10 0 1.257e-09 0 1.26e-09 0.0005 1.263e-09 0 1.857e-09 0 1.86e-09 0.0005 1.863e-09 0 2.457e-09 0 2.46e-09 0.0005 2.463e-09 0 3.057e-09 0 3.06e-09 0.0005 3.063e-09 0 3.657e-09 0 3.66e-09 0.0005 3.663e-09 0 4.257e-09 0 4.26e-09 0.0005 4.263e-09 0 4.857e-09 0 4.86e-09 0.0005 4.863e-09 0 5.457e-09 0 5.46e-09 0.0005 5.463e-09 0 6.057e-09 0 6.06e-09 0.0005 6.063e-09 0 6.657e-09 0 6.66e-09 0.0005 6.663e-09 0 7.257e-09 0 7.26e-09 0.0005 7.263e-09 0 7.857e-09 0 7.86e-09 0.0005 7.863e-09 0 8.457e-09 0 8.46e-09 0.0005 8.463e-09 0 9.057e-09 0 9.06e-09 0.0005 9.063e-09 0 9.657e-09 0 9.66e-09 0.0005 9.663e-09 0 1.0257e-08 0 1.026e-08 0.0005 1.0263e-08 0 1.0857e-08 0 1.086e-08 0.0005 1.0863e-08 0 1.1457e-08 0 1.146e-08 0.0005 1.1463e-08 0)
IDATA_B|B 0 B  PWL(0 0 1.017e-09 0 1.02e-09 0.0005 1.023e-09 0 1.317e-09 0 1.32e-09 0.0005 1.323e-09 0 2.217e-09 0 2.22e-09 0.0005 2.223e-09 0 2.517e-09 0 2.52e-09 0.0005 2.523e-09 0 3.417e-09 0 3.42e-09 0.0005 3.423e-09 0 3.717e-09 0 3.72e-09 0.0005 3.723e-09 0 4.617e-09 0 4.62e-09 0.0005 4.623e-09 0 4.917e-09 0 4.92e-09 0.0005 4.923e-09 0 5.817e-09 0 5.82e-09 0.0005 5.823e-09 0 6.117e-09 0 6.12e-09 0.0005 6.123e-09 0 7.017e-09 0 7.02e-09 0.0005 7.023e-09 0 7.317e-09 0 7.32e-09 0.0005 7.323e-09 0 8.217e-09 0 8.22e-09 0.0005 8.223e-09 0 8.517e-09 0 8.52e-09 0.0005 8.523e-09 0 9.417e-09 0 9.42e-09 0.0005 9.423e-09 0 9.717e-09 0 9.72e-09 0.0005 9.723e-09 0 1.0617e-08 0 1.062e-08 0.0005 1.0623e-08 0 1.0917e-08 0 1.092e-08 0.0005 1.0923e-08 0 1.1817e-08 0 1.182e-08 0.0005 1.1823e-08 0)
IDATA_C|T 0 C  PWL(0 0 1.677e-09 0 1.68e-09 0.0005 1.683e-09 0 1.977e-09 0 1.98e-09 0.0005 1.983e-09 0 2.277e-09 0 2.28e-09 0.0005 2.283e-09 0 2.577e-09 0 2.58e-09 0.0005 2.583e-09 0 4.077e-09 0 4.08e-09 0.0005 4.083e-09 0 4.377e-09 0 4.38e-09 0.0005 4.383e-09 0 4.677e-09 0 4.68e-09 0.0005 4.683e-09 0 4.977e-09 0 4.98e-09 0.0005 4.983e-09 0 6.477e-09 0 6.48e-09 0.0005 6.483e-09 0 6.777e-09 0 6.78e-09 0.0005 6.783e-09 0 7.077e-09 0 7.08e-09 0.0005 7.083e-09 0 7.377e-09 0 7.38e-09 0.0005 7.383e-09 0 8.877e-09 0 8.88e-09 0.0005 8.883e-09 0 9.177e-09 0 9.18e-09 0.0005 9.183e-09 0 9.477e-09 0 9.48e-09 0.0005 9.483e-09 0 9.777e-09 0 9.78e-09 0.0005 9.783e-09 0 1.1277e-08 0 1.128e-08 0.0005 1.1283e-08 0 1.1577e-08 0 1.158e-08 0.0005 1.1583e-08 0 1.1877e-08 0 1.188e-08 0.0005 1.1883e-08 0)
IDATA_D|T 0 D  PWL(0 0 2.937e-09 0 2.94e-09 0.0005 2.943e-09 0 3.237e-09 0 3.24e-09 0.0005 3.243e-09 0 3.537e-09 0 3.54e-09 0.0005 3.543e-09 0 3.837e-09 0 3.84e-09 0.0005 3.843e-09 0 4.137e-09 0 4.14e-09 0.0005 4.143e-09 0 4.437e-09 0 4.44e-09 0.0005 4.443e-09 0 4.737e-09 0 4.74e-09 0.0005 4.743e-09 0 5.037e-09 0 5.04e-09 0.0005 5.043e-09 0 7.737e-09 0 7.74e-09 0.0005 7.743e-09 0 8.037e-09 0 8.04e-09 0.0005 8.043e-09 0 8.337e-09 0 8.34e-09 0.0005 8.343e-09 0 8.637e-09 0 8.64e-09 0.0005 8.643e-09 0 8.937e-09 0 8.94e-09 0.0005 8.943e-09 0 9.237e-09 0 9.24e-09 0.0005 9.243e-09 0 9.537e-09 0 9.54e-09 0.0005 9.543e-09 0 9.837e-09 0 9.84e-09 0.0005 9.843e-09 0)
B_AND_1|1 _AND_1|1 _AND_1|2 JJMIT AREA=2.5
B_AND_1|2 _AND_1|4 _AND_1|5 JJMIT AREA=1.7857142857142858
B_AND_1|3 _AND_1|5 _AND_1|6 JJMIT AREA=2.5
B_AND_1|4 _AND_1|8 _AND_1|9 JJMIT AREA=1.7857142857142858
B_AND_1|5 _AND_1|8 _AND_1|11 JJMIT AREA=2.5
B_AND_1|6 _AND_1|12 _AND_1|13 JJMIT AREA=1.7857142857142858
B_AND_1|7 _AND_1|14 _AND_1|15 JJMIT AREA=2.5
B_AND_1|8 _AND_1|17 _AND_1|18 JJMIT AREA=1.7857142857142858
B_AND_1|9 _AND_1|18 _AND_1|19 JJMIT AREA=2.5
B_AND_1|10 _AND_1|21 _AND_1|22 JJMIT AREA=1.7857142857142858
B_AND_1|11 _AND_1|21 _AND_1|23 JJMIT AREA=2.5
B_AND_1|12 _AND_1|24 _AND_1|13 JJMIT AREA=1.7857142857142858
B_AND_1|13 _AND_1|25 _AND_1|26 JJMIT AREA=2.5
B_AND_1|14 _AND_1|31 _AND_1|32 JJMIT AREA=2.5
B_AND_1|15 _AND_1|28 _AND_1|29 JJMIT AREA=2.5
I_AND_1|B1 0 _AND_1|3  PWL(0 0 5e-12 0.000175)
I_AND_1|B2 0 _AND_1|7  PWL(0 0 5e-12 0.000175)
I_AND_1|B3 0 _AND_1|16  PWL(0 0 5e-12 0.000175)
I_AND_1|B4 0 _AND_1|20  PWL(0 0 5e-12 0.000175)
I_AND_1|B5 0 _AND_1|27  PWL(0 0 5e-12 0.000175)
I_AND_1|B6 0 _AND_1|33  PWL(0 0 5e-12 0.000175)
I_AND_1|B7 0 _AND_1|30  PWL(0 0 5e-12 0.000175)
L_AND_1|B1 _AND_1|3 _AND_1|1  2e-12
L_AND_1|B2 _AND_1|7 _AND_1|5  2e-12
L_AND_1|B3 _AND_1|16 _AND_1|14  2e-12
L_AND_1|B4 _AND_1|20 _AND_1|18  2e-12
L_AND_1|B5 _AND_1|27 _AND_1|25  2e-12
L_AND_1|B6 _AND_1|30 _AND_1|28  2e-12
L_AND_1|B7 _AND_1|33 _AND_1|31  2e-12
L_AND_1|P1 _AND_1|2 0  2e-13
L_AND_1|P3 _AND_1|6 0  2e-13
L_AND_1|P5 _AND_1|11 0  2e-13
L_AND_1|P7 _AND_1|15 0  2e-13
L_AND_1|P9 _AND_1|19 0  2e-13
L_AND_1|P11 _AND_1|23 0  2e-13
L_AND_1|P13 _AND_1|26 0  2e-13
L_AND_1|P14 _AND_1|32 0  2e-13
L_AND_1|P15 _AND_1|29 0  2e-13
L_AND_1|1 A _AND_1|1  2.067833848e-12
L_AND_1|2 _AND_1|1 _AND_1|4  4.135667696e-12
L_AND_1|3 _AND_1|5 _AND_1|8  8.271335392e-12
L_AND_1|4 _AND_1|9 _AND_1|10  1e-12
L_AND_1|5 _AND_1|8 _AND_1|12  4.135667696e-12
L_AND_1|6 B _AND_1|14  2.067833848e-12
L_AND_1|7 _AND_1|14 _AND_1|17  4.135667696e-12
L_AND_1|8 _AND_1|18 _AND_1|21  8.271335392e-12
L_AND_1|9 _AND_1|22 _AND_1|10  1e-12
L_AND_1|10 _AND_1|21 _AND_1|24  4.135667696e-12
L_AND_1|11 T1 _AND_1|25  2.067833848e-12
L_AND_1|12 _AND_1|25 _AND_1|31  4.135667696e-12
L_AND_1|13 _AND_1|31 _AND_1|10  1e-12
L_AND_1|14 _AND_1|13 _AND_1|28  1e-12
L_AND_1|15 _AND_1|28 AB0  2.067833848e-12
R_AND_1|B1 _AND_1|1 _AND_1|101  2.7439617672
L_AND_1|RB1 _AND_1|101 0  1.550338398468e-12
R_AND_1|B2 _AND_1|4 _AND_1|104  3.84154647408
L_AND_1|RB2 _AND_1|104 _AND_1|5  2.1704737578552e-12
R_AND_1|B3 _AND_1|5 _AND_1|105  2.7439617672
L_AND_1|RB3 _AND_1|105 0  1.550338398468e-12
R_AND_1|B4 _AND_1|8 _AND_1|109  3.84154647408
L_AND_1|RB4 _AND_1|109 _AND_1|9  2.1704737578552e-12
R_AND_1|B5 _AND_1|8 _AND_1|108  2.7439617672
L_AND_1|RB5 _AND_1|108 0  1.550338398468e-12
R_AND_1|B6 _AND_1|12 _AND_1|112  3.84154647408
L_AND_1|RB6 _AND_1|112 _AND_1|13  2.1704737578552e-12
R_AND_1|B7 _AND_1|14 _AND_1|114  2.7439617672
L_AND_1|RB7 _AND_1|114 0  1.550338398468e-12
R_AND_1|B8 _AND_1|17 _AND_1|117  3.84154647408
L_AND_1|RB8 _AND_1|117 _AND_1|18  2.1704737578552e-12
R_AND_1|B9 _AND_1|18 _AND_1|118  2.7439617672
L_AND_1|RB9 _AND_1|118 0  1.550338398468e-12
R_AND_1|B10 _AND_1|21 _AND_1|122  3.84154647408
L_AND_1|RB10 _AND_1|122 _AND_1|22  2.1704737578552e-12
R_AND_1|B11 _AND_1|21 _AND_1|121  2.7439617672
L_AND_1|RB11 _AND_1|121 0  1.550338398468e-12
R_AND_1|B12 _AND_1|24 _AND_1|124  3.84154647408
L_AND_1|RB12 _AND_1|124 _AND_1|13  2.1704737578552e-12
R_AND_1|B13 _AND_1|25 _AND_1|125  2.7439617672
L_AND_1|RB13 _AND_1|125 0  1.550338398468e-12
R_AND_1|B14 _AND_1|31 _AND_1|131  2.7439617672
L_AND_1|RB14 _AND_1|131 0  1.550338398468e-12
R_AND_1|B15 _AND_1|28 _AND_1|128  2.7439617672
L_AND_1|RB15 _AND_1|128 0  1.550338398468e-12
B_AND_2|1 _AND_2|1 _AND_2|2 JJMIT AREA=2.5
B_AND_2|2 _AND_2|4 _AND_2|5 JJMIT AREA=1.7857142857142858
B_AND_2|3 _AND_2|5 _AND_2|6 JJMIT AREA=2.5
B_AND_2|4 _AND_2|8 _AND_2|9 JJMIT AREA=1.7857142857142858
B_AND_2|5 _AND_2|8 _AND_2|11 JJMIT AREA=2.5
B_AND_2|6 _AND_2|12 _AND_2|13 JJMIT AREA=1.7857142857142858
B_AND_2|7 _AND_2|14 _AND_2|15 JJMIT AREA=2.5
B_AND_2|8 _AND_2|17 _AND_2|18 JJMIT AREA=1.7857142857142858
B_AND_2|9 _AND_2|18 _AND_2|19 JJMIT AREA=2.5
B_AND_2|10 _AND_2|21 _AND_2|22 JJMIT AREA=1.7857142857142858
B_AND_2|11 _AND_2|21 _AND_2|23 JJMIT AREA=2.5
B_AND_2|12 _AND_2|24 _AND_2|13 JJMIT AREA=1.7857142857142858
B_AND_2|13 _AND_2|25 _AND_2|26 JJMIT AREA=2.5
B_AND_2|14 _AND_2|31 _AND_2|32 JJMIT AREA=2.5
B_AND_2|15 _AND_2|28 _AND_2|29 JJMIT AREA=2.5
I_AND_2|B1 0 _AND_2|3  PWL(0 0 5e-12 0.000175)
I_AND_2|B2 0 _AND_2|7  PWL(0 0 5e-12 0.000175)
I_AND_2|B3 0 _AND_2|16  PWL(0 0 5e-12 0.000175)
I_AND_2|B4 0 _AND_2|20  PWL(0 0 5e-12 0.000175)
I_AND_2|B5 0 _AND_2|27  PWL(0 0 5e-12 0.000175)
I_AND_2|B6 0 _AND_2|33  PWL(0 0 5e-12 0.000175)
I_AND_2|B7 0 _AND_2|30  PWL(0 0 5e-12 0.000175)
L_AND_2|B1 _AND_2|3 _AND_2|1  2e-12
L_AND_2|B2 _AND_2|7 _AND_2|5  2e-12
L_AND_2|B3 _AND_2|16 _AND_2|14  2e-12
L_AND_2|B4 _AND_2|20 _AND_2|18  2e-12
L_AND_2|B5 _AND_2|27 _AND_2|25  2e-12
L_AND_2|B6 _AND_2|30 _AND_2|28  2e-12
L_AND_2|B7 _AND_2|33 _AND_2|31  2e-12
L_AND_2|P1 _AND_2|2 0  2e-13
L_AND_2|P3 _AND_2|6 0  2e-13
L_AND_2|P5 _AND_2|11 0  2e-13
L_AND_2|P7 _AND_2|15 0  2e-13
L_AND_2|P9 _AND_2|19 0  2e-13
L_AND_2|P11 _AND_2|23 0  2e-13
L_AND_2|P13 _AND_2|26 0  2e-13
L_AND_2|P14 _AND_2|32 0  2e-13
L_AND_2|P15 _AND_2|29 0  2e-13
L_AND_2|1 C _AND_2|1  2.067833848e-12
L_AND_2|2 _AND_2|1 _AND_2|4  4.135667696e-12
L_AND_2|3 _AND_2|5 _AND_2|8  8.271335392e-12
L_AND_2|4 _AND_2|9 _AND_2|10  1e-12
L_AND_2|5 _AND_2|8 _AND_2|12  4.135667696e-12
L_AND_2|6 D _AND_2|14  2.067833848e-12
L_AND_2|7 _AND_2|14 _AND_2|17  4.135667696e-12
L_AND_2|8 _AND_2|18 _AND_2|21  8.271335392e-12
L_AND_2|9 _AND_2|22 _AND_2|10  1e-12
L_AND_2|10 _AND_2|21 _AND_2|24  4.135667696e-12
L_AND_2|11 T1 _AND_2|25  2.067833848e-12
L_AND_2|12 _AND_2|25 _AND_2|31  4.135667696e-12
L_AND_2|13 _AND_2|31 _AND_2|10  1e-12
L_AND_2|14 _AND_2|13 _AND_2|28  1e-12
L_AND_2|15 _AND_2|28 CD0  2.067833848e-12
R_AND_2|B1 _AND_2|1 _AND_2|101  2.7439617672
L_AND_2|RB1 _AND_2|101 0  1.550338398468e-12
R_AND_2|B2 _AND_2|4 _AND_2|104  3.84154647408
L_AND_2|RB2 _AND_2|104 _AND_2|5  2.1704737578552e-12
R_AND_2|B3 _AND_2|5 _AND_2|105  2.7439617672
L_AND_2|RB3 _AND_2|105 0  1.550338398468e-12
R_AND_2|B4 _AND_2|8 _AND_2|109  3.84154647408
L_AND_2|RB4 _AND_2|109 _AND_2|9  2.1704737578552e-12
R_AND_2|B5 _AND_2|8 _AND_2|108  2.7439617672
L_AND_2|RB5 _AND_2|108 0  1.550338398468e-12
R_AND_2|B6 _AND_2|12 _AND_2|112  3.84154647408
L_AND_2|RB6 _AND_2|112 _AND_2|13  2.1704737578552e-12
R_AND_2|B7 _AND_2|14 _AND_2|114  2.7439617672
L_AND_2|RB7 _AND_2|114 0  1.550338398468e-12
R_AND_2|B8 _AND_2|17 _AND_2|117  3.84154647408
L_AND_2|RB8 _AND_2|117 _AND_2|18  2.1704737578552e-12
R_AND_2|B9 _AND_2|18 _AND_2|118  2.7439617672
L_AND_2|RB9 _AND_2|118 0  1.550338398468e-12
R_AND_2|B10 _AND_2|21 _AND_2|122  3.84154647408
L_AND_2|RB10 _AND_2|122 _AND_2|22  2.1704737578552e-12
R_AND_2|B11 _AND_2|21 _AND_2|121  2.7439617672
L_AND_2|RB11 _AND_2|121 0  1.550338398468e-12
R_AND_2|B12 _AND_2|24 _AND_2|124  3.84154647408
L_AND_2|RB12 _AND_2|124 _AND_2|13  2.1704737578552e-12
R_AND_2|B13 _AND_2|25 _AND_2|125  2.7439617672
L_AND_2|RB13 _AND_2|125 0  1.550338398468e-12
R_AND_2|B14 _AND_2|31 _AND_2|131  2.7439617672
L_AND_2|RB14 _AND_2|131 0  1.550338398468e-12
R_AND_2|B15 _AND_2|28 _AND_2|128  2.7439617672
L_AND_2|RB15 _AND_2|128 0  1.550338398468e-12
BD1|1 D1|1 D1|2 JJMIT AREA=2.5
BD1|2 D1|4 D1|5 JJMIT AREA=2.5
BD1|3 D1|7 D1|8 JJMIT AREA=2.5
BD1|4 D1|10 D1|11 JJMIT AREA=2.5
ID1|B1 0 D1|3  PWL(0 0 5e-12 0.000175)
ID1|B2 0 D1|6  PWL(0 0 5e-12 0.0002375)
ID1|B3 0 D1|9  PWL(0 0 5e-12 0.0002375)
ID1|B4 0 D1|12  PWL(0 0 5e-12 0.000175)
LD1|1 AB0 D1|1  2.067833848e-12
LD1|2 D1|1 D1|4  4.135667696e-12
LD1|3 D1|4 D1|7  4.135667696e-12
LD1|4 D1|7 D1|10  4.135667696e-12
LD1|5 D1|10 AB1  2.067833848e-12
LD1|P1 D1|2 0  5e-13
LD1|P2 D1|5 0  5e-13
LD1|P3 D1|8 0  5e-13
LD1|P4 D1|11 0  5e-13
LD1|B1 D1|1 D1|3  2e-12
LD1|B2 D1|4 D1|6  2e-12
LD1|B3 D1|7 D1|9  2e-12
LD1|B4 D1|10 D1|12  2e-12
RD1|B1 D1|1 D1|101  2.7439617672
RD1|B2 D1|4 D1|104  2.7439617672
RD1|B3 D1|7 D1|107  2.7439617672
RD1|B4 D1|10 D1|110  2.7439617672
LD1|RB1 D1|101 0  2.050338398468e-12
LD1|RB2 D1|104 0  2.050338398468e-12
LD1|RB3 D1|107 0  2.050338398468e-12
LD1|RB4 D1|110 0  2.050338398468e-12
BD2|1 D2|1 D2|2 JJMIT AREA=2.5
BD2|2 D2|4 D2|5 JJMIT AREA=2.5
BD2|3 D2|7 D2|8 JJMIT AREA=2.5
BD2|4 D2|10 D2|11 JJMIT AREA=2.5
ID2|B1 0 D2|3  PWL(0 0 5e-12 0.000175)
ID2|B2 0 D2|6  PWL(0 0 5e-12 0.0002375)
ID2|B3 0 D2|9  PWL(0 0 5e-12 0.0002375)
ID2|B4 0 D2|12  PWL(0 0 5e-12 0.000175)
LD2|1 CD0 D2|1  2.067833848e-12
LD2|2 D2|1 D2|4  4.135667696e-12
LD2|3 D2|4 D2|7  4.135667696e-12
LD2|4 D2|7 D2|10  4.135667696e-12
LD2|5 D2|10 CD1  2.067833848e-12
LD2|P1 D2|2 0  5e-13
LD2|P2 D2|5 0  5e-13
LD2|P3 D2|8 0  5e-13
LD2|P4 D2|11 0  5e-13
LD2|B1 D2|1 D2|3  2e-12
LD2|B2 D2|4 D2|6  2e-12
LD2|B3 D2|7 D2|9  2e-12
LD2|B4 D2|10 D2|12  2e-12
RD2|B1 D2|1 D2|101  2.7439617672
RD2|B2 D2|4 D2|104  2.7439617672
RD2|B3 D2|7 D2|107  2.7439617672
RD2|B4 D2|10 D2|110  2.7439617672
LD2|RB1 D2|101 0  2.050338398468e-12
LD2|RB2 D2|104 0  2.050338398468e-12
LD2|RB3 D2|107 0  2.050338398468e-12
LD2|RB4 D2|110 0  2.050338398468e-12
BD3|1 D3|1 D3|2 JJMIT AREA=2.5
BD3|2 D3|6 D3|7 JJMIT AREA=2.5
ID3|B1 0 D3|5  0.00035
LD3|1 AB1 D3|1  2.067833848e-12
LD3|2 D3|1 D3|4  2.067833848e-12
LD3|3 D3|4 D3|6  2.067833848e-12
LD3|4 D3|6 AB  2.067833848e-12
LD3|P1 D3|2 0  2e-13
LD3|P2 D3|7 0  2e-13
LD3|B1 D3|5 D3|4  2e-12
RD3|B1 D3|1 D3|3  2.7439617672
RD3|B2 D3|6 D3|8  2.7439617672
LD3|RB1 D3|3 0  1.750338398468e-12
LD3|RB2 D3|8 0  1.750338398468e-12
BD4|1 D4|1 D4|2 JJMIT AREA=2.5
BD4|2 D4|6 D4|7 JJMIT AREA=2.5
ID4|B1 0 D4|5  0.00035
LD4|1 CD1 D4|1  2.067833848e-12
LD4|2 D4|1 D4|4  2.067833848e-12
LD4|3 D4|4 D4|6  2.067833848e-12
LD4|4 D4|6 CD  2.067833848e-12
LD4|P1 D4|2 0  2e-13
LD4|P2 D4|7 0  2e-13
LD4|B1 D4|5 D4|4  2e-12
RD4|B1 D4|1 D4|3  2.7439617672
RD4|B2 D4|6 D4|8  2.7439617672
LD4|RB1 D4|3 0  1.750338398468e-12
LD4|RB2 D4|8 0  1.750338398468e-12
IT2|T 0 T2  PWL(0 0 2.97e-10 0 3e-10 0.0005 3.03e-10 0 5.97e-10 0 6e-10 0.0005 6.03e-10 0 8.97e-10 0 9e-10 0.0005 9.03e-10 0 1.197e-09 0 1.2e-09 0.0005 1.203e-09 0 1.497e-09 0 1.5e-09 0.0005 1.503e-09 0 1.797e-09 0 1.8e-09 0.0005 1.803e-09 0 2.097e-09 0 2.1e-09 0.0005 2.103e-09 0 2.397e-09 0 2.4e-09 0.0005 2.403e-09 0 2.697e-09 0 2.7e-09 0.0005 2.703e-09 0 2.997e-09 0 3e-09 0.0005 3.003e-09 0 3.297e-09 0 3.3e-09 0.0005 3.303e-09 0 3.597e-09 0 3.6e-09 0.0005 3.603e-09 0 3.897e-09 0 3.9e-09 0.0005 3.903e-09 0 4.197e-09 0 4.2e-09 0.0005 4.203e-09 0 4.497e-09 0 4.5e-09 0.0005 4.503e-09 0 4.797e-09 0 4.8e-09 0.0005 4.803e-09 0 5.097e-09 0 5.1e-09 0.0005 5.103e-09 0 5.397e-09 0 5.4e-09 0.0005 5.403e-09 0 5.697e-09 0 5.7e-09 0.0005 5.703e-09 0 5.997e-09 0 6e-09 0.0005 6.003e-09 0 6.297e-09 0 6.3e-09 0.0005 6.303e-09 0 6.597e-09 0 6.6e-09 0.0005 6.603e-09 0 6.897e-09 0 6.9e-09 0.0005 6.903e-09 0 7.197e-09 0 7.2e-09 0.0005 7.203e-09 0 7.497e-09 0 7.5e-09 0.0005 7.503e-09 0 7.797e-09 0 7.8e-09 0.0005 7.803e-09 0 8.097e-09 0 8.1e-09 0.0005 8.103e-09 0 8.397e-09 0 8.4e-09 0.0005 8.403e-09 0 8.697e-09 0 8.7e-09 0.0005 8.703e-09 0 8.997e-09 0 9e-09 0.0005 9.003e-09 0 9.297e-09 0 9.3e-09 0.0005 9.303e-09 0 9.597e-09 0 9.6e-09 0.0005 9.603e-09 0 9.897e-09 0 9.9e-09 0.0005 9.903e-09 0 1.0197e-08 0 1.02e-08 0.0005 1.0203e-08 0 1.0497e-08 0 1.05e-08 0.0005 1.0503e-08 0 1.0797e-08 0 1.08e-08 0.0005 1.0803e-08 0 1.1097e-08 0 1.11e-08 0.0005 1.1103e-08 0 1.1397e-08 0 1.14e-08 0.0005 1.1403e-08 0 1.1697e-08 0 1.17e-08 0.0005 1.1703e-08 0)
B_XOR|1 _XOR|1 _XOR|2 JJMIT AREA=2.5
B_XOR|2 _XOR|4 _XOR|5 JJMIT AREA=2.5
B_XOR|3 _XOR|25 _XOR|6 JJMIT AREA=2.5
B_XOR|4 _XOR|9 _XOR|10 JJMIT AREA=2.5
B_XOR|5 _XOR|12 _XOR|13 JJMIT AREA=2.5
B_XOR|6 _XOR|26 _XOR|14 JJMIT AREA=2.5
B_XOR|7 _XOR|27 _XOR|16 JJMIT AREA=2.0
B_XOR|8 _XOR|17 _XOR|18 JJMIT AREA=2.5
B_XOR|9 _XOR|20 _XOR|16 JJMIT AREA=2.0
B_XOR|10 _XOR|16 _XOR|21 JJMIT AREA=2.5
B_XOR|11 _XOR|22 _XOR|23 JJMIT AREA=2.5
I_XOR|B1 0 _XOR|3  0.00017499999999999997
I_XOR|B2 0 _XOR|7  0.00017499999999999997
I_XOR|B3 0 _XOR|11  0.00017499999999999997
I_XOR|B4 0 _XOR|15  0.00017499999999999997
I_XOR|B5 0 _XOR|19  0.00017499999999999997
I_XOR|B6 0 _XOR|24  0.00017499999999999997
L_XOR|B1 _XOR|3 _XOR|1  2e-12
L_XOR|B2 _XOR|7 _XOR|6  2e-12
L_XOR|B3 _XOR|11 _XOR|9  2e-12
L_XOR|B4 _XOR|15 _XOR|14  2e-12
L_XOR|B5 _XOR|19 _XOR|17  2e-12
L_XOR|B6 _XOR|24 _XOR|22  2e-12
L_XOR|1 AB _XOR|1  2.067833848e-12
L_XOR|2 _XOR|1 _XOR|4  4.135667696e-12
L_XOR|3 _XOR|4 _XOR|25  1.2e-12
L_XOR|4 _XOR|6 _XOR|8  8.271335392e-12
L_XOR|5 CD _XOR|9  2.067833848e-12
L_XOR|6 _XOR|9 _XOR|12  4.135667696e-12
L_XOR|7 _XOR|12 _XOR|26  1.2e-12
L_XOR|8 _XOR|14 _XOR|8  8.271335392e-12
L_XOR|9 _XOR|8 _XOR|27  1.2e-12
L_XOR|10 T2 _XOR|17  2.067833848e-12
L_XOR|11 _XOR|17 _XOR|20  4.135667696e-12
L_XOR|12 _XOR|16 _XOR|22  4.135667696e-12
L_XOR|13 _XOR|22 ABXCD0  2.067833848e-12
L_XOR|P1 _XOR|2 0  5e-13
L_XOR|P2 _XOR|5 0  5e-13
L_XOR|P4 _XOR|10 0  5e-13
L_XOR|P5 _XOR|13 0  5e-13
L_XOR|P8 _XOR|18 0  5e-13
L_XOR|P10 _XOR|21 0  5e-13
L_XOR|P11 _XOR|23 0  5e-13
R_XOR|B1 _XOR|1 _XOR|101  2.7439617672
L_XOR|RB1 _XOR|101 0  2.050338398468e-12
R_XOR|B2 _XOR|4 _XOR|104  2.7439617672
L_XOR|RB2 _XOR|104 0  2.050338398468e-12
R_XOR|B3 _XOR|4 _XOR|106  2.7439617672
L_XOR|RB3 _XOR|106 _XOR|6  2.050338398468e-12
R_XOR|B4 _XOR|9 _XOR|109  2.7439617672
L_XOR|RB4 _XOR|109 0  2.050338398468e-12
R_XOR|B5 _XOR|12 _XOR|112  2.7439617672
L_XOR|RB5 _XOR|112 0  2.050338398468e-12
R_XOR|B6 _XOR|12 _XOR|114  2.7439617672
L_XOR|RB6 _XOR|114 _XOR|14  2.050338398468e-12
R_XOR|B7 _XOR|8 _XOR|108  3.429952209
L_XOR|RB7 _XOR|108 _XOR|16  2.437922998085e-12
R_XOR|B8 _XOR|17 _XOR|117  2.7439617672
L_XOR|RB8 _XOR|117 0  2.050338398468e-12
R_XOR|B9 _XOR|20 _XOR|120  3.429952209
L_XOR|RB9 _XOR|120 _XOR|16  2.437922998085e-12
R_XOR|B10 _XOR|16 _XOR|116  2.7439617672
L_XOR|RB10 _XOR|116 0  2.050338398468e-12
R_XOR|B11 _XOR|22 _XOR|122  2.7439617672
L_XOR|RB11 _XOR|122 0  2.050338398468e-12
LJTLOUT|1 ABXCD0 JTLOUT|1  2.067833848e-12
LJTLOUT|2 JTLOUT|1 JTLOUT|4  2.067833848e-12
LJTLOUT|3 JTLOUT|4 JTLOUT|6  2.067833848e-12
LJTLOUT|4 JTLOUT|6 ABXCD  2.067833848e-12
BJTLOUT|1|1 JTLOUT|1 JTLOUT|1|MID_SERIES JJMIT AREA=2.5
LJTLOUT|1|P JTLOUT|1|MID_SERIES 0  2e-13
RJTLOUT|1|B JTLOUT|1 JTLOUT|1|MID_SHUNT  2.7439617672
LJTLOUT|1|RB JTLOUT|1|MID_SHUNT 0  1.750338398468e-12
LJTLOUT|B|B JTLOUT|4 JTLOUT|B|MID  2e-12
IJTLOUT|B|B 0 JTLOUT|B|MID  0.0005
BJTLOUT|2|1 JTLOUT|6 JTLOUT|2|MID_SERIES JJMIT AREA=2.5
LJTLOUT|2|P JTLOUT|2|MID_SERIES 0  2e-13
RJTLOUT|2|B JTLOUT|6 JTLOUT|2|MID_SHUNT  2.7439617672
LJTLOUT|2|RB JTLOUT|2|MID_SHUNT 0  1.750338398468e-12
.print DEVI ROUT
.print DEVI IT1|T
.print DEVI IDATA_A|A
.print DEVI IDATA_B|B
.print DEVI IDATA_C|T
.print DEVI IDATA_D|T
.print DEVI B_AND_1|1
.print DEVI B_AND_1|2
.print DEVI B_AND_1|3
.print DEVI B_AND_1|4
.print DEVI B_AND_1|5
.print DEVI B_AND_1|6
.print DEVI B_AND_1|7
.print DEVI B_AND_1|8
.print DEVI B_AND_1|9
.print DEVI B_AND_1|10
.print DEVI B_AND_1|11
.print DEVI B_AND_1|12
.print DEVI B_AND_1|13
.print DEVI B_AND_1|14
.print DEVI B_AND_1|15
.print DEVI I_AND_1|B1
.print DEVI I_AND_1|B2
.print DEVI I_AND_1|B3
.print DEVI I_AND_1|B4
.print DEVI I_AND_1|B5
.print DEVI I_AND_1|B6
.print DEVI I_AND_1|B7
.print DEVI L_AND_1|B1
.print DEVI L_AND_1|B2
.print DEVI L_AND_1|B3
.print DEVI L_AND_1|B4
.print DEVI L_AND_1|B5
.print DEVI L_AND_1|B6
.print DEVI L_AND_1|B7
.print DEVI L_AND_1|P1
.print DEVI L_AND_1|P3
.print DEVI L_AND_1|P5
.print DEVI L_AND_1|P7
.print DEVI L_AND_1|P9
.print DEVI L_AND_1|P11
.print DEVI L_AND_1|P13
.print DEVI L_AND_1|P14
.print DEVI L_AND_1|P15
.print DEVI L_AND_1|1
.print DEVI L_AND_1|2
.print DEVI L_AND_1|3
.print DEVI L_AND_1|4
.print DEVI L_AND_1|5
.print DEVI L_AND_1|6
.print DEVI L_AND_1|7
.print DEVI L_AND_1|8
.print DEVI L_AND_1|9
.print DEVI L_AND_1|10
.print DEVI L_AND_1|11
.print DEVI L_AND_1|12
.print DEVI L_AND_1|13
.print DEVI L_AND_1|14
.print DEVI L_AND_1|15
.print DEVI R_AND_1|B1
.print DEVI L_AND_1|RB1
.print DEVI R_AND_1|B2
.print DEVI L_AND_1|RB2
.print DEVI R_AND_1|B3
.print DEVI L_AND_1|RB3
.print DEVI R_AND_1|B4
.print DEVI L_AND_1|RB4
.print DEVI R_AND_1|B5
.print DEVI L_AND_1|RB5
.print DEVI R_AND_1|B6
.print DEVI L_AND_1|RB6
.print DEVI R_AND_1|B7
.print DEVI L_AND_1|RB7
.print DEVI R_AND_1|B8
.print DEVI L_AND_1|RB8
.print DEVI R_AND_1|B9
.print DEVI L_AND_1|RB9
.print DEVI R_AND_1|B10
.print DEVI L_AND_1|RB10
.print DEVI R_AND_1|B11
.print DEVI L_AND_1|RB11
.print DEVI R_AND_1|B12
.print DEVI L_AND_1|RB12
.print DEVI R_AND_1|B13
.print DEVI L_AND_1|RB13
.print DEVI R_AND_1|B14
.print DEVI L_AND_1|RB14
.print DEVI R_AND_1|B15
.print DEVI L_AND_1|RB15
.print DEVI B_AND_2|1
.print DEVI B_AND_2|2
.print DEVI B_AND_2|3
.print DEVI B_AND_2|4
.print DEVI B_AND_2|5
.print DEVI B_AND_2|6
.print DEVI B_AND_2|7
.print DEVI B_AND_2|8
.print DEVI B_AND_2|9
.print DEVI B_AND_2|10
.print DEVI B_AND_2|11
.print DEVI B_AND_2|12
.print DEVI B_AND_2|13
.print DEVI B_AND_2|14
.print DEVI B_AND_2|15
.print DEVI I_AND_2|B1
.print DEVI I_AND_2|B2
.print DEVI I_AND_2|B3
.print DEVI I_AND_2|B4
.print DEVI I_AND_2|B5
.print DEVI I_AND_2|B6
.print DEVI I_AND_2|B7
.print DEVI L_AND_2|B1
.print DEVI L_AND_2|B2
.print DEVI L_AND_2|B3
.print DEVI L_AND_2|B4
.print DEVI L_AND_2|B5
.print DEVI L_AND_2|B6
.print DEVI L_AND_2|B7
.print DEVI L_AND_2|P1
.print DEVI L_AND_2|P3
.print DEVI L_AND_2|P5
.print DEVI L_AND_2|P7
.print DEVI L_AND_2|P9
.print DEVI L_AND_2|P11
.print DEVI L_AND_2|P13
.print DEVI L_AND_2|P14
.print DEVI L_AND_2|P15
.print DEVI L_AND_2|1
.print DEVI L_AND_2|2
.print DEVI L_AND_2|3
.print DEVI L_AND_2|4
.print DEVI L_AND_2|5
.print DEVI L_AND_2|6
.print DEVI L_AND_2|7
.print DEVI L_AND_2|8
.print DEVI L_AND_2|9
.print DEVI L_AND_2|10
.print DEVI L_AND_2|11
.print DEVI L_AND_2|12
.print DEVI L_AND_2|13
.print DEVI L_AND_2|14
.print DEVI L_AND_2|15
.print DEVI R_AND_2|B1
.print DEVI L_AND_2|RB1
.print DEVI R_AND_2|B2
.print DEVI L_AND_2|RB2
.print DEVI R_AND_2|B3
.print DEVI L_AND_2|RB3
.print DEVI R_AND_2|B4
.print DEVI L_AND_2|RB4
.print DEVI R_AND_2|B5
.print DEVI L_AND_2|RB5
.print DEVI R_AND_2|B6
.print DEVI L_AND_2|RB6
.print DEVI R_AND_2|B7
.print DEVI L_AND_2|RB7
.print DEVI R_AND_2|B8
.print DEVI L_AND_2|RB8
.print DEVI R_AND_2|B9
.print DEVI L_AND_2|RB9
.print DEVI R_AND_2|B10
.print DEVI L_AND_2|RB10
.print DEVI R_AND_2|B11
.print DEVI L_AND_2|RB11
.print DEVI R_AND_2|B12
.print DEVI L_AND_2|RB12
.print DEVI R_AND_2|B13
.print DEVI L_AND_2|RB13
.print DEVI R_AND_2|B14
.print DEVI L_AND_2|RB14
.print DEVI R_AND_2|B15
.print DEVI L_AND_2|RB15
.print DEVI BD1|1
.print DEVI BD1|2
.print DEVI BD1|3
.print DEVI BD1|4
.print DEVI ID1|B1
.print DEVI ID1|B2
.print DEVI ID1|B3
.print DEVI ID1|B4
.print DEVI LD1|1
.print DEVI LD1|2
.print DEVI LD1|3
.print DEVI LD1|4
.print DEVI LD1|5
.print DEVI LD1|P1
.print DEVI LD1|P2
.print DEVI LD1|P3
.print DEVI LD1|P4
.print DEVI LD1|B1
.print DEVI LD1|B2
.print DEVI LD1|B3
.print DEVI LD1|B4
.print DEVI RD1|B1
.print DEVI RD1|B2
.print DEVI RD1|B3
.print DEVI RD1|B4
.print DEVI LD1|RB1
.print DEVI LD1|RB2
.print DEVI LD1|RB3
.print DEVI LD1|RB4
.print DEVI BD2|1
.print DEVI BD2|2
.print DEVI BD2|3
.print DEVI BD2|4
.print DEVI ID2|B1
.print DEVI ID2|B2
.print DEVI ID2|B3
.print DEVI ID2|B4
.print DEVI LD2|1
.print DEVI LD2|2
.print DEVI LD2|3
.print DEVI LD2|4
.print DEVI LD2|5
.print DEVI LD2|P1
.print DEVI LD2|P2
.print DEVI LD2|P3
.print DEVI LD2|P4
.print DEVI LD2|B1
.print DEVI LD2|B2
.print DEVI LD2|B3
.print DEVI LD2|B4
.print DEVI RD2|B1
.print DEVI RD2|B2
.print DEVI RD2|B3
.print DEVI RD2|B4
.print DEVI LD2|RB1
.print DEVI LD2|RB2
.print DEVI LD2|RB3
.print DEVI LD2|RB4
.print DEVI BD3|1
.print DEVI BD3|2
.print DEVI ID3|B1
.print DEVI LD3|1
.print DEVI LD3|2
.print DEVI LD3|3
.print DEVI LD3|4
.print DEVI LD3|P1
.print DEVI LD3|P2
.print DEVI LD3|B1
.print DEVI RD3|B1
.print DEVI RD3|B2
.print DEVI LD3|RB1
.print DEVI LD3|RB2
.print DEVI BD4|1
.print DEVI BD4|2
.print DEVI ID4|B1
.print DEVI LD4|1
.print DEVI LD4|2
.print DEVI LD4|3
.print DEVI LD4|4
.print DEVI LD4|P1
.print DEVI LD4|P2
.print DEVI LD4|B1
.print DEVI RD4|B1
.print DEVI RD4|B2
.print DEVI LD4|RB1
.print DEVI LD4|RB2
.print DEVI IT2|T
.print DEVI B_XOR|1
.print DEVI B_XOR|2
.print DEVI B_XOR|3
.print DEVI B_XOR|4
.print DEVI B_XOR|5
.print DEVI B_XOR|6
.print DEVI B_XOR|7
.print DEVI B_XOR|8
.print DEVI B_XOR|9
.print DEVI B_XOR|10
.print DEVI B_XOR|11
.print DEVI I_XOR|B1
.print DEVI I_XOR|B2
.print DEVI I_XOR|B3
.print DEVI I_XOR|B4
.print DEVI I_XOR|B5
.print DEVI I_XOR|B6
.print DEVI L_XOR|B1
.print DEVI L_XOR|B2
.print DEVI L_XOR|B3
.print DEVI L_XOR|B4
.print DEVI L_XOR|B5
.print DEVI L_XOR|B6
.print DEVI L_XOR|1
.print DEVI L_XOR|2
.print DEVI L_XOR|3
.print DEVI L_XOR|4
.print DEVI L_XOR|5
.print DEVI L_XOR|6
.print DEVI L_XOR|7
.print DEVI L_XOR|8
.print DEVI L_XOR|9
.print DEVI L_XOR|10
.print DEVI L_XOR|11
.print DEVI L_XOR|12
.print DEVI L_XOR|13
.print DEVI L_XOR|P1
.print DEVI L_XOR|P2
.print DEVI L_XOR|P4
.print DEVI L_XOR|P5
.print DEVI L_XOR|P8
.print DEVI L_XOR|P10
.print DEVI L_XOR|P11
.print DEVI R_XOR|B1
.print DEVI L_XOR|RB1
.print DEVI R_XOR|B2
.print DEVI L_XOR|RB2
.print DEVI R_XOR|B3
.print DEVI L_XOR|RB3
.print DEVI R_XOR|B4
.print DEVI L_XOR|RB4
.print DEVI R_XOR|B5
.print DEVI L_XOR|RB5
.print DEVI R_XOR|B6
.print DEVI L_XOR|RB6
.print DEVI R_XOR|B7
.print DEVI L_XOR|RB7
.print DEVI R_XOR|B8
.print DEVI L_XOR|RB8
.print DEVI R_XOR|B9
.print DEVI L_XOR|RB9
.print DEVI R_XOR|B10
.print DEVI L_XOR|RB10
.print DEVI R_XOR|B11
.print DEVI L_XOR|RB11
.print DEVI LJTLOUT|1
.print DEVI LJTLOUT|2
.print DEVI LJTLOUT|3
.print DEVI LJTLOUT|4
.print DEVI BJTLOUT|1|1
.print DEVI LJTLOUT|1|P
.print DEVI RJTLOUT|1|B
.print DEVI LJTLOUT|1|RB
.print DEVI LJTLOUT|B|B
.print DEVI IJTLOUT|B|B
.print DEVI BJTLOUT|2|1
.print DEVI LJTLOUT|2|P
.print DEVI RJTLOUT|2|B
.print DEVI LJTLOUT|2|RB
.print V D2|107
.print V D3|3
.print V _AND_1|128
.print V _AND_1|24
.print V D3|7
.print V _AND_1|9
.print V _AND_1|117
.print V _AND_2|32
.print V _AND_1|32
.print V _AND_1|26
.print V _AND_1|27
.print V _XOR|19
.print V D2|9
.print V CD1
.print V _AND_2|105
.print V _XOR|9
.print V _AND_2|16
.print V D
.print V D3|1
.print V _XOR|117
.print V _XOR|27
.print V _AND_2|118
.print V AB1
.print V JTLOUT|6
.print V D4|1
.print V _XOR|26
.print V _AND_1|114
.print V _AND_2|18
.print V _AND_1|5
.print V _AND_2|125
.print V _AND_2|131
.print V _AND_2|21
.print V D2|2
.print V _AND_2|11
.print V D1|1
.print V D4|6
.print V _AND_2|121
.print V _XOR|108
.print V _AND_1|1
.print V D3|8
.print V _AND_1|15
.print V _XOR|3
.print V _AND_2|112
.print V _XOR|116
.print V AB
.print V D2|10
.print V _XOR|13
.print V _XOR|5
.print V JTLOUT|1
.print V _AND_1|21
.print V _AND_2|5
.print V _XOR|122
.print V ABXCD0
.print V _AND_2|8
.print V D1|12
.print V _XOR|114
.print V _AND_2|3
.print V _AND_2|4
.print V D3|4
.print V JTLOUT|2|MID_SERIES
.print V _AND_1|20
.print V _XOR|101
.print V _AND_1|12
.print V _AND_1|31
.print V _AND_2|23
.print V _XOR|112
.print V _AND_1|121
.print V _AND_1|6
.print V JTLOUT|1|MID_SERIES
.print V _AND_2|12
.print V _XOR|24
.print V _AND_1|23
.print V _XOR|16
.print V D2|110
.print V _XOR|23
.print V _AND_1|104
.print V _AND_2|9
.print V _AND_1|22
.print V _AND_2|15
.print V D1|10
.print V D2|12
.print V D4|4
.print V _AND_2|33
.print V _AND_2|2
.print V _AND_1|125
.print V _XOR|109
.print V ABXCD
.print V D3|5
.print V _XOR|20
.print V D3|6
.print V D2|101
.print V _AND_2|14
.print V _XOR|4
.print V D2|104
.print V D1|110
.print V _AND_1|4
.print V A
.print V D4|2
.print V _AND_1|13
.print V _XOR|25
.print V _AND_2|22
.print V _XOR|18
.print V _AND_1|131
.print V _AND_1|30
.print V _AND_2|7
.print V D4|3
.print V _XOR|120
.print V _AND_1|17
.print V D2|6
.print V B
.print V D1|7
.print V _AND_1|28
.print V T2
.print V AB0
.print V _XOR|14
.print V D1|107
.print V D4|5
.print V _AND_1|7
.print V _AND_1|25
.print V D1|104
.print V _AND_2|101
.print V _XOR|2
.print V D2|11
.print V _AND_1|109
.print V _XOR|11
.print V _AND_2|124
.print V T1
.print V D1|3
.print V D1|2
.print V _XOR|10
.print V D4|7
.print V _XOR|8
.print V _AND_1|8
.print V _AND_2|30
.print V _AND_1|112
.print V CD
.print V JTLOUT|1|MID_SHUNT
.print V _AND_2|19
.print V _XOR|1
.print V _AND_2|13
.print V _AND_2|17
.print V JTLOUT|4
.print V _AND_2|24
.print V _XOR|104
.print V CD0
.print V JTLOUT|2|MID_SHUNT
.print V _XOR|17
.print V _AND_1|105
.print V _AND_2|25
.print V D1|101
.print V _AND_1|101
.print V D1|8
.print V _XOR|12
.print V D2|1
.print V _XOR|15
.print V D1|11
.print V C
.print V _XOR|6
.print V D2|7
.print V _XOR|7
.print V _AND_1|122
.print V _AND_1|3
.print V _AND_1|118
.print V D1|9
.print V D3|2
.print V D2|5
.print V _AND_1|18
.print V _AND_1|29
.print V _AND_2|27
.print V _AND_1|11
.print V _AND_2|6
.print V _AND_2|28
.print V _AND_2|108
.print V _AND_2|31
.print V _AND_2|26
.print V _AND_2|114
.print V _AND_1|16
.print V D2|3
.print V _AND_1|14
.print V D4|8
.print V _AND_2|29
.print V _AND_2|128
.print V D1|6
.print V _AND_2|10
.print V D1|5
.print V _XOR|106
.print V _XOR|22
.print V _AND_2|109
.print V D1|4
.print V _AND_2|20
.print V _AND_1|108
.print V _AND_1|19
.print V _AND_1|33
.print V JTLOUT|B|MID
.print V _XOR|21
.print V _AND_2|1
.print V D2|4
.print V D2|8
.print V _AND_1|10
.print V _AND_2|117
.print V _AND_2|104
.print V _AND_1|124
.print V _AND_2|122
.print V _AND_1|2
.print DEVP B_AND_1|1
.print DEVP B_AND_1|2
.print DEVP B_AND_1|3
.print DEVP B_AND_1|4
.print DEVP B_AND_1|5
.print DEVP B_AND_1|6
.print DEVP B_AND_1|7
.print DEVP B_AND_1|8
.print DEVP B_AND_1|9
.print DEVP B_AND_1|10
.print DEVP B_AND_1|11
.print DEVP B_AND_1|12
.print DEVP B_AND_1|13
.print DEVP B_AND_1|14
.print DEVP B_AND_1|15
.print DEVP B_AND_2|1
.print DEVP B_AND_2|2
.print DEVP B_AND_2|3
.print DEVP B_AND_2|4
.print DEVP B_AND_2|5
.print DEVP B_AND_2|6
.print DEVP B_AND_2|7
.print DEVP B_AND_2|8
.print DEVP B_AND_2|9
.print DEVP B_AND_2|10
.print DEVP B_AND_2|11
.print DEVP B_AND_2|12
.print DEVP B_AND_2|13
.print DEVP B_AND_2|14
.print DEVP B_AND_2|15
.print DEVP BD1|1
.print DEVP BD1|2
.print DEVP BD1|3
.print DEVP BD1|4
.print DEVP BD2|1
.print DEVP BD2|2
.print DEVP BD2|3
.print DEVP BD2|4
.print DEVP BD3|1
.print DEVP BD3|2
.print DEVP BD4|1
.print DEVP BD4|2
.print DEVP B_XOR|1
.print DEVP B_XOR|2
.print DEVP B_XOR|3
.print DEVP B_XOR|4
.print DEVP B_XOR|5
.print DEVP B_XOR|6
.print DEVP B_XOR|7
.print DEVP B_XOR|8
.print DEVP B_XOR|9
.print DEVP B_XOR|10
.print DEVP B_XOR|11
.print DEVP BJTLOUT|1|1
.print DEVP BJTLOUT|2|1
