
.include /Users/brainkz/Documents/GitHub/SFQ_gate_Exploration/jj_library.cir
.include /Users/brainkz/Documents/GitHub/SFQ/sunmagnetics_library.cir



.subckt	pg_init	a	b	clk	pout	gout
  * Need	3	clocks	here
  X_spl_a	a	a1	a2	spl2
  X_spl_b	b	b1	b2	spl2

  X_dff_a	a1	clk	a1_sync	dff
  X_dff_b	b1	clk	b1_sync	dff
  
  X_xor	a2	b2	clk	pout	xor
  X_and	a1_sync	b1_sync	gout	merge	mbias=0.2
.ends

.subckt	B_pg	P0  G0  P1  G1  clk pout    gout
  * Need 4 clocks here
  X_spl_g1	G1	G1_copy_1	G1_copy_2	spl2
  X_spl_p1	P1	P1_copy_1	P1_copy_2	spl2
  
  X_pg	P1_copy_1	G1_copy_1	pg	merge	mbias=1
  X_gg	G0          G1_copy_2	gg	merge	mbias=1

  X_dff_p0	P0	        clk	P0_sync	dff
  X_dff_p1	P1_copy_2	clk	P1_sync	dff
  X_dff_pg    pg          clk pg_sync dff
  X_dff_gg    gg          clk gg_sync dff

  X_and_g	pg_sync	gg_sync	gout	merge	mbias=0.2
  X_and_p	P0_sync	P1_sync	pout	merge	mbias=0.2
.ends

.subckt	W_pg	pin  gin  clk pout    gout
  * Need 2 clocks here
  Xp	    pin     clk	    pout	dff
  Xg	    gin     clk	    gout	dff
.ends

.subckt	B_g         G0  P1  G1  clk          gout
  * Need 2 clocks here
  X_spl_g1	G1	G1_copy_1	G1_copy_2	spl2
  
  X_pg	P1   G1_copy_1	pg	merge	mbias=1
  X_gg	G0   G1_copy_2	gg	merge	mbias=1

  X_dff_pg    pg          clk pg_sync dff
  X_dff_gg    gg          clk gg_sync dff

  X_and_g	pg_sync	gg_sync	gout	merge	mbias=0.2
.ends

.param tclock=200e-12
.param OS=tclock/40
.param step=0.08
*  Input signals
  Xa0_ a0_ data_sig_a_r clk_offset=OS do_factor=step*2+step*0 Tck=tclock
  Xb0_ b0_ data_sig_b_r clk_offset=OS do_factor=step*3+step*0 Tck=tclock
  Xa1_ a1_ data_sig_c_r clk_offset=OS do_factor=step*4+step*0 Tck=tclock
  Xb1_ b1_ data_sig_d_r clk_offset=OS do_factor=step*5+step*0 Tck=tclock
  Xa2_ a2_ data_sig_e_r clk_offset=OS do_factor=step*6+step*0 Tck=tclock
  Xb2_ b2_ data_sig_f_r clk_offset=OS do_factor=step*7+step*0 Tck=tclock
  Xa3_ a3_ data_sig_g_r clk_offset=OS do_factor=step*8+step*0 Tck=tclock
  Xb3_ b3_ data_sig_h_r clk_offset=OS do_factor=step*9+step*0 Tck=tclock
* 
* Cycle 0
  xt00_ T00_ clk_sig clk_offset=OS*4 factor=3 Tck=tclock
  Xi0_ a0_ b0_ T00_ iP0_0_ iG0_0_ pg_init
  
  Xt01_ T01_ clk_sig clk_offset=OS*4 factor=3 Tck=tclock
  Xi1_ a1_ b1_ T01_ iP1_0_ iG1_0_ pg_init
  
  Xt02_ T02_ clk_sig clk_offset=OS*4 factor=3 Tck=tclock
  Xi2_ a2_ b2_ T02_ iP2_0_ iG2_0_ pg_init
  
  Xt03_ T03_ clk_sig clk_offset=OS*4 factor=3 Tck=tclock
  Xi3_ a3_ b3_ T03_ iP3_0_ iG3_0_ pg_init
* 

*  Output Resistors
*   R_ip0_     iP0_0_  0   1
*   R_ig0_     iG0_0_  0   1
*   R_ip1_     iP1_0_  0   1
*   R_ig1_     iG1_0_  0   1
*   R_ip2_     iP2_0_  0   1
*   R_ig2_     iG2_0_  0   1
*   R_ip3_     iP3_0_  0   1
*   R_ig3_     iG3_0_  0   1
*   .tran 1e-12 64000e-12
*   .end
* 
* Splitters at level 0
  * Splitting 0
*   Xspl_iP0_0 iP0_0 iP0_0_to0 iP0_0_to1           spl2
  Xspl_iG0_0_ iG0_0_ iG0_0_to0_ iG0_0_to1_           spl2
  * Splitting 1
  Xspl_iP1_0_ iP1_0_ iP1_0_to1_           iP1_0_out_ spl2
  * Splitting 2
  Xspl_iP2_0_ iP2_0_ iP2_0_to2_ iP2_0_to3_ iP2_0_out_ spl3
  Xspl_iG2_0_ iG2_0_ iG2_0_to2_ iG2_0_to3_           spl2
  * Splitting 3
  Xspl_iP3_0_ iP3_0_ iP3_0_to1_           iP3_0_out_ spl2
* 
*   
  * R_ip0_to0     iP0_0_to0  0   1
  * R_ip0_to1     iP0_0_to1  0   1
  * R_ig0_to0     iG0_0_to0  0   1
  * R_ig0_to1     iG0_0_to1  0   1
  * R_ip1_to1     iP1_0_to1  0   1
  * R_ip1_out     iP1_0_out  0   1
  * R_ip1     iP1_0  0   1
  * R_ig1     iG1_0  0   1
  * R_ip2_to2     iP2_0_to2  0   1
  * R_ip2_to3     iP2_0_to3  0   1
  * R_ip2_out     iP2_0_out  0   1
  * R_ig2_to2     iG2_0_to2  0   1
  * R_ig2_to3     iG2_0_to3  0   1
  * R_ip3_to1     iP3_0_to1  0   1
  * R_ip3_out     iP3_0_out  0   1
  * R_ig3     iG3_0  0   1
  * .tran 1e-12 64000e-12
  * .end
* 

*  Cycle 1
  Xt04_ T04_ clk_sig clk_offset=OS*3 factor=2 Tck=tclock
*   X_pg0_01 iP0_0_to0 iG0_0_to0                 T04 P0_1 G0_1 W_pg
  X_pg0_01_ iP0_0_     iG0_0_to0_                 T04_ P0_1_ G0_1_ W_pg

  Xt05_ T05_ clk_sig clk_offset=OS*3 factor=2 Tck=tclock
*   X_pg1_01 iP0_0_to1 iG0_0_to1 iP1_0_to1 iG1_0 T05 P1_1 G1_1 B_pg
  X_pg1_01_           iG0_0_to1_ iP1_0_to1_ iG1_0_ T05_      G1_1_ B_g

  Xt06_ T06_ clk_sig clk_offset=OS*3 factor=2 Tck=tclock
  X_pg2_01_ iP2_0_to2_ iG2_0_to2_                 T06_ P2_1_ G2_1_ W_pg

  Xt07_ T07_ clk_sig clk_offset=OS*3 factor=4 Tck=tclock
  X_pg3_01_ iP2_0_to3_ iG2_0_to3_ iP3_0_to1_ iG3_0_ T07_ P3_1_ G3_1_ B_pg

  Xd01_ D01_ clk_sig clk_offset=OS*3 factor=1 Tck=tclock
  X_dff_ip1_01_  iP1_0_out_   D01_ iP1_1_out_   dff

  Xd02_ D02_ clk_sig clk_offset=OS*3 factor=1 Tck=tclock
*   Xbuf_ip2_01   iP2_0_out       iP2_0_tmp     LSMITLL_BUFF
  X_dff_ip2_01_  iP2_0_out_   D02_ iP2_1_out_   dff

  Xd03_ D03_ clk_sig clk_offset=OS*3 factor=1 Tck=tclock
  X_dff_ip3_01_  iP3_0_out_   D03_ iP3_1_out_   dff
* 

* Splitters at level 1
  * Splitting 0
  * Splitting 1
*   Xspl_P1_1   P1_1    P1_1_to1    P1_1_to2    P1_1_to3    spl3
  Xspl_G1_1_   G1_1_    G1_1_to1_    G1_1_to2_    G1_1_to3_    spl3
  * Splitting 2
  * Splitting 3
* 
* 
      R_p0_1     P0_1  0   1
      R_g0_1     G0_1  0   1
      R_p1_1_to1     P1_1_to1  0   1
      R_p1_1_to2     P1_1_to2  0   1
      R_p1_1_to3     P1_1_to3  0   1
      R_g1_1_to1     G1_1_to1  0   1
      R_g1_1_to2     G1_1_to2  0   1
      R_g1_1_to3     G1_1_to3  0   1
      R_p2_1     P2_1  0   1
      R_g2_1     G2_1  0   1
      R_p3_1     P3_1  0   1
      R_g3_1     G3_1  0   1
      R_ip1_1     iP1_1_out  0   1
      R_ip2_1     iP2_1_out  0   1
      R_ip3_1     iP3_1_out  0   1
      .tran 1e-12 54000e-12
      .end
* 

*  Cycle 2
  Xt08 T08 clk_sig clk_offset=OS*2 factor=2 Tck=tclock
  X_pg0_12  P0_1      G0_1                 T08 P0_2 G0_2 W_pg

  Xt09 T09 clk_sig clk_offset=OS*2 factor=1 Tck=tclock
*   X_pg1_12  P1_1_to1  G1_1_to1             T09 P1_2 G1_2 W_pg
  X_pg1_12            G1_1_to1             T09      G1_2 dff

  Xt10 T10 clk_sig clk_offset=OS*2 factor=2 Tck=tclock
*   X_pg2_12  P1_1_to2  G1_1_to2  P2_1  G2_1 T10 P2_2 G2_2 B_pg
  X_pg2_12            G1_1_to2  P2_1  G2_1 T10      G2_2 B_g

  Xt11 T11 clk_sig clk_offset=OS*2 factor=2 Tck=tclock
*   X_pg3_12  P1_1_to3  G1_1_to3  P3_1  G3_1 T11 P3_2 G3_2 B_pg
  X_pg3_12            G1_1_to3  P3_1  G3_1 T11      G3_2 B_g

  Xd11 D11 clk_sig clk_offset=OS*2 factor=1 Tck=tclock
  X_dff_ip1_12  iP1_1_out   D11 iP1_2_out   dff

  Xd12 D12 clk_sig clk_offset=OS*2 factor=1 Tck=tclock
*   Xbuf_ip2_12   iP2_1_out       iP2_1_tmp     LSMITLL_BUFF
  X_dff_ip2_12  iP2_1_out   D12 iP2_2_out   dff

  Xd13 D13 clk_sig clk_offset=OS*2 factor=1 Tck=tclock
  X_dff_ip3_12  iP3_1_out   D13 iP3_2_out   dff 
* 
*
    * R_p0_2     P0_2  0   1
    * R_g0_2     G0_2  0   1
    * R_p1_2     P1_2  0   1
    * R_g1_2     G1_2  0   1
    * R_p2_2     P2_2  0   1
    * R_g2_2     G2_2  0   1
    * R_p3_2     P3_2  0   1
    * R_g3_2     G3_2  0   1
    * R_ip1_2     iP1_2_out  0   1
    * R_ip2_2     iP2_2_out  0   1
    * R_ip3_2     iP3_2_out  0   1
    * .tran 2e-12 54000e-12
    * .end 
*

* Final processing
  * Bit 0
  Xt12 T12 clk_sig clk_offset=OS*1 factor=1 Tck=tclock
  X_s0  P0_2                T12 s0  dff
  R_s0  s0      0   1
*   R_c1  G0_2    0   1
  Xt13 T13 clk_sig clk_offset=OS*1 factor=1 Tck=tclock
  Xbuf_G0_2_tmp   G0_2         G0_2_tmp     LSMITLL_BUFF
  Xbuf_G0_2   G0_2_tmp     G0_2_buf     jtl
  Xbuf_iP1_2_tmp iP1_2_out    iP1_2_tmp     LSMITLL_BUFF
  Xbuf_iP1_2 iP1_2_tmp    iP1_2_out_buf jtl
  X_s1	G0_2_buf	iP1_2_out_buf	T13	s1	xor t_scaling=1 main_scaling=0.8 bottom_scaling=0.8
  R_s1  s1      0   1
*   R_c2  G1_2    0   1
  Xt14 T14 clk_sig clk_offset=OS*1 factor=1 Tck=tclock
  Xbuf_G1_2_tmp   G1_2         G1_2_tmp     LSMITLL_BUFF
  Xbuf_G1_2   G1_2_tmp     G1_2_buf     jtl
  Xbuf_iP2_2_tmp iP2_2_out    iP2_2_tmp     LSMITLL_BUFF
  Xbuf_iP2_2 iP2_2_tmp    iP2_2_out_buf jtl
  X_s2	G1_2_buf	iP2_2_out_buf	T14	s2	xor t_scaling=1 main_scaling=0.8 bottom_scaling=0.8
  R_s2  s2    0   1
*   R_c3  G2_2    0   1
  Xt15 T15 clk_sig clk_offset=OS*1 factor=1 Tck=tclock
  Xbuf_G2_2_tmp   G2_2         G2_2_tmp     LSMITLL_BUFF
  Xbuf_G2_2   G2_2_tmp     G2_2_buf     jtl
*   Xbuf_iP3_2_tmp iP3_2_out    iP3_2_tmp     LSMITLL_BUFF
*   Xbuf_iP3_2 iP3_2_tmp    iP3_2_out_buf jtl
  X_s3	G2_2_tmp	iP3_2_out	T15	s3	xor t_scaling=1 main_scaling=0.9 bottom_scaling=0.9
  R_s3  s3    0   1
*   R_c4  G3_2    0   1
  Xt16 T16 clk_sig clk_offset=OS*1 factor=1 Tck=tclock
  X_s4  G3_2                T16 s4  dff
  R_s4  s4      0   1
* 
    * R_p0_2     P0_2  0   1
    * R_g0_2     G0_2  0   1
    * R_p1_2     P1_2  0   1
    * R_g1_2     G1_2  0   1
    * R_p2_2     P2_2  0   1
    * R_g2_2     G2_2  0   1
    * R_p3_2     P3_2  0   1
    * R_g3_2     G3_2  0   1
    * R_ip1_2     iP1_2_out  0   1
    * R_ip2_2     iP2_2_out  0   1
    * R_ip3_2     iP3_2_out  0   1
    * .tran 1e-12 52000e-12
    * .tran 1e-12 39000e-12
    .tran 1e-12 52000e-12
    .end 


* *   
*   R_ip0      P0_1  0   1
*   R_ig0      G0_1  0   1
*   R_ip1     iP1_0  0   1
*   R_ig1     iG1_0  0   1
*   R_ip2     iP2_0  0   1
*   R_ig2     iG2_0  0   1
*   R_ip3     iP3_0  0   1
*   R_ig3     iG3_0  0   1
* * 

